---   Background Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: smario_traspas_patron.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_MARIO_TRASPAS_BG is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_MARIO_TRASPAS_BG;

architecture BEHAVIORAL of ROM_PTABLE_MARIO_TRASPAS_BG is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table both color planes
    "00111000", --    0 -  0x0  :   56 - 0x38 -- Background 0x0
    "01001100", --    1 -  0x1  :   76 - 0x4c
    "11000110", --    2 -  0x2  :  198 - 0xc6
    "11000110", --    3 -  0x3  :  198 - 0xc6
    "11000110", --    4 -  0x4  :  198 - 0xc6
    "01100100", --    5 -  0x5  :  100 - 0x64
    "00111000", --    6 -  0x6  :   56 - 0x38
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00011000", --   16 - 0x10  :   24 - 0x18 -- Background 0x1
    "00111000", --   17 - 0x11  :   56 - 0x38
    "00011000", --   18 - 0x12  :   24 - 0x18
    "00011000", --   19 - 0x13  :   24 - 0x18
    "00011000", --   20 - 0x14  :   24 - 0x18
    "00011000", --   21 - 0x15  :   24 - 0x18
    "01111110", --   22 - 0x16  :  126 - 0x7e
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "01111100", --   32 - 0x20  :  124 - 0x7c -- Background 0x2
    "11000110", --   33 - 0x21  :  198 - 0xc6
    "00001110", --   34 - 0x22  :   14 - 0xe
    "00111100", --   35 - 0x23  :   60 - 0x3c
    "01111000", --   36 - 0x24  :  120 - 0x78
    "11100000", --   37 - 0x25  :  224 - 0xe0
    "11111110", --   38 - 0x26  :  254 - 0xfe
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "01111110", --   48 - 0x30  :  126 - 0x7e -- Background 0x3
    "00001100", --   49 - 0x31  :   12 - 0xc
    "00011000", --   50 - 0x32  :   24 - 0x18
    "00111100", --   51 - 0x33  :   60 - 0x3c
    "00000110", --   52 - 0x34  :    6 - 0x6
    "11000110", --   53 - 0x35  :  198 - 0xc6
    "01111100", --   54 - 0x36  :  124 - 0x7c
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- plane 1
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00011100", --   64 - 0x40  :   28 - 0x1c -- Background 0x4
    "00111100", --   65 - 0x41  :   60 - 0x3c
    "01101100", --   66 - 0x42  :  108 - 0x6c
    "11001100", --   67 - 0x43  :  204 - 0xcc
    "11111110", --   68 - 0x44  :  254 - 0xfe
    "00001100", --   69 - 0x45  :   12 - 0xc
    "00001100", --   70 - 0x46  :   12 - 0xc
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- plane 1
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "11111100", --   80 - 0x50  :  252 - 0xfc -- Background 0x5
    "11000000", --   81 - 0x51  :  192 - 0xc0
    "11111100", --   82 - 0x52  :  252 - 0xfc
    "00000110", --   83 - 0x53  :    6 - 0x6
    "00000110", --   84 - 0x54  :    6 - 0x6
    "11000110", --   85 - 0x55  :  198 - 0xc6
    "01111100", --   86 - 0x56  :  124 - 0x7c
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- plane 1
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00111100", --   96 - 0x60  :   60 - 0x3c -- Background 0x6
    "01100000", --   97 - 0x61  :   96 - 0x60
    "11000000", --   98 - 0x62  :  192 - 0xc0
    "11111100", --   99 - 0x63  :  252 - 0xfc
    "11000110", --  100 - 0x64  :  198 - 0xc6
    "11000110", --  101 - 0x65  :  198 - 0xc6
    "01111100", --  102 - 0x66  :  124 - 0x7c
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- plane 1
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11111110", --  112 - 0x70  :  254 - 0xfe -- Background 0x7
    "11000110", --  113 - 0x71  :  198 - 0xc6
    "00001100", --  114 - 0x72  :   12 - 0xc
    "00011000", --  115 - 0x73  :   24 - 0x18
    "00110000", --  116 - 0x74  :   48 - 0x30
    "00110000", --  117 - 0x75  :   48 - 0x30
    "00110000", --  118 - 0x76  :   48 - 0x30
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- plane 1
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "01111100", --  128 - 0x80  :  124 - 0x7c -- Background 0x8
    "11000110", --  129 - 0x81  :  198 - 0xc6
    "11000110", --  130 - 0x82  :  198 - 0xc6
    "01111100", --  131 - 0x83  :  124 - 0x7c
    "11000110", --  132 - 0x84  :  198 - 0xc6
    "11000110", --  133 - 0x85  :  198 - 0xc6
    "01111100", --  134 - 0x86  :  124 - 0x7c
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- plane 1
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01111100", --  144 - 0x90  :  124 - 0x7c -- Background 0x9
    "11000110", --  145 - 0x91  :  198 - 0xc6
    "11000110", --  146 - 0x92  :  198 - 0xc6
    "01111110", --  147 - 0x93  :  126 - 0x7e
    "00000110", --  148 - 0x94  :    6 - 0x6
    "00001100", --  149 - 0x95  :   12 - 0xc
    "01111000", --  150 - 0x96  :  120 - 0x78
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- plane 1
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00111000", --  160 - 0xa0  :   56 - 0x38 -- Background 0xa
    "01101100", --  161 - 0xa1  :  108 - 0x6c
    "11000110", --  162 - 0xa2  :  198 - 0xc6
    "11000110", --  163 - 0xa3  :  198 - 0xc6
    "11111110", --  164 - 0xa4  :  254 - 0xfe
    "11000110", --  165 - 0xa5  :  198 - 0xc6
    "11000110", --  166 - 0xa6  :  198 - 0xc6
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- plane 1
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11111100", --  176 - 0xb0  :  252 - 0xfc -- Background 0xb
    "11000110", --  177 - 0xb1  :  198 - 0xc6
    "11000110", --  178 - 0xb2  :  198 - 0xc6
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11000110", --  180 - 0xb4  :  198 - 0xc6
    "11000110", --  181 - 0xb5  :  198 - 0xc6
    "11111100", --  182 - 0xb6  :  252 - 0xfc
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- plane 1
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00111100", --  192 - 0xc0  :   60 - 0x3c -- Background 0xc
    "01100110", --  193 - 0xc1  :  102 - 0x66
    "11000000", --  194 - 0xc2  :  192 - 0xc0
    "11000000", --  195 - 0xc3  :  192 - 0xc0
    "11000000", --  196 - 0xc4  :  192 - 0xc0
    "01100110", --  197 - 0xc5  :  102 - 0x66
    "00111100", --  198 - 0xc6  :   60 - 0x3c
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- plane 1
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "11111000", --  208 - 0xd0  :  248 - 0xf8 -- Background 0xd
    "11001100", --  209 - 0xd1  :  204 - 0xcc
    "11000110", --  210 - 0xd2  :  198 - 0xc6
    "11000110", --  211 - 0xd3  :  198 - 0xc6
    "11000110", --  212 - 0xd4  :  198 - 0xc6
    "11001100", --  213 - 0xd5  :  204 - 0xcc
    "11111000", --  214 - 0xd6  :  248 - 0xf8
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- plane 1
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "11111110", --  224 - 0xe0  :  254 - 0xfe -- Background 0xe
    "11000000", --  225 - 0xe1  :  192 - 0xc0
    "11000000", --  226 - 0xe2  :  192 - 0xc0
    "11111100", --  227 - 0xe3  :  252 - 0xfc
    "11000000", --  228 - 0xe4  :  192 - 0xc0
    "11000000", --  229 - 0xe5  :  192 - 0xc0
    "11111110", --  230 - 0xe6  :  254 - 0xfe
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- plane 1
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11111110", --  240 - 0xf0  :  254 - 0xfe -- Background 0xf
    "11000000", --  241 - 0xf1  :  192 - 0xc0
    "11000000", --  242 - 0xf2  :  192 - 0xc0
    "11111100", --  243 - 0xf3  :  252 - 0xfc
    "11000000", --  244 - 0xf4  :  192 - 0xc0
    "11000000", --  245 - 0xf5  :  192 - 0xc0
    "11000000", --  246 - 0xf6  :  192 - 0xc0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- plane 1
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00111110", --  256 - 0x100  :   62 - 0x3e -- Background 0x10
    "01100000", --  257 - 0x101  :   96 - 0x60
    "11000000", --  258 - 0x102  :  192 - 0xc0
    "11001110", --  259 - 0x103  :  206 - 0xce
    "11000110", --  260 - 0x104  :  198 - 0xc6
    "01100110", --  261 - 0x105  :  102 - 0x66
    "00111110", --  262 - 0x106  :   62 - 0x3e
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- plane 1
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "11000110", --  272 - 0x110  :  198 - 0xc6 -- Background 0x11
    "11000110", --  273 - 0x111  :  198 - 0xc6
    "11000110", --  274 - 0x112  :  198 - 0xc6
    "11111110", --  275 - 0x113  :  254 - 0xfe
    "11000110", --  276 - 0x114  :  198 - 0xc6
    "11000110", --  277 - 0x115  :  198 - 0xc6
    "11000110", --  278 - 0x116  :  198 - 0xc6
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- plane 1
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "01111110", --  288 - 0x120  :  126 - 0x7e -- Background 0x12
    "00011000", --  289 - 0x121  :   24 - 0x18
    "00011000", --  290 - 0x122  :   24 - 0x18
    "00011000", --  291 - 0x123  :   24 - 0x18
    "00011000", --  292 - 0x124  :   24 - 0x18
    "00011000", --  293 - 0x125  :   24 - 0x18
    "01111110", --  294 - 0x126  :  126 - 0x7e
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- plane 1
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00011110", --  304 - 0x130  :   30 - 0x1e -- Background 0x13
    "00000110", --  305 - 0x131  :    6 - 0x6
    "00000110", --  306 - 0x132  :    6 - 0x6
    "00000110", --  307 - 0x133  :    6 - 0x6
    "11000110", --  308 - 0x134  :  198 - 0xc6
    "11000110", --  309 - 0x135  :  198 - 0xc6
    "01111100", --  310 - 0x136  :  124 - 0x7c
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- plane 1
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "11000110", --  320 - 0x140  :  198 - 0xc6 -- Background 0x14
    "11001100", --  321 - 0x141  :  204 - 0xcc
    "11011000", --  322 - 0x142  :  216 - 0xd8
    "11110000", --  323 - 0x143  :  240 - 0xf0
    "11111000", --  324 - 0x144  :  248 - 0xf8
    "11011100", --  325 - 0x145  :  220 - 0xdc
    "11001110", --  326 - 0x146  :  206 - 0xce
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- plane 1
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "01100000", --  336 - 0x150  :   96 - 0x60 -- Background 0x15
    "01100000", --  337 - 0x151  :   96 - 0x60
    "01100000", --  338 - 0x152  :   96 - 0x60
    "01100000", --  339 - 0x153  :   96 - 0x60
    "01100000", --  340 - 0x154  :   96 - 0x60
    "01100000", --  341 - 0x155  :   96 - 0x60
    "01111110", --  342 - 0x156  :  126 - 0x7e
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0 -- plane 1
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "11000110", --  352 - 0x160  :  198 - 0xc6 -- Background 0x16
    "11101110", --  353 - 0x161  :  238 - 0xee
    "11111110", --  354 - 0x162  :  254 - 0xfe
    "11111110", --  355 - 0x163  :  254 - 0xfe
    "11010110", --  356 - 0x164  :  214 - 0xd6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "11000110", --  358 - 0x166  :  198 - 0xc6
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- plane 1
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "11000110", --  368 - 0x170  :  198 - 0xc6 -- Background 0x17
    "11100110", --  369 - 0x171  :  230 - 0xe6
    "11110110", --  370 - 0x172  :  246 - 0xf6
    "11111110", --  371 - 0x173  :  254 - 0xfe
    "11011110", --  372 - 0x174  :  222 - 0xde
    "11001110", --  373 - 0x175  :  206 - 0xce
    "11000110", --  374 - 0x176  :  198 - 0xc6
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- plane 1
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "01111100", --  384 - 0x180  :  124 - 0x7c -- Background 0x18
    "11000110", --  385 - 0x181  :  198 - 0xc6
    "11000110", --  386 - 0x182  :  198 - 0xc6
    "11000110", --  387 - 0x183  :  198 - 0xc6
    "11000110", --  388 - 0x184  :  198 - 0xc6
    "11000110", --  389 - 0x185  :  198 - 0xc6
    "01111100", --  390 - 0x186  :  124 - 0x7c
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- plane 1
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "11111100", --  400 - 0x190  :  252 - 0xfc -- Background 0x19
    "11000110", --  401 - 0x191  :  198 - 0xc6
    "11000110", --  402 - 0x192  :  198 - 0xc6
    "11000110", --  403 - 0x193  :  198 - 0xc6
    "11111100", --  404 - 0x194  :  252 - 0xfc
    "11000000", --  405 - 0x195  :  192 - 0xc0
    "11000000", --  406 - 0x196  :  192 - 0xc0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- plane 1
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "01111100", --  416 - 0x1a0  :  124 - 0x7c -- Background 0x1a
    "11000110", --  417 - 0x1a1  :  198 - 0xc6
    "11000110", --  418 - 0x1a2  :  198 - 0xc6
    "11000110", --  419 - 0x1a3  :  198 - 0xc6
    "11011110", --  420 - 0x1a4  :  222 - 0xde
    "11001100", --  421 - 0x1a5  :  204 - 0xcc
    "01111010", --  422 - 0x1a6  :  122 - 0x7a
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- plane 1
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "11111100", --  432 - 0x1b0  :  252 - 0xfc -- Background 0x1b
    "11000110", --  433 - 0x1b1  :  198 - 0xc6
    "11000110", --  434 - 0x1b2  :  198 - 0xc6
    "11001110", --  435 - 0x1b3  :  206 - 0xce
    "11111000", --  436 - 0x1b4  :  248 - 0xf8
    "11011100", --  437 - 0x1b5  :  220 - 0xdc
    "11001110", --  438 - 0x1b6  :  206 - 0xce
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- plane 1
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "01111000", --  448 - 0x1c0  :  120 - 0x78 -- Background 0x1c
    "11001100", --  449 - 0x1c1  :  204 - 0xcc
    "11000000", --  450 - 0x1c2  :  192 - 0xc0
    "01111100", --  451 - 0x1c3  :  124 - 0x7c
    "00000110", --  452 - 0x1c4  :    6 - 0x6
    "11000110", --  453 - 0x1c5  :  198 - 0xc6
    "01111100", --  454 - 0x1c6  :  124 - 0x7c
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- plane 1
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "01111110", --  464 - 0x1d0  :  126 - 0x7e -- Background 0x1d
    "00011000", --  465 - 0x1d1  :   24 - 0x18
    "00011000", --  466 - 0x1d2  :   24 - 0x18
    "00011000", --  467 - 0x1d3  :   24 - 0x18
    "00011000", --  468 - 0x1d4  :   24 - 0x18
    "00011000", --  469 - 0x1d5  :   24 - 0x18
    "00011000", --  470 - 0x1d6  :   24 - 0x18
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- plane 1
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "11000110", --  480 - 0x1e0  :  198 - 0xc6 -- Background 0x1e
    "11000110", --  481 - 0x1e1  :  198 - 0xc6
    "11000110", --  482 - 0x1e2  :  198 - 0xc6
    "11000110", --  483 - 0x1e3  :  198 - 0xc6
    "11000110", --  484 - 0x1e4  :  198 - 0xc6
    "11000110", --  485 - 0x1e5  :  198 - 0xc6
    "01111100", --  486 - 0x1e6  :  124 - 0x7c
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- plane 1
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "11000110", --  496 - 0x1f0  :  198 - 0xc6 -- Background 0x1f
    "11000110", --  497 - 0x1f1  :  198 - 0xc6
    "11000110", --  498 - 0x1f2  :  198 - 0xc6
    "11101110", --  499 - 0x1f3  :  238 - 0xee
    "01111100", --  500 - 0x1f4  :  124 - 0x7c
    "00111000", --  501 - 0x1f5  :   56 - 0x38
    "00010000", --  502 - 0x1f6  :   16 - 0x10
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- plane 1
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "11000110", --  512 - 0x200  :  198 - 0xc6 -- Background 0x20
    "11000110", --  513 - 0x201  :  198 - 0xc6
    "11010110", --  514 - 0x202  :  214 - 0xd6
    "11111110", --  515 - 0x203  :  254 - 0xfe
    "11111110", --  516 - 0x204  :  254 - 0xfe
    "11101110", --  517 - 0x205  :  238 - 0xee
    "11000110", --  518 - 0x206  :  198 - 0xc6
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "11000110", --  528 - 0x210  :  198 - 0xc6 -- Background 0x21
    "11101110", --  529 - 0x211  :  238 - 0xee
    "01111100", --  530 - 0x212  :  124 - 0x7c
    "00111000", --  531 - 0x213  :   56 - 0x38
    "01111100", --  532 - 0x214  :  124 - 0x7c
    "11101110", --  533 - 0x215  :  238 - 0xee
    "11000110", --  534 - 0x216  :  198 - 0xc6
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- plane 1
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01100110", --  544 - 0x220  :  102 - 0x66 -- Background 0x22
    "01100110", --  545 - 0x221  :  102 - 0x66
    "01100110", --  546 - 0x222  :  102 - 0x66
    "00111100", --  547 - 0x223  :   60 - 0x3c
    "00011000", --  548 - 0x224  :   24 - 0x18
    "00011000", --  549 - 0x225  :   24 - 0x18
    "00011000", --  550 - 0x226  :   24 - 0x18
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- plane 1
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "11111110", --  560 - 0x230  :  254 - 0xfe -- Background 0x23
    "00001110", --  561 - 0x231  :   14 - 0xe
    "00011100", --  562 - 0x232  :   28 - 0x1c
    "00111000", --  563 - 0x233  :   56 - 0x38
    "01110000", --  564 - 0x234  :  112 - 0x70
    "11100000", --  565 - 0x235  :  224 - 0xe0
    "11111110", --  566 - 0x236  :  254 - 0xfe
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- plane 1
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x24
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- plane 1
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "11111111", --  592 - 0x250  :  255 - 0xff -- Background 0x25
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111111", --  595 - 0x253  :  255 - 0xff
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "11111111", --  598 - 0x256  :  255 - 0xff
    "11111111", --  599 - 0x257  :  255 - 0xff
    "00000000", --  600 - 0x258  :    0 - 0x0 -- plane 1
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x26
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "11111111", --  616 - 0x268  :  255 - 0xff -- plane 1
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11111111", --  620 - 0x26c  :  255 - 0xff
    "11111111", --  621 - 0x26d  :  255 - 0xff
    "11111111", --  622 - 0x26e  :  255 - 0xff
    "11111111", --  623 - 0x26f  :  255 - 0xff
    "11111111", --  624 - 0x270  :  255 - 0xff -- Background 0x27
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11111111", --  626 - 0x272  :  255 - 0xff
    "11111111", --  627 - 0x273  :  255 - 0xff
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111111", --  629 - 0x275  :  255 - 0xff
    "11111111", --  630 - 0x276  :  255 - 0xff
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11111111", --  632 - 0x278  :  255 - 0xff -- plane 1
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11111111", --  634 - 0x27a  :  255 - 0xff
    "11111111", --  635 - 0x27b  :  255 - 0xff
    "11111111", --  636 - 0x27c  :  255 - 0xff
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11111111", --  638 - 0x27e  :  255 - 0xff
    "11111111", --  639 - 0x27f  :  255 - 0xff
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x28
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "01111110", --  643 - 0x283  :  126 - 0x7e
    "01111110", --  644 - 0x284  :  126 - 0x7e
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x29
    "00000000", --  657 - 0x291  :    0 - 0x0
    "01000100", --  658 - 0x292  :   68 - 0x44
    "00101000", --  659 - 0x293  :   40 - 0x28
    "00010000", --  660 - 0x294  :   16 - 0x10
    "00101000", --  661 - 0x295  :   40 - 0x28
    "01000100", --  662 - 0x296  :   68 - 0x44
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- plane 1
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "11111111", --  672 - 0x2a0  :  255 - 0xff -- Background 0x2a
    "11111111", --  673 - 0x2a1  :  255 - 0xff
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111111", --  679 - 0x2a7  :  255 - 0xff
    "01111111", --  680 - 0x2a8  :  127 - 0x7f -- plane 1
    "01111111", --  681 - 0x2a9  :  127 - 0x7f
    "01111111", --  682 - 0x2aa  :  127 - 0x7f
    "01111111", --  683 - 0x2ab  :  127 - 0x7f
    "01111111", --  684 - 0x2ac  :  127 - 0x7f
    "01111111", --  685 - 0x2ad  :  127 - 0x7f
    "01111111", --  686 - 0x2ae  :  127 - 0x7f
    "01111111", --  687 - 0x2af  :  127 - 0x7f
    "00011000", --  688 - 0x2b0  :   24 - 0x18 -- Background 0x2b
    "00111100", --  689 - 0x2b1  :   60 - 0x3c
    "00111100", --  690 - 0x2b2  :   60 - 0x3c
    "00111100", --  691 - 0x2b3  :   60 - 0x3c
    "00011000", --  692 - 0x2b4  :   24 - 0x18
    "00011000", --  693 - 0x2b5  :   24 - 0x18
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00011000", --  695 - 0x2b7  :   24 - 0x18
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- plane 1
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Background 0x2c
    "01111111", --  705 - 0x2c1  :  127 - 0x7f
    "01111111", --  706 - 0x2c2  :  127 - 0x7f
    "01111111", --  707 - 0x2c3  :  127 - 0x7f
    "01111111", --  708 - 0x2c4  :  127 - 0x7f
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11100011", --  710 - 0x2c6  :  227 - 0xe3
    "11000001", --  711 - 0x2c7  :  193 - 0xc1
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- plane 1
    "10000000", --  713 - 0x2c9  :  128 - 0x80
    "10000000", --  714 - 0x2ca  :  128 - 0x80
    "10000000", --  715 - 0x2cb  :  128 - 0x80
    "10000000", --  716 - 0x2cc  :  128 - 0x80
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00011100", --  718 - 0x2ce  :   28 - 0x1c
    "00111110", --  719 - 0x2cf  :   62 - 0x3e
    "10000000", --  720 - 0x2d0  :  128 - 0x80 -- Background 0x2d
    "10000000", --  721 - 0x2d1  :  128 - 0x80
    "10000000", --  722 - 0x2d2  :  128 - 0x80
    "11000001", --  723 - 0x2d3  :  193 - 0xc1
    "11100011", --  724 - 0x2d4  :  227 - 0xe3
    "11111111", --  725 - 0x2d5  :  255 - 0xff
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "01111111", --  728 - 0x2d8  :  127 - 0x7f -- plane 1
    "01111111", --  729 - 0x2d9  :  127 - 0x7f
    "01111111", --  730 - 0x2da  :  127 - 0x7f
    "00111110", --  731 - 0x2db  :   62 - 0x3e
    "00011100", --  732 - 0x2dc  :   28 - 0x1c
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00111000", --  736 - 0x2e0  :   56 - 0x38 -- Background 0x2e
    "01111100", --  737 - 0x2e1  :  124 - 0x7c
    "01111100", --  738 - 0x2e2  :  124 - 0x7c
    "01111100", --  739 - 0x2e3  :  124 - 0x7c
    "01111100", --  740 - 0x2e4  :  124 - 0x7c
    "01111100", --  741 - 0x2e5  :  124 - 0x7c
    "00111000", --  742 - 0x2e6  :   56 - 0x38
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00001000", --  744 - 0x2e8  :    8 - 0x8 -- plane 1
    "00000100", --  745 - 0x2e9  :    4 - 0x4
    "00000100", --  746 - 0x2ea  :    4 - 0x4
    "00000100", --  747 - 0x2eb  :    4 - 0x4
    "00000100", --  748 - 0x2ec  :    4 - 0x4
    "00000100", --  749 - 0x2ed  :    4 - 0x4
    "00001000", --  750 - 0x2ee  :    8 - 0x8
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000011", --  752 - 0x2f0  :    3 - 0x3 -- Background 0x2f
    "00000110", --  753 - 0x2f1  :    6 - 0x6
    "00001100", --  754 - 0x2f2  :   12 - 0xc
    "00001100", --  755 - 0x2f3  :   12 - 0xc
    "00001000", --  756 - 0x2f4  :    8 - 0x8
    "00001000", --  757 - 0x2f5  :    8 - 0x8
    "00000100", --  758 - 0x2f6  :    4 - 0x4
    "00000011", --  759 - 0x2f7  :    3 - 0x3
    "00000011", --  760 - 0x2f8  :    3 - 0x3 -- plane 1
    "00000101", --  761 - 0x2f9  :    5 - 0x5
    "00001011", --  762 - 0x2fa  :   11 - 0xb
    "00001011", --  763 - 0x2fb  :   11 - 0xb
    "00001111", --  764 - 0x2fc  :   15 - 0xf
    "00001111", --  765 - 0x2fd  :   15 - 0xf
    "00000111", --  766 - 0x2fe  :    7 - 0x7
    "00000011", --  767 - 0x2ff  :    3 - 0x3
    "00000001", --  768 - 0x300  :    1 - 0x1 -- Background 0x30
    "00000010", --  769 - 0x301  :    2 - 0x2
    "00000100", --  770 - 0x302  :    4 - 0x4
    "00001000", --  771 - 0x303  :    8 - 0x8
    "00010000", --  772 - 0x304  :   16 - 0x10
    "00100000", --  773 - 0x305  :   32 - 0x20
    "01000000", --  774 - 0x306  :   64 - 0x40
    "10000000", --  775 - 0x307  :  128 - 0x80
    "00000001", --  776 - 0x308  :    1 - 0x1 -- plane 1
    "00000011", --  777 - 0x309  :    3 - 0x3
    "00000111", --  778 - 0x30a  :    7 - 0x7
    "00001111", --  779 - 0x30b  :   15 - 0xf
    "00011111", --  780 - 0x30c  :   31 - 0x1f
    "00111111", --  781 - 0x30d  :   63 - 0x3f
    "01111111", --  782 - 0x30e  :  127 - 0x7f
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Background 0x31
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000111", --  789 - 0x315  :    7 - 0x7
    "00111000", --  790 - 0x316  :   56 - 0x38
    "11000000", --  791 - 0x317  :  192 - 0xc0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- plane 1
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000111", --  797 - 0x31d  :    7 - 0x7
    "00111111", --  798 - 0x31e  :   63 - 0x3f
    "11111111", --  799 - 0x31f  :  255 - 0xff
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x32
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "11100000", --  805 - 0x325  :  224 - 0xe0
    "00011100", --  806 - 0x326  :   28 - 0x1c
    "00000011", --  807 - 0x327  :    3 - 0x3
    "00000000", --  808 - 0x328  :    0 - 0x0 -- plane 1
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "11100000", --  813 - 0x32d  :  224 - 0xe0
    "11111100", --  814 - 0x32e  :  252 - 0xfc
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "10000000", --  816 - 0x330  :  128 - 0x80 -- Background 0x33
    "01000000", --  817 - 0x331  :   64 - 0x40
    "00100000", --  818 - 0x332  :   32 - 0x20
    "00010000", --  819 - 0x333  :   16 - 0x10
    "00001000", --  820 - 0x334  :    8 - 0x8
    "00000100", --  821 - 0x335  :    4 - 0x4
    "00000010", --  822 - 0x336  :    2 - 0x2
    "00000001", --  823 - 0x337  :    1 - 0x1
    "10000000", --  824 - 0x338  :  128 - 0x80 -- plane 1
    "11000000", --  825 - 0x339  :  192 - 0xc0
    "11100000", --  826 - 0x33a  :  224 - 0xe0
    "11110000", --  827 - 0x33b  :  240 - 0xf0
    "11111000", --  828 - 0x33c  :  248 - 0xf8
    "11111100", --  829 - 0x33d  :  252 - 0xfc
    "11111110", --  830 - 0x33e  :  254 - 0xfe
    "11111111", --  831 - 0x33f  :  255 - 0xff
    "00000100", --  832 - 0x340  :    4 - 0x4 -- Background 0x34
    "00001110", --  833 - 0x341  :   14 - 0xe
    "00001110", --  834 - 0x342  :   14 - 0xe
    "00001110", --  835 - 0x343  :   14 - 0xe
    "01101110", --  836 - 0x344  :  110 - 0x6e
    "01100100", --  837 - 0x345  :  100 - 0x64
    "01100000", --  838 - 0x346  :   96 - 0x60
    "01100000", --  839 - 0x347  :   96 - 0x60
    "11111111", --  840 - 0x348  :  255 - 0xff -- plane 1
    "11111111", --  841 - 0x349  :  255 - 0xff
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111111", --  843 - 0x34b  :  255 - 0xff
    "11111111", --  844 - 0x34c  :  255 - 0xff
    "11111111", --  845 - 0x34d  :  255 - 0xff
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "00000111", --  848 - 0x350  :    7 - 0x7 -- Background 0x35
    "00001111", --  849 - 0x351  :   15 - 0xf
    "00011111", --  850 - 0x352  :   31 - 0x1f
    "00011111", --  851 - 0x353  :   31 - 0x1f
    "01111111", --  852 - 0x354  :  127 - 0x7f
    "11111111", --  853 - 0x355  :  255 - 0xff
    "11111111", --  854 - 0x356  :  255 - 0xff
    "01111111", --  855 - 0x357  :  127 - 0x7f
    "00000111", --  856 - 0x358  :    7 - 0x7 -- plane 1
    "00001000", --  857 - 0x359  :    8 - 0x8
    "00010000", --  858 - 0x35a  :   16 - 0x10
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "01100000", --  860 - 0x35c  :   96 - 0x60
    "10000000", --  861 - 0x35d  :  128 - 0x80
    "10000000", --  862 - 0x35e  :  128 - 0x80
    "01000000", --  863 - 0x35f  :   64 - 0x40
    "00000011", --  864 - 0x360  :    3 - 0x3 -- Background 0x36
    "00000111", --  865 - 0x361  :    7 - 0x7
    "00011111", --  866 - 0x362  :   31 - 0x1f
    "00111111", --  867 - 0x363  :   63 - 0x3f
    "00111111", --  868 - 0x364  :   63 - 0x3f
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "01111001", --  870 - 0x366  :  121 - 0x79
    "11110111", --  871 - 0x367  :  247 - 0xf7
    "00000011", --  872 - 0x368  :    3 - 0x3 -- plane 1
    "00000100", --  873 - 0x369  :    4 - 0x4
    "00011000", --  874 - 0x36a  :   24 - 0x18
    "00100000", --  875 - 0x36b  :   32 - 0x20
    "00100000", --  876 - 0x36c  :   32 - 0x20
    "00100000", --  877 - 0x36d  :   32 - 0x20
    "01000110", --  878 - 0x36e  :   70 - 0x46
    "10001000", --  879 - 0x36f  :  136 - 0x88
    "11000000", --  880 - 0x370  :  192 - 0xc0 -- Background 0x37
    "11100000", --  881 - 0x371  :  224 - 0xe0
    "11110000", --  882 - 0x372  :  240 - 0xf0
    "11110100", --  883 - 0x373  :  244 - 0xf4
    "11111110", --  884 - 0x374  :  254 - 0xfe
    "10111111", --  885 - 0x375  :  191 - 0xbf
    "11011111", --  886 - 0x376  :  223 - 0xdf
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11000000", --  888 - 0x378  :  192 - 0xc0 -- plane 1
    "00100000", --  889 - 0x379  :   32 - 0x20
    "00010000", --  890 - 0x37a  :   16 - 0x10
    "00010100", --  891 - 0x37b  :   20 - 0x14
    "00001010", --  892 - 0x37c  :   10 - 0xa
    "01000001", --  893 - 0x37d  :   65 - 0x41
    "00100001", --  894 - 0x37e  :   33 - 0x21
    "00000001", --  895 - 0x37f  :    1 - 0x1
    "10010000", --  896 - 0x380  :  144 - 0x90 -- Background 0x38
    "10111000", --  897 - 0x381  :  184 - 0xb8
    "11111000", --  898 - 0x382  :  248 - 0xf8
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111111", --  900 - 0x384  :  255 - 0xff
    "11111111", --  901 - 0x385  :  255 - 0xff
    "11111111", --  902 - 0x386  :  255 - 0xff
    "11111110", --  903 - 0x387  :  254 - 0xfe
    "10010000", --  904 - 0x388  :  144 - 0x90 -- plane 1
    "10101000", --  905 - 0x389  :  168 - 0xa8
    "01001000", --  906 - 0x38a  :   72 - 0x48
    "00001010", --  907 - 0x38b  :   10 - 0xa
    "00000101", --  908 - 0x38c  :    5 - 0x5
    "00000001", --  909 - 0x38d  :    1 - 0x1
    "00000001", --  910 - 0x38e  :    1 - 0x1
    "00000010", --  911 - 0x38f  :    2 - 0x2
    "00111011", --  912 - 0x390  :   59 - 0x3b -- Background 0x39
    "00011101", --  913 - 0x391  :   29 - 0x1d
    "00001110", --  914 - 0x392  :   14 - 0xe
    "00001111", --  915 - 0x393  :   15 - 0xf
    "00000111", --  916 - 0x394  :    7 - 0x7
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00100100", --  920 - 0x398  :   36 - 0x24 -- plane 1
    "00010010", --  921 - 0x399  :   18 - 0x12
    "00001001", --  922 - 0x39a  :    9 - 0x9
    "00001000", --  923 - 0x39b  :    8 - 0x8
    "00000111", --  924 - 0x39c  :    7 - 0x7
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "11111111", --  928 - 0x3a0  :  255 - 0xff -- Background 0x3a
    "10111111", --  929 - 0x3a1  :  191 - 0xbf
    "00011100", --  930 - 0x3a2  :   28 - 0x1c
    "11000000", --  931 - 0x3a3  :  192 - 0xc0
    "11110011", --  932 - 0x3a4  :  243 - 0xf3
    "11111111", --  933 - 0x3a5  :  255 - 0xff
    "01111110", --  934 - 0x3a6  :  126 - 0x7e
    "00011100", --  935 - 0x3a7  :   28 - 0x1c
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "01000000", --  937 - 0x3a9  :   64 - 0x40
    "11100011", --  938 - 0x3aa  :  227 - 0xe3
    "00111111", --  939 - 0x3ab  :   63 - 0x3f
    "00001100", --  940 - 0x3ac  :   12 - 0xc
    "10000001", --  941 - 0x3ad  :  129 - 0x81
    "01100010", --  942 - 0x3ae  :   98 - 0x62
    "00011100", --  943 - 0x3af  :   28 - 0x1c
    "10111111", --  944 - 0x3b0  :  191 - 0xbf -- Background 0x3b
    "01111111", --  945 - 0x3b1  :  127 - 0x7f
    "00111101", --  946 - 0x3b2  :   61 - 0x3d
    "10000011", --  947 - 0x3b3  :  131 - 0x83
    "11000111", --  948 - 0x3b4  :  199 - 0xc7
    "11111111", --  949 - 0x3b5  :  255 - 0xff
    "11111111", --  950 - 0x3b6  :  255 - 0xff
    "00111100", --  951 - 0x3b7  :   60 - 0x3c
    "01000000", --  952 - 0x3b8  :   64 - 0x40 -- plane 1
    "10000000", --  953 - 0x3b9  :  128 - 0x80
    "11000010", --  954 - 0x3ba  :  194 - 0xc2
    "01111100", --  955 - 0x3bb  :  124 - 0x7c
    "00111000", --  956 - 0x3bc  :   56 - 0x38
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "11000011", --  958 - 0x3be  :  195 - 0xc3
    "00111100", --  959 - 0x3bf  :   60 - 0x3c
    "11111100", --  960 - 0x3c0  :  252 - 0xfc -- Background 0x3c
    "11111110", --  961 - 0x3c1  :  254 - 0xfe
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111110", --  963 - 0x3c3  :  254 - 0xfe
    "11111110", --  964 - 0x3c4  :  254 - 0xfe
    "11111000", --  965 - 0x3c5  :  248 - 0xf8
    "01100000", --  966 - 0x3c6  :   96 - 0x60
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000100", --  968 - 0x3c8  :    4 - 0x4 -- plane 1
    "00000010", --  969 - 0x3c9  :    2 - 0x2
    "00000001", --  970 - 0x3ca  :    1 - 0x1
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000110", --  972 - 0x3cc  :    6 - 0x6
    "10011000", --  973 - 0x3cd  :  152 - 0x98
    "01100000", --  974 - 0x3ce  :   96 - 0x60
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "11000000", --  976 - 0x3d0  :  192 - 0xc0 -- Background 0x3d
    "00100000", --  977 - 0x3d1  :   32 - 0x20
    "00010000", --  978 - 0x3d2  :   16 - 0x10
    "00010000", --  979 - 0x3d3  :   16 - 0x10
    "00010000", --  980 - 0x3d4  :   16 - 0x10
    "00010000", --  981 - 0x3d5  :   16 - 0x10
    "00100000", --  982 - 0x3d6  :   32 - 0x20
    "11000000", --  983 - 0x3d7  :  192 - 0xc0
    "11000000", --  984 - 0x3d8  :  192 - 0xc0 -- plane 1
    "11100000", --  985 - 0x3d9  :  224 - 0xe0
    "11110000", --  986 - 0x3da  :  240 - 0xf0
    "11110000", --  987 - 0x3db  :  240 - 0xf0
    "11110000", --  988 - 0x3dc  :  240 - 0xf0
    "11110000", --  989 - 0x3dd  :  240 - 0xf0
    "11100000", --  990 - 0x3de  :  224 - 0xe0
    "11000000", --  991 - 0x3df  :  192 - 0xc0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00111111", --  996 - 0x3e4  :   63 - 0x3f
    "01111111", --  997 - 0x3e5  :  127 - 0x7f
    "11100000", --  998 - 0x3e6  :  224 - 0xe0
    "11000000", --  999 - 0x3e7  :  192 - 0xc0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00011100", -- 1006 - 0x3ee  :   28 - 0x1c
    "00111110", -- 1007 - 0x3ef  :   62 - 0x3e
    "10001000", -- 1008 - 0x3f0  :  136 - 0x88 -- Background 0x3f
    "10011100", -- 1009 - 0x3f1  :  156 - 0x9c
    "10001000", -- 1010 - 0x3f2  :  136 - 0x88
    "10000000", -- 1011 - 0x3f3  :  128 - 0x80
    "10000000", -- 1012 - 0x3f4  :  128 - 0x80
    "10000000", -- 1013 - 0x3f5  :  128 - 0x80
    "10000000", -- 1014 - 0x3f6  :  128 - 0x80
    "10000000", -- 1015 - 0x3f7  :  128 - 0x80
    "01111111", -- 1016 - 0x3f8  :  127 - 0x7f -- plane 1
    "01111111", -- 1017 - 0x3f9  :  127 - 0x7f
    "01111111", -- 1018 - 0x3fa  :  127 - 0x7f
    "00111110", -- 1019 - 0x3fb  :   62 - 0x3e
    "00011100", -- 1020 - 0x3fc  :   28 - 0x1c
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "11111110", -- 1024 - 0x400  :  254 - 0xfe -- Background 0x40
    "11111110", -- 1025 - 0x401  :  254 - 0xfe
    "11111110", -- 1026 - 0x402  :  254 - 0xfe
    "11111110", -- 1027 - 0x403  :  254 - 0xfe
    "11111110", -- 1028 - 0x404  :  254 - 0xfe
    "11111110", -- 1029 - 0x405  :  254 - 0xfe
    "11111110", -- 1030 - 0x406  :  254 - 0xfe
    "11111110", -- 1031 - 0x407  :  254 - 0xfe
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- plane 1
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11111111", -- 1035 - 0x40b  :  255 - 0xff
    "11111111", -- 1036 - 0x40c  :  255 - 0xff
    "11111111", -- 1037 - 0x40d  :  255 - 0xff
    "11111111", -- 1038 - 0x40e  :  255 - 0xff
    "11111111", -- 1039 - 0x40f  :  255 - 0xff
    "00001000", -- 1040 - 0x410  :    8 - 0x8 -- Background 0x41
    "00010100", -- 1041 - 0x411  :   20 - 0x14
    "00100100", -- 1042 - 0x412  :   36 - 0x24
    "11000100", -- 1043 - 0x413  :  196 - 0xc4
    "00000011", -- 1044 - 0x414  :    3 - 0x3
    "01000000", -- 1045 - 0x415  :   64 - 0x40
    "10100001", -- 1046 - 0x416  :  161 - 0xa1
    "00100110", -- 1047 - 0x417  :   38 - 0x26
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- plane 1
    "00001000", -- 1049 - 0x419  :    8 - 0x8
    "00011000", -- 1050 - 0x41a  :   24 - 0x18
    "00111000", -- 1051 - 0x41b  :   56 - 0x38
    "11111100", -- 1052 - 0x41c  :  252 - 0xfc
    "10111111", -- 1053 - 0x41d  :  191 - 0xbf
    "01011110", -- 1054 - 0x41e  :   94 - 0x5e
    "11011001", -- 1055 - 0x41f  :  217 - 0xd9
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Background 0x42
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "01111111", -- 1060 - 0x424  :  127 - 0x7f
    "01111111", -- 1061 - 0x425  :  127 - 0x7f
    "01111111", -- 1062 - 0x426  :  127 - 0x7f
    "01111111", -- 1063 - 0x427  :  127 - 0x7f
    "10000001", -- 1064 - 0x428  :  129 - 0x81 -- plane 1
    "10000001", -- 1065 - 0x429  :  129 - 0x81
    "10000001", -- 1066 - 0x42a  :  129 - 0x81
    "10000001", -- 1067 - 0x42b  :  129 - 0x81
    "10000001", -- 1068 - 0x42c  :  129 - 0x81
    "10000001", -- 1069 - 0x42d  :  129 - 0x81
    "10000001", -- 1070 - 0x42e  :  129 - 0x81
    "10000001", -- 1071 - 0x42f  :  129 - 0x81
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Background 0x43
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11111111", -- 1078 - 0x436  :  255 - 0xff
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "00000001", -- 1080 - 0x438  :    1 - 0x1 -- plane 1
    "00000001", -- 1081 - 0x439  :    1 - 0x1
    "00000001", -- 1082 - 0x43a  :    1 - 0x1
    "00000001", -- 1083 - 0x43b  :    1 - 0x1
    "00000001", -- 1084 - 0x43c  :    1 - 0x1
    "00000001", -- 1085 - 0x43d  :    1 - 0x1
    "00000001", -- 1086 - 0x43e  :    1 - 0x1
    "00000001", -- 1087 - 0x43f  :    1 - 0x1
    "01111111", -- 1088 - 0x440  :  127 - 0x7f -- Background 0x44
    "10000000", -- 1089 - 0x441  :  128 - 0x80
    "10000000", -- 1090 - 0x442  :  128 - 0x80
    "10011000", -- 1091 - 0x443  :  152 - 0x98
    "10011100", -- 1092 - 0x444  :  156 - 0x9c
    "10001100", -- 1093 - 0x445  :  140 - 0x8c
    "10000000", -- 1094 - 0x446  :  128 - 0x80
    "10000000", -- 1095 - 0x447  :  128 - 0x80
    "00000000", -- 1096 - 0x448  :    0 - 0x0 -- plane 1
    "01111111", -- 1097 - 0x449  :  127 - 0x7f
    "01111111", -- 1098 - 0x44a  :  127 - 0x7f
    "01100111", -- 1099 - 0x44b  :  103 - 0x67
    "01100111", -- 1100 - 0x44c  :  103 - 0x67
    "01111111", -- 1101 - 0x44d  :  127 - 0x7f
    "01111111", -- 1102 - 0x44e  :  127 - 0x7f
    "01111111", -- 1103 - 0x44f  :  127 - 0x7f
    "11111111", -- 1104 - 0x450  :  255 - 0xff -- Background 0x45
    "00000001", -- 1105 - 0x451  :    1 - 0x1
    "00000001", -- 1106 - 0x452  :    1 - 0x1
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "00010000", -- 1108 - 0x454  :   16 - 0x10
    "00010000", -- 1109 - 0x455  :   16 - 0x10
    "00010000", -- 1110 - 0x456  :   16 - 0x10
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "00000000", -- 1112 - 0x458  :    0 - 0x0 -- plane 1
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "11111111", -- 1117 - 0x45d  :  255 - 0xff
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11111111", -- 1119 - 0x45f  :  255 - 0xff
    "10000000", -- 1120 - 0x460  :  128 - 0x80 -- Background 0x46
    "10000000", -- 1121 - 0x461  :  128 - 0x80
    "10000000", -- 1122 - 0x462  :  128 - 0x80
    "10000000", -- 1123 - 0x463  :  128 - 0x80
    "10000000", -- 1124 - 0x464  :  128 - 0x80
    "10000000", -- 1125 - 0x465  :  128 - 0x80
    "10000000", -- 1126 - 0x466  :  128 - 0x80
    "10000000", -- 1127 - 0x467  :  128 - 0x80
    "01111111", -- 1128 - 0x468  :  127 - 0x7f -- plane 1
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "01111111", -- 1130 - 0x46a  :  127 - 0x7f
    "01111111", -- 1131 - 0x46b  :  127 - 0x7f
    "01111111", -- 1132 - 0x46c  :  127 - 0x7f
    "01111111", -- 1133 - 0x46d  :  127 - 0x7f
    "01111111", -- 1134 - 0x46e  :  127 - 0x7f
    "01111111", -- 1135 - 0x46f  :  127 - 0x7f
    "00000001", -- 1136 - 0x470  :    1 - 0x1 -- Background 0x47
    "00000001", -- 1137 - 0x471  :    1 - 0x1
    "00000001", -- 1138 - 0x472  :    1 - 0x1
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "00010000", -- 1140 - 0x474  :   16 - 0x10
    "00010000", -- 1141 - 0x475  :   16 - 0x10
    "00010000", -- 1142 - 0x476  :   16 - 0x10
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- plane 1
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111111", -- 1146 - 0x47a  :  255 - 0xff
    "11111111", -- 1147 - 0x47b  :  255 - 0xff
    "11111111", -- 1148 - 0x47c  :  255 - 0xff
    "11111111", -- 1149 - 0x47d  :  255 - 0xff
    "11111111", -- 1150 - 0x47e  :  255 - 0xff
    "11111111", -- 1151 - 0x47f  :  255 - 0xff
    "11111111", -- 1152 - 0x480  :  255 - 0xff -- Background 0x48
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- plane 1
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "11111111", -- 1163 - 0x48b  :  255 - 0xff
    "11111111", -- 1164 - 0x48c  :  255 - 0xff
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11111110", -- 1168 - 0x490  :  254 - 0xfe -- Background 0x49
    "00000001", -- 1169 - 0x491  :    1 - 0x1
    "00000001", -- 1170 - 0x492  :    1 - 0x1
    "00011001", -- 1171 - 0x493  :   25 - 0x19
    "00011101", -- 1172 - 0x494  :   29 - 0x1d
    "00001101", -- 1173 - 0x495  :   13 - 0xd
    "00000001", -- 1174 - 0x496  :    1 - 0x1
    "00000001", -- 1175 - 0x497  :    1 - 0x1
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- plane 1
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11100111", -- 1179 - 0x49b  :  231 - 0xe7
    "11100111", -- 1180 - 0x49c  :  231 - 0xe7
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "00000001", -- 1184 - 0x4a0  :    1 - 0x1 -- Background 0x4a
    "00000001", -- 1185 - 0x4a1  :    1 - 0x1
    "00000001", -- 1186 - 0x4a2  :    1 - 0x1
    "00000001", -- 1187 - 0x4a3  :    1 - 0x1
    "00000001", -- 1188 - 0x4a4  :    1 - 0x1
    "00000001", -- 1189 - 0x4a5  :    1 - 0x1
    "00000001", -- 1190 - 0x4a6  :    1 - 0x1
    "00000001", -- 1191 - 0x4a7  :    1 - 0x1
    "11111111", -- 1192 - 0x4a8  :  255 - 0xff -- plane 1
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "11111111", -- 1194 - 0x4aa  :  255 - 0xff
    "11111111", -- 1195 - 0x4ab  :  255 - 0xff
    "11111111", -- 1196 - 0x4ac  :  255 - 0xff
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "11111111", -- 1198 - 0x4ae  :  255 - 0xff
    "11111111", -- 1199 - 0x4af  :  255 - 0xff
    "00111111", -- 1200 - 0x4b0  :   63 - 0x3f -- Background 0x4b
    "01111111", -- 1201 - 0x4b1  :  127 - 0x7f
    "01111111", -- 1202 - 0x4b2  :  127 - 0x7f
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "11111111", -- 1204 - 0x4b4  :  255 - 0xff
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111111", -- 1206 - 0x4b6  :  255 - 0xff
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "00111111", -- 1208 - 0x4b8  :   63 - 0x3f -- plane 1
    "01100000", -- 1209 - 0x4b9  :   96 - 0x60
    "01000000", -- 1210 - 0x4ba  :   64 - 0x40
    "11000000", -- 1211 - 0x4bb  :  192 - 0xc0
    "10000000", -- 1212 - 0x4bc  :  128 - 0x80
    "10000000", -- 1213 - 0x4bd  :  128 - 0x80
    "10000000", -- 1214 - 0x4be  :  128 - 0x80
    "10000000", -- 1215 - 0x4bf  :  128 - 0x80
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x4c
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "01111110", -- 1222 - 0x4c6  :  126 - 0x7e
    "00111100", -- 1223 - 0x4c7  :   60 - 0x3c
    "10000000", -- 1224 - 0x4c8  :  128 - 0x80 -- plane 1
    "10000000", -- 1225 - 0x4c9  :  128 - 0x80
    "10000000", -- 1226 - 0x4ca  :  128 - 0x80
    "10000000", -- 1227 - 0x4cb  :  128 - 0x80
    "10000000", -- 1228 - 0x4cc  :  128 - 0x80
    "10000001", -- 1229 - 0x4cd  :  129 - 0x81
    "01000010", -- 1230 - 0x4ce  :   66 - 0x42
    "00111100", -- 1231 - 0x4cf  :   60 - 0x3c
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Background 0x4d
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11111111", -- 1235 - 0x4d3  :  255 - 0xff
    "11111111", -- 1236 - 0x4d4  :  255 - 0xff
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11111111", -- 1238 - 0x4d6  :  255 - 0xff
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- plane 1
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Background 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "11111111", -- 1250 - 0x4e2  :  255 - 0xff
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111110", -- 1254 - 0x4e6  :  254 - 0xfe
    "01111100", -- 1255 - 0x4e7  :  124 - 0x7c
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000001", -- 1261 - 0x4ed  :    1 - 0x1
    "10000010", -- 1262 - 0x4ee  :  130 - 0x82
    "01111100", -- 1263 - 0x4ef  :  124 - 0x7c
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Background 0x4f
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11111111", -- 1266 - 0x4f2  :  255 - 0xff
    "11111111", -- 1267 - 0x4f3  :  255 - 0xff
    "11111111", -- 1268 - 0x4f4  :  255 - 0xff
    "11111111", -- 1269 - 0x4f5  :  255 - 0xff
    "11111110", -- 1270 - 0x4f6  :  254 - 0xfe
    "01111100", -- 1271 - 0x4f7  :  124 - 0x7c
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000001", -- 1277 - 0x4fd  :    1 - 0x1
    "10000011", -- 1278 - 0x4fe  :  131 - 0x83
    "11111111", -- 1279 - 0x4ff  :  255 - 0xff
    "11111000", -- 1280 - 0x500  :  248 - 0xf8 -- Background 0x50
    "11111100", -- 1281 - 0x501  :  252 - 0xfc
    "11111110", -- 1282 - 0x502  :  254 - 0xfe
    "11111110", -- 1283 - 0x503  :  254 - 0xfe
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "11111000", -- 1288 - 0x508  :  248 - 0xf8 -- plane 1
    "00000100", -- 1289 - 0x509  :    4 - 0x4
    "00000010", -- 1290 - 0x50a  :    2 - 0x2
    "00000010", -- 1291 - 0x50b  :    2 - 0x2
    "00000001", -- 1292 - 0x50c  :    1 - 0x1
    "00000001", -- 1293 - 0x50d  :    1 - 0x1
    "00000001", -- 1294 - 0x50e  :    1 - 0x1
    "00000001", -- 1295 - 0x50f  :    1 - 0x1
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Background 0x51
    "11111111", -- 1297 - 0x511  :  255 - 0xff
    "11111111", -- 1298 - 0x512  :  255 - 0xff
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "11111111", -- 1300 - 0x514  :  255 - 0xff
    "11111111", -- 1301 - 0x515  :  255 - 0xff
    "01111110", -- 1302 - 0x516  :  126 - 0x7e
    "00111100", -- 1303 - 0x517  :   60 - 0x3c
    "00000001", -- 1304 - 0x518  :    1 - 0x1 -- plane 1
    "00000001", -- 1305 - 0x519  :    1 - 0x1
    "00000001", -- 1306 - 0x51a  :    1 - 0x1
    "00000001", -- 1307 - 0x51b  :    1 - 0x1
    "00000001", -- 1308 - 0x51c  :    1 - 0x1
    "10000001", -- 1309 - 0x51d  :  129 - 0x81
    "01000010", -- 1310 - 0x51e  :   66 - 0x42
    "00111100", -- 1311 - 0x51f  :   60 - 0x3c
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Background 0x52
    "00001000", -- 1313 - 0x521  :    8 - 0x8
    "00001000", -- 1314 - 0x522  :    8 - 0x8
    "00001000", -- 1315 - 0x523  :    8 - 0x8
    "00010000", -- 1316 - 0x524  :   16 - 0x10
    "00010000", -- 1317 - 0x525  :   16 - 0x10
    "00010000", -- 1318 - 0x526  :   16 - 0x10
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "11111111", -- 1320 - 0x528  :  255 - 0xff -- plane 1
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11111111", -- 1325 - 0x52d  :  255 - 0xff
    "11111111", -- 1326 - 0x52e  :  255 - 0xff
    "11111111", -- 1327 - 0x52f  :  255 - 0xff
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0x53
    "01111111", -- 1329 - 0x531  :  127 - 0x7f
    "01111111", -- 1330 - 0x532  :  127 - 0x7f
    "01111000", -- 1331 - 0x533  :  120 - 0x78
    "01110011", -- 1332 - 0x534  :  115 - 0x73
    "01110011", -- 1333 - 0x535  :  115 - 0x73
    "01110011", -- 1334 - 0x536  :  115 - 0x73
    "01111111", -- 1335 - 0x537  :  127 - 0x7f
    "01111111", -- 1336 - 0x538  :  127 - 0x7f -- plane 1
    "10000000", -- 1337 - 0x539  :  128 - 0x80
    "10100000", -- 1338 - 0x53a  :  160 - 0xa0
    "10000111", -- 1339 - 0x53b  :  135 - 0x87
    "10001111", -- 1340 - 0x53c  :  143 - 0x8f
    "10001110", -- 1341 - 0x53d  :  142 - 0x8e
    "10001110", -- 1342 - 0x53e  :  142 - 0x8e
    "10000110", -- 1343 - 0x53f  :  134 - 0x86
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Background 0x54
    "11111111", -- 1345 - 0x541  :  255 - 0xff
    "11111111", -- 1346 - 0x542  :  255 - 0xff
    "00111111", -- 1347 - 0x543  :   63 - 0x3f
    "10011111", -- 1348 - 0x544  :  159 - 0x9f
    "10011111", -- 1349 - 0x545  :  159 - 0x9f
    "10011111", -- 1350 - 0x546  :  159 - 0x9f
    "00011111", -- 1351 - 0x547  :   31 - 0x1f
    "11111110", -- 1352 - 0x548  :  254 - 0xfe -- plane 1
    "00000001", -- 1353 - 0x549  :    1 - 0x1
    "00000101", -- 1354 - 0x54a  :    5 - 0x5
    "11000001", -- 1355 - 0x54b  :  193 - 0xc1
    "11100001", -- 1356 - 0x54c  :  225 - 0xe1
    "01110001", -- 1357 - 0x54d  :  113 - 0x71
    "01110001", -- 1358 - 0x54e  :  113 - 0x71
    "11110001", -- 1359 - 0x54f  :  241 - 0xf1
    "01111110", -- 1360 - 0x550  :  126 - 0x7e -- Background 0x55
    "01111110", -- 1361 - 0x551  :  126 - 0x7e
    "01111111", -- 1362 - 0x552  :  127 - 0x7f
    "01111110", -- 1363 - 0x553  :  126 - 0x7e
    "01111110", -- 1364 - 0x554  :  126 - 0x7e
    "01111111", -- 1365 - 0x555  :  127 - 0x7f
    "01111111", -- 1366 - 0x556  :  127 - 0x7f
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "10000001", -- 1368 - 0x558  :  129 - 0x81 -- plane 1
    "10000001", -- 1369 - 0x559  :  129 - 0x81
    "10000000", -- 1370 - 0x55a  :  128 - 0x80
    "10000001", -- 1371 - 0x55b  :  129 - 0x81
    "10000001", -- 1372 - 0x55c  :  129 - 0x81
    "10100000", -- 1373 - 0x55d  :  160 - 0xa0
    "10000000", -- 1374 - 0x55e  :  128 - 0x80
    "11111111", -- 1375 - 0x55f  :  255 - 0xff
    "01111111", -- 1376 - 0x560  :  127 - 0x7f -- Background 0x56
    "01111111", -- 1377 - 0x561  :  127 - 0x7f
    "11111111", -- 1378 - 0x562  :  255 - 0xff
    "01111111", -- 1379 - 0x563  :  127 - 0x7f
    "01111111", -- 1380 - 0x564  :  127 - 0x7f
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "11111111", -- 1382 - 0x566  :  255 - 0xff
    "11111111", -- 1383 - 0x567  :  255 - 0xff
    "11110001", -- 1384 - 0x568  :  241 - 0xf1 -- plane 1
    "11000001", -- 1385 - 0x569  :  193 - 0xc1
    "11000001", -- 1386 - 0x56a  :  193 - 0xc1
    "10000001", -- 1387 - 0x56b  :  129 - 0x81
    "11000001", -- 1388 - 0x56c  :  193 - 0xc1
    "11000101", -- 1389 - 0x56d  :  197 - 0xc5
    "00000001", -- 1390 - 0x56e  :    1 - 0x1
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "01111111", -- 1392 - 0x570  :  127 - 0x7f -- Background 0x57
    "10000000", -- 1393 - 0x571  :  128 - 0x80
    "10100000", -- 1394 - 0x572  :  160 - 0xa0
    "10000000", -- 1395 - 0x573  :  128 - 0x80
    "10000000", -- 1396 - 0x574  :  128 - 0x80
    "10000000", -- 1397 - 0x575  :  128 - 0x80
    "10000000", -- 1398 - 0x576  :  128 - 0x80
    "10000000", -- 1399 - 0x577  :  128 - 0x80
    "01111111", -- 1400 - 0x578  :  127 - 0x7f -- plane 1
    "11111111", -- 1401 - 0x579  :  255 - 0xff
    "11111111", -- 1402 - 0x57a  :  255 - 0xff
    "11111111", -- 1403 - 0x57b  :  255 - 0xff
    "11111111", -- 1404 - 0x57c  :  255 - 0xff
    "11111111", -- 1405 - 0x57d  :  255 - 0xff
    "11111111", -- 1406 - 0x57e  :  255 - 0xff
    "11111111", -- 1407 - 0x57f  :  255 - 0xff
    "11111110", -- 1408 - 0x580  :  254 - 0xfe -- Background 0x58
    "00000001", -- 1409 - 0x581  :    1 - 0x1
    "00000101", -- 1410 - 0x582  :    5 - 0x5
    "00000001", -- 1411 - 0x583  :    1 - 0x1
    "00000001", -- 1412 - 0x584  :    1 - 0x1
    "00000001", -- 1413 - 0x585  :    1 - 0x1
    "00000001", -- 1414 - 0x586  :    1 - 0x1
    "00000001", -- 1415 - 0x587  :    1 - 0x1
    "11111110", -- 1416 - 0x588  :  254 - 0xfe -- plane 1
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11111111", -- 1418 - 0x58a  :  255 - 0xff
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11111111", -- 1421 - 0x58d  :  255 - 0xff
    "11111111", -- 1422 - 0x58e  :  255 - 0xff
    "11111111", -- 1423 - 0x58f  :  255 - 0xff
    "10000000", -- 1424 - 0x590  :  128 - 0x80 -- Background 0x59
    "10000000", -- 1425 - 0x591  :  128 - 0x80
    "10000000", -- 1426 - 0x592  :  128 - 0x80
    "10000000", -- 1427 - 0x593  :  128 - 0x80
    "10000000", -- 1428 - 0x594  :  128 - 0x80
    "10100000", -- 1429 - 0x595  :  160 - 0xa0
    "10000000", -- 1430 - 0x596  :  128 - 0x80
    "01111111", -- 1431 - 0x597  :  127 - 0x7f
    "11111111", -- 1432 - 0x598  :  255 - 0xff -- plane 1
    "11111111", -- 1433 - 0x599  :  255 - 0xff
    "11111111", -- 1434 - 0x59a  :  255 - 0xff
    "11111111", -- 1435 - 0x59b  :  255 - 0xff
    "11111111", -- 1436 - 0x59c  :  255 - 0xff
    "11111111", -- 1437 - 0x59d  :  255 - 0xff
    "11111111", -- 1438 - 0x59e  :  255 - 0xff
    "01111111", -- 1439 - 0x59f  :  127 - 0x7f
    "00000001", -- 1440 - 0x5a0  :    1 - 0x1 -- Background 0x5a
    "00000001", -- 1441 - 0x5a1  :    1 - 0x1
    "00000001", -- 1442 - 0x5a2  :    1 - 0x1
    "00000001", -- 1443 - 0x5a3  :    1 - 0x1
    "00000001", -- 1444 - 0x5a4  :    1 - 0x1
    "00000101", -- 1445 - 0x5a5  :    5 - 0x5
    "00000001", -- 1446 - 0x5a6  :    1 - 0x1
    "11111110", -- 1447 - 0x5a7  :  254 - 0xfe
    "11111111", -- 1448 - 0x5a8  :  255 - 0xff -- plane 1
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111111", -- 1450 - 0x5aa  :  255 - 0xff
    "11111111", -- 1451 - 0x5ab  :  255 - 0xff
    "11111111", -- 1452 - 0x5ac  :  255 - 0xff
    "11111111", -- 1453 - 0x5ad  :  255 - 0xff
    "11111111", -- 1454 - 0x5ae  :  255 - 0xff
    "11111110", -- 1455 - 0x5af  :  254 - 0xfe
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "11111100", -- 1460 - 0x5b4  :  252 - 0xfc
    "11111110", -- 1461 - 0x5b5  :  254 - 0xfe
    "00000111", -- 1462 - 0x5b6  :    7 - 0x7
    "00000011", -- 1463 - 0x5b7  :    3 - 0x3
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00111000", -- 1470 - 0x5be  :   56 - 0x38
    "01111100", -- 1471 - 0x5bf  :  124 - 0x7c
    "00010001", -- 1472 - 0x5c0  :   17 - 0x11 -- Background 0x5c
    "00111001", -- 1473 - 0x5c1  :   57 - 0x39
    "00010001", -- 1474 - 0x5c2  :   17 - 0x11
    "00000001", -- 1475 - 0x5c3  :    1 - 0x1
    "00000001", -- 1476 - 0x5c4  :    1 - 0x1
    "00000001", -- 1477 - 0x5c5  :    1 - 0x1
    "00000001", -- 1478 - 0x5c6  :    1 - 0x1
    "00000001", -- 1479 - 0x5c7  :    1 - 0x1
    "11111110", -- 1480 - 0x5c8  :  254 - 0xfe -- plane 1
    "11111110", -- 1481 - 0x5c9  :  254 - 0xfe
    "11111110", -- 1482 - 0x5ca  :  254 - 0xfe
    "01111100", -- 1483 - 0x5cb  :  124 - 0x7c
    "00111000", -- 1484 - 0x5cc  :   56 - 0x38
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "11101111", -- 1488 - 0x5d0  :  239 - 0xef -- Background 0x5d
    "00101000", -- 1489 - 0x5d1  :   40 - 0x28
    "00101000", -- 1490 - 0x5d2  :   40 - 0x28
    "00101000", -- 1491 - 0x5d3  :   40 - 0x28
    "00101000", -- 1492 - 0x5d4  :   40 - 0x28
    "00101000", -- 1493 - 0x5d5  :   40 - 0x28
    "11101111", -- 1494 - 0x5d6  :  239 - 0xef
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00100000", -- 1496 - 0x5d8  :   32 - 0x20 -- plane 1
    "11100111", -- 1497 - 0x5d9  :  231 - 0xe7
    "11100111", -- 1498 - 0x5da  :  231 - 0xe7
    "11100111", -- 1499 - 0x5db  :  231 - 0xe7
    "11100111", -- 1500 - 0x5dc  :  231 - 0xe7
    "11100111", -- 1501 - 0x5dd  :  231 - 0xe7
    "11101111", -- 1502 - 0x5de  :  239 - 0xef
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "11111110", -- 1504 - 0x5e0  :  254 - 0xfe -- Background 0x5e
    "10000010", -- 1505 - 0x5e1  :  130 - 0x82
    "10000010", -- 1506 - 0x5e2  :  130 - 0x82
    "10000010", -- 1507 - 0x5e3  :  130 - 0x82
    "10000010", -- 1508 - 0x5e4  :  130 - 0x82
    "10000010", -- 1509 - 0x5e5  :  130 - 0x82
    "11111110", -- 1510 - 0x5e6  :  254 - 0xfe
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000010", -- 1512 - 0x5e8  :    2 - 0x2 -- plane 1
    "01111110", -- 1513 - 0x5e9  :  126 - 0x7e
    "01111110", -- 1514 - 0x5ea  :  126 - 0x7e
    "01111110", -- 1515 - 0x5eb  :  126 - 0x7e
    "01111110", -- 1516 - 0x5ec  :  126 - 0x7e
    "01111110", -- 1517 - 0x5ed  :  126 - 0x7e
    "11111110", -- 1518 - 0x5ee  :  254 - 0xfe
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "10000000", -- 1520 - 0x5f0  :  128 - 0x80 -- Background 0x5f
    "10000000", -- 1521 - 0x5f1  :  128 - 0x80
    "10000000", -- 1522 - 0x5f2  :  128 - 0x80
    "10011000", -- 1523 - 0x5f3  :  152 - 0x98
    "10011100", -- 1524 - 0x5f4  :  156 - 0x9c
    "10001100", -- 1525 - 0x5f5  :  140 - 0x8c
    "10000000", -- 1526 - 0x5f6  :  128 - 0x80
    "01111111", -- 1527 - 0x5f7  :  127 - 0x7f
    "01111111", -- 1528 - 0x5f8  :  127 - 0x7f -- plane 1
    "01111111", -- 1529 - 0x5f9  :  127 - 0x7f
    "01111111", -- 1530 - 0x5fa  :  127 - 0x7f
    "01100111", -- 1531 - 0x5fb  :  103 - 0x67
    "01100111", -- 1532 - 0x5fc  :  103 - 0x67
    "01111111", -- 1533 - 0x5fd  :  127 - 0x7f
    "01111111", -- 1534 - 0x5fe  :  127 - 0x7f
    "01111111", -- 1535 - 0x5ff  :  127 - 0x7f
    "11111111", -- 1536 - 0x600  :  255 - 0xff -- Background 0x60
    "11111111", -- 1537 - 0x601  :  255 - 0xff
    "10000011", -- 1538 - 0x602  :  131 - 0x83
    "11110011", -- 1539 - 0x603  :  243 - 0xf3
    "11110011", -- 1540 - 0x604  :  243 - 0xf3
    "11110011", -- 1541 - 0x605  :  243 - 0xf3
    "11110011", -- 1542 - 0x606  :  243 - 0xf3
    "11110011", -- 1543 - 0x607  :  243 - 0xf3
    "11111111", -- 1544 - 0x608  :  255 - 0xff -- plane 1
    "10000000", -- 1545 - 0x609  :  128 - 0x80
    "11111100", -- 1546 - 0x60a  :  252 - 0xfc
    "10001100", -- 1547 - 0x60b  :  140 - 0x8c
    "10001100", -- 1548 - 0x60c  :  140 - 0x8c
    "10001100", -- 1549 - 0x60d  :  140 - 0x8c
    "10001100", -- 1550 - 0x60e  :  140 - 0x8c
    "10001100", -- 1551 - 0x60f  :  140 - 0x8c
    "11111111", -- 1552 - 0x610  :  255 - 0xff -- Background 0x61
    "11111111", -- 1553 - 0x611  :  255 - 0xff
    "11110000", -- 1554 - 0x612  :  240 - 0xf0
    "11110110", -- 1555 - 0x613  :  246 - 0xf6
    "11110110", -- 1556 - 0x614  :  246 - 0xf6
    "11110110", -- 1557 - 0x615  :  246 - 0xf6
    "11110110", -- 1558 - 0x616  :  246 - 0xf6
    "11110110", -- 1559 - 0x617  :  246 - 0xf6
    "11111111", -- 1560 - 0x618  :  255 - 0xff -- plane 1
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00001111", -- 1562 - 0x61a  :   15 - 0xf
    "00001001", -- 1563 - 0x61b  :    9 - 0x9
    "00001001", -- 1564 - 0x61c  :    9 - 0x9
    "00001001", -- 1565 - 0x61d  :    9 - 0x9
    "00001001", -- 1566 - 0x61e  :    9 - 0x9
    "00001001", -- 1567 - 0x61f  :    9 - 0x9
    "11111111", -- 1568 - 0x620  :  255 - 0xff -- Background 0x62
    "11111111", -- 1569 - 0x621  :  255 - 0xff
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "11111111", -- 1576 - 0x628  :  255 - 0xff -- plane 1
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "11111111", -- 1578 - 0x62a  :  255 - 0xff
    "11111111", -- 1579 - 0x62b  :  255 - 0xff
    "11111111", -- 1580 - 0x62c  :  255 - 0xff
    "11111111", -- 1581 - 0x62d  :  255 - 0xff
    "11111111", -- 1582 - 0x62e  :  255 - 0xff
    "11111111", -- 1583 - 0x62f  :  255 - 0xff
    "11111111", -- 1584 - 0x630  :  255 - 0xff -- Background 0x63
    "11111111", -- 1585 - 0x631  :  255 - 0xff
    "00000001", -- 1586 - 0x632  :    1 - 0x1
    "01010111", -- 1587 - 0x633  :   87 - 0x57
    "00101111", -- 1588 - 0x634  :   47 - 0x2f
    "01010111", -- 1589 - 0x635  :   87 - 0x57
    "00101111", -- 1590 - 0x636  :   47 - 0x2f
    "01010111", -- 1591 - 0x637  :   87 - 0x57
    "11111111", -- 1592 - 0x638  :  255 - 0xff -- plane 1
    "00000001", -- 1593 - 0x639  :    1 - 0x1
    "11111111", -- 1594 - 0x63a  :  255 - 0xff
    "10101001", -- 1595 - 0x63b  :  169 - 0xa9
    "11010001", -- 1596 - 0x63c  :  209 - 0xd1
    "10101001", -- 1597 - 0x63d  :  169 - 0xa9
    "11010001", -- 1598 - 0x63e  :  209 - 0xd1
    "10101001", -- 1599 - 0x63f  :  169 - 0xa9
    "11110011", -- 1600 - 0x640  :  243 - 0xf3 -- Background 0x64
    "11110011", -- 1601 - 0x641  :  243 - 0xf3
    "11110011", -- 1602 - 0x642  :  243 - 0xf3
    "11110011", -- 1603 - 0x643  :  243 - 0xf3
    "11110011", -- 1604 - 0x644  :  243 - 0xf3
    "11110011", -- 1605 - 0x645  :  243 - 0xf3
    "11111111", -- 1606 - 0x646  :  255 - 0xff
    "00111111", -- 1607 - 0x647  :   63 - 0x3f
    "10001100", -- 1608 - 0x648  :  140 - 0x8c -- plane 1
    "10001100", -- 1609 - 0x649  :  140 - 0x8c
    "10001100", -- 1610 - 0x64a  :  140 - 0x8c
    "10001100", -- 1611 - 0x64b  :  140 - 0x8c
    "10001100", -- 1612 - 0x64c  :  140 - 0x8c
    "10001100", -- 1613 - 0x64d  :  140 - 0x8c
    "11111111", -- 1614 - 0x64e  :  255 - 0xff
    "00111111", -- 1615 - 0x64f  :   63 - 0x3f
    "11110110", -- 1616 - 0x650  :  246 - 0xf6 -- Background 0x65
    "11110110", -- 1617 - 0x651  :  246 - 0xf6
    "11110110", -- 1618 - 0x652  :  246 - 0xf6
    "11110110", -- 1619 - 0x653  :  246 - 0xf6
    "11110110", -- 1620 - 0x654  :  246 - 0xf6
    "11110110", -- 1621 - 0x655  :  246 - 0xf6
    "11111111", -- 1622 - 0x656  :  255 - 0xff
    "11111111", -- 1623 - 0x657  :  255 - 0xff
    "00001001", -- 1624 - 0x658  :    9 - 0x9 -- plane 1
    "00001001", -- 1625 - 0x659  :    9 - 0x9
    "00001001", -- 1626 - 0x65a  :    9 - 0x9
    "00001001", -- 1627 - 0x65b  :    9 - 0x9
    "00001001", -- 1628 - 0x65c  :    9 - 0x9
    "00001001", -- 1629 - 0x65d  :    9 - 0x9
    "11111111", -- 1630 - 0x65e  :  255 - 0xff
    "11111111", -- 1631 - 0x65f  :  255 - 0xff
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Background 0x66
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "11111111", -- 1639 - 0x667  :  255 - 0xff
    "11111111", -- 1640 - 0x668  :  255 - 0xff -- plane 1
    "11111111", -- 1641 - 0x669  :  255 - 0xff
    "11111111", -- 1642 - 0x66a  :  255 - 0xff
    "11111111", -- 1643 - 0x66b  :  255 - 0xff
    "11111111", -- 1644 - 0x66c  :  255 - 0xff
    "11111111", -- 1645 - 0x66d  :  255 - 0xff
    "11111111", -- 1646 - 0x66e  :  255 - 0xff
    "11111111", -- 1647 - 0x66f  :  255 - 0xff
    "00101111", -- 1648 - 0x670  :   47 - 0x2f -- Background 0x67
    "01010111", -- 1649 - 0x671  :   87 - 0x57
    "00101111", -- 1650 - 0x672  :   47 - 0x2f
    "01010111", -- 1651 - 0x673  :   87 - 0x57
    "00101111", -- 1652 - 0x674  :   47 - 0x2f
    "01010111", -- 1653 - 0x675  :   87 - 0x57
    "11111111", -- 1654 - 0x676  :  255 - 0xff
    "11111100", -- 1655 - 0x677  :  252 - 0xfc
    "11010001", -- 1656 - 0x678  :  209 - 0xd1 -- plane 1
    "10101001", -- 1657 - 0x679  :  169 - 0xa9
    "11010001", -- 1658 - 0x67a  :  209 - 0xd1
    "10101001", -- 1659 - 0x67b  :  169 - 0xa9
    "11010001", -- 1660 - 0x67c  :  209 - 0xd1
    "10101001", -- 1661 - 0x67d  :  169 - 0xa9
    "11111111", -- 1662 - 0x67e  :  255 - 0xff
    "11111100", -- 1663 - 0x67f  :  252 - 0xfc
    "00111100", -- 1664 - 0x680  :   60 - 0x3c -- Background 0x68
    "00111100", -- 1665 - 0x681  :   60 - 0x3c
    "00111100", -- 1666 - 0x682  :   60 - 0x3c
    "00111100", -- 1667 - 0x683  :   60 - 0x3c
    "00111100", -- 1668 - 0x684  :   60 - 0x3c
    "00111100", -- 1669 - 0x685  :   60 - 0x3c
    "00111100", -- 1670 - 0x686  :   60 - 0x3c
    "00111100", -- 1671 - 0x687  :   60 - 0x3c
    "00100011", -- 1672 - 0x688  :   35 - 0x23 -- plane 1
    "00100011", -- 1673 - 0x689  :   35 - 0x23
    "00100011", -- 1674 - 0x68a  :   35 - 0x23
    "00100011", -- 1675 - 0x68b  :   35 - 0x23
    "00100011", -- 1676 - 0x68c  :   35 - 0x23
    "00100011", -- 1677 - 0x68d  :   35 - 0x23
    "00100011", -- 1678 - 0x68e  :   35 - 0x23
    "00100011", -- 1679 - 0x68f  :   35 - 0x23
    "11111011", -- 1680 - 0x690  :  251 - 0xfb -- Background 0x69
    "11111011", -- 1681 - 0x691  :  251 - 0xfb
    "11111011", -- 1682 - 0x692  :  251 - 0xfb
    "11111011", -- 1683 - 0x693  :  251 - 0xfb
    "11111011", -- 1684 - 0x694  :  251 - 0xfb
    "11111011", -- 1685 - 0x695  :  251 - 0xfb
    "11111011", -- 1686 - 0x696  :  251 - 0xfb
    "11111011", -- 1687 - 0x697  :  251 - 0xfb
    "00000100", -- 1688 - 0x698  :    4 - 0x4 -- plane 1
    "00000100", -- 1689 - 0x699  :    4 - 0x4
    "00000100", -- 1690 - 0x69a  :    4 - 0x4
    "00000100", -- 1691 - 0x69b  :    4 - 0x4
    "00000100", -- 1692 - 0x69c  :    4 - 0x4
    "00000100", -- 1693 - 0x69d  :    4 - 0x4
    "00000100", -- 1694 - 0x69e  :    4 - 0x4
    "00000100", -- 1695 - 0x69f  :    4 - 0x4
    "10111100", -- 1696 - 0x6a0  :  188 - 0xbc -- Background 0x6a
    "01011100", -- 1697 - 0x6a1  :   92 - 0x5c
    "10111100", -- 1698 - 0x6a2  :  188 - 0xbc
    "01011100", -- 1699 - 0x6a3  :   92 - 0x5c
    "10111100", -- 1700 - 0x6a4  :  188 - 0xbc
    "01011100", -- 1701 - 0x6a5  :   92 - 0x5c
    "10111100", -- 1702 - 0x6a6  :  188 - 0xbc
    "01011100", -- 1703 - 0x6a7  :   92 - 0x5c
    "01000100", -- 1704 - 0x6a8  :   68 - 0x44 -- plane 1
    "10100100", -- 1705 - 0x6a9  :  164 - 0xa4
    "01000100", -- 1706 - 0x6aa  :   68 - 0x44
    "10100100", -- 1707 - 0x6ab  :  164 - 0xa4
    "01000100", -- 1708 - 0x6ac  :   68 - 0x44
    "10100100", -- 1709 - 0x6ad  :  164 - 0xa4
    "01000100", -- 1710 - 0x6ae  :   68 - 0x44
    "10100100", -- 1711 - 0x6af  :  164 - 0xa4
    "00011111", -- 1712 - 0x6b0  :   31 - 0x1f -- Background 0x6b
    "00100000", -- 1713 - 0x6b1  :   32 - 0x20
    "01000000", -- 1714 - 0x6b2  :   64 - 0x40
    "01000000", -- 1715 - 0x6b3  :   64 - 0x40
    "10000000", -- 1716 - 0x6b4  :  128 - 0x80
    "10000000", -- 1717 - 0x6b5  :  128 - 0x80
    "10000000", -- 1718 - 0x6b6  :  128 - 0x80
    "10000001", -- 1719 - 0x6b7  :  129 - 0x81
    "00011111", -- 1720 - 0x6b8  :   31 - 0x1f -- plane 1
    "00111111", -- 1721 - 0x6b9  :   63 - 0x3f
    "01111111", -- 1722 - 0x6ba  :  127 - 0x7f
    "01111111", -- 1723 - 0x6bb  :  127 - 0x7f
    "11111111", -- 1724 - 0x6bc  :  255 - 0xff
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111110", -- 1727 - 0x6bf  :  254 - 0xfe
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Background 0x6c
    "10000000", -- 1729 - 0x6c1  :  128 - 0x80
    "10000000", -- 1730 - 0x6c2  :  128 - 0x80
    "11000000", -- 1731 - 0x6c3  :  192 - 0xc0
    "11111111", -- 1732 - 0x6c4  :  255 - 0xff
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111110", -- 1734 - 0x6c6  :  254 - 0xfe
    "11111110", -- 1735 - 0x6c7  :  254 - 0xfe
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- plane 1
    "01111111", -- 1737 - 0x6c9  :  127 - 0x7f
    "01111111", -- 1738 - 0x6ca  :  127 - 0x7f
    "00111111", -- 1739 - 0x6cb  :   63 - 0x3f
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000001", -- 1742 - 0x6ce  :    1 - 0x1
    "00000001", -- 1743 - 0x6cf  :    1 - 0x1
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Background 0x6d
    "01111111", -- 1745 - 0x6d1  :  127 - 0x7f
    "01111111", -- 1746 - 0x6d2  :  127 - 0x7f
    "11111111", -- 1747 - 0x6d3  :  255 - 0xff
    "11111111", -- 1748 - 0x6d4  :  255 - 0xff
    "00000111", -- 1749 - 0x6d5  :    7 - 0x7
    "00000011", -- 1750 - 0x6d6  :    3 - 0x3
    "00000011", -- 1751 - 0x6d7  :    3 - 0x3
    "11111111", -- 1752 - 0x6d8  :  255 - 0xff -- plane 1
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "10000000", -- 1754 - 0x6da  :  128 - 0x80
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "11111000", -- 1757 - 0x6dd  :  248 - 0xf8
    "11111100", -- 1758 - 0x6de  :  252 - 0xfc
    "11111100", -- 1759 - 0x6df  :  252 - 0xfc
    "11111111", -- 1760 - 0x6e0  :  255 - 0xff -- Background 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "10000001", -- 1765 - 0x6e5  :  129 - 0x81
    "11000011", -- 1766 - 0x6e6  :  195 - 0xc3
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "11111111", -- 1768 - 0x6e8  :  255 - 0xff -- plane 1
    "11111111", -- 1769 - 0x6e9  :  255 - 0xff
    "11111111", -- 1770 - 0x6ea  :  255 - 0xff
    "11111111", -- 1771 - 0x6eb  :  255 - 0xff
    "11111111", -- 1772 - 0x6ec  :  255 - 0xff
    "01111110", -- 1773 - 0x6ed  :  126 - 0x7e
    "00111100", -- 1774 - 0x6ee  :   60 - 0x3c
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11111000", -- 1776 - 0x6f0  :  248 - 0xf8 -- Background 0x6f
    "11111100", -- 1777 - 0x6f1  :  252 - 0xfc
    "11111110", -- 1778 - 0x6f2  :  254 - 0xfe
    "11111110", -- 1779 - 0x6f3  :  254 - 0xfe
    "11100011", -- 1780 - 0x6f4  :  227 - 0xe3
    "11000001", -- 1781 - 0x6f5  :  193 - 0xc1
    "10000001", -- 1782 - 0x6f6  :  129 - 0x81
    "10000001", -- 1783 - 0x6f7  :  129 - 0x81
    "11111000", -- 1784 - 0x6f8  :  248 - 0xf8 -- plane 1
    "00000100", -- 1785 - 0x6f9  :    4 - 0x4
    "00000010", -- 1786 - 0x6fa  :    2 - 0x2
    "00000010", -- 1787 - 0x6fb  :    2 - 0x2
    "00011101", -- 1788 - 0x6fc  :   29 - 0x1d
    "00111111", -- 1789 - 0x6fd  :   63 - 0x3f
    "01111111", -- 1790 - 0x6fe  :  127 - 0x7f
    "01111111", -- 1791 - 0x6ff  :  127 - 0x7f
    "10000011", -- 1792 - 0x700  :  131 - 0x83 -- Background 0x70
    "11111111", -- 1793 - 0x701  :  255 - 0xff
    "11111111", -- 1794 - 0x702  :  255 - 0xff
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "11111111", -- 1796 - 0x704  :  255 - 0xff
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "01111111", -- 1798 - 0x706  :  127 - 0x7f
    "00011111", -- 1799 - 0x707  :   31 - 0x1f
    "11111100", -- 1800 - 0x708  :  252 - 0xfc -- plane 1
    "10000000", -- 1801 - 0x709  :  128 - 0x80
    "10000000", -- 1802 - 0x70a  :  128 - 0x80
    "10000000", -- 1803 - 0x70b  :  128 - 0x80
    "10000000", -- 1804 - 0x70c  :  128 - 0x80
    "10000000", -- 1805 - 0x70d  :  128 - 0x80
    "01100000", -- 1806 - 0x70e  :   96 - 0x60
    "00011111", -- 1807 - 0x70f  :   31 - 0x1f
    "11111100", -- 1808 - 0x710  :  252 - 0xfc -- Background 0x71
    "11111100", -- 1809 - 0x711  :  252 - 0xfc
    "11111100", -- 1810 - 0x712  :  252 - 0xfc
    "11111100", -- 1811 - 0x713  :  252 - 0xfc
    "11111110", -- 1812 - 0x714  :  254 - 0xfe
    "11111110", -- 1813 - 0x715  :  254 - 0xfe
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "00000011", -- 1816 - 0x718  :    3 - 0x3 -- plane 1
    "00000011", -- 1817 - 0x719  :    3 - 0x3
    "00000011", -- 1818 - 0x71a  :    3 - 0x3
    "00000011", -- 1819 - 0x71b  :    3 - 0x3
    "00000001", -- 1820 - 0x71c  :    1 - 0x1
    "00000001", -- 1821 - 0x71d  :    1 - 0x1
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "00000001", -- 1824 - 0x720  :    1 - 0x1 -- Background 0x72
    "00000001", -- 1825 - 0x721  :    1 - 0x1
    "00000001", -- 1826 - 0x722  :    1 - 0x1
    "00000001", -- 1827 - 0x723  :    1 - 0x1
    "00000011", -- 1828 - 0x724  :    3 - 0x3
    "00000011", -- 1829 - 0x725  :    3 - 0x3
    "00000111", -- 1830 - 0x726  :    7 - 0x7
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111110", -- 1832 - 0x728  :  254 - 0xfe -- plane 1
    "11111110", -- 1833 - 0x729  :  254 - 0xfe
    "11111110", -- 1834 - 0x72a  :  254 - 0xfe
    "11111110", -- 1835 - 0x72b  :  254 - 0xfe
    "11111100", -- 1836 - 0x72c  :  252 - 0xfc
    "11111100", -- 1837 - 0x72d  :  252 - 0xfc
    "11111000", -- 1838 - 0x72e  :  248 - 0xf8
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Background 0x73
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11111111", -- 1843 - 0x733  :  255 - 0xff
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11111111", -- 1845 - 0x735  :  255 - 0xff
    "11111111", -- 1846 - 0x736  :  255 - 0xff
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- plane 1
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "10000001", -- 1856 - 0x740  :  129 - 0x81 -- Background 0x74
    "11000001", -- 1857 - 0x741  :  193 - 0xc1
    "11100011", -- 1858 - 0x742  :  227 - 0xe3
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111110", -- 1863 - 0x747  :  254 - 0xfe
    "01111111", -- 1864 - 0x748  :  127 - 0x7f -- plane 1
    "00111111", -- 1865 - 0x749  :   63 - 0x3f
    "00011101", -- 1866 - 0x74a  :   29 - 0x1d
    "00000001", -- 1867 - 0x74b  :    1 - 0x1
    "00000001", -- 1868 - 0x74c  :    1 - 0x1
    "00000001", -- 1869 - 0x74d  :    1 - 0x1
    "00000011", -- 1870 - 0x74e  :    3 - 0x3
    "11111110", -- 1871 - 0x74f  :  254 - 0xfe
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Background 0x75
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111011", -- 1877 - 0x755  :  251 - 0xfb
    "10110101", -- 1878 - 0x756  :  181 - 0xb5
    "11001110", -- 1879 - 0x757  :  206 - 0xce
    "10000000", -- 1880 - 0x758  :  128 - 0x80 -- plane 1
    "10000000", -- 1881 - 0x759  :  128 - 0x80
    "10000000", -- 1882 - 0x75a  :  128 - 0x80
    "10000000", -- 1883 - 0x75b  :  128 - 0x80
    "10000000", -- 1884 - 0x75c  :  128 - 0x80
    "10000100", -- 1885 - 0x75d  :  132 - 0x84
    "11001010", -- 1886 - 0x75e  :  202 - 0xca
    "10110001", -- 1887 - 0x75f  :  177 - 0xb1
    "11111111", -- 1888 - 0x760  :  255 - 0xff -- Background 0x76
    "11111111", -- 1889 - 0x761  :  255 - 0xff
    "11111111", -- 1890 - 0x762  :  255 - 0xff
    "11111111", -- 1891 - 0x763  :  255 - 0xff
    "11111111", -- 1892 - 0x764  :  255 - 0xff
    "11011111", -- 1893 - 0x765  :  223 - 0xdf
    "10101101", -- 1894 - 0x766  :  173 - 0xad
    "01110011", -- 1895 - 0x767  :  115 - 0x73
    "00000001", -- 1896 - 0x768  :    1 - 0x1 -- plane 1
    "00000001", -- 1897 - 0x769  :    1 - 0x1
    "00000001", -- 1898 - 0x76a  :    1 - 0x1
    "00000001", -- 1899 - 0x76b  :    1 - 0x1
    "00000001", -- 1900 - 0x76c  :    1 - 0x1
    "00100001", -- 1901 - 0x76d  :   33 - 0x21
    "01010011", -- 1902 - 0x76e  :   83 - 0x53
    "10001101", -- 1903 - 0x76f  :  141 - 0x8d
    "01110111", -- 1904 - 0x770  :  119 - 0x77 -- Background 0x77
    "01110111", -- 1905 - 0x771  :  119 - 0x77
    "01110111", -- 1906 - 0x772  :  119 - 0x77
    "01110111", -- 1907 - 0x773  :  119 - 0x77
    "01110111", -- 1908 - 0x774  :  119 - 0x77
    "01110111", -- 1909 - 0x775  :  119 - 0x77
    "01110111", -- 1910 - 0x776  :  119 - 0x77
    "01110111", -- 1911 - 0x777  :  119 - 0x77
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- plane 1
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "01110111", -- 1916 - 0x77c  :  119 - 0x77
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11111111", -- 1919 - 0x77f  :  255 - 0xff
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- plane 1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "01110111", -- 1936 - 0x790  :  119 - 0x77 -- Background 0x79
    "01110111", -- 1937 - 0x791  :  119 - 0x77
    "01110111", -- 1938 - 0x792  :  119 - 0x77
    "01110111", -- 1939 - 0x793  :  119 - 0x77
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- plane 1
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "01110111", -- 1947 - 0x79b  :  119 - 0x77
    "01110111", -- 1948 - 0x79c  :  119 - 0x77
    "01110111", -- 1949 - 0x79d  :  119 - 0x77
    "01110111", -- 1950 - 0x79e  :  119 - 0x77
    "01110111", -- 1951 - 0x79f  :  119 - 0x77
    "00000001", -- 1952 - 0x7a0  :    1 - 0x1 -- Background 0x7a
    "00000001", -- 1953 - 0x7a1  :    1 - 0x1
    "00000001", -- 1954 - 0x7a2  :    1 - 0x1
    "00011001", -- 1955 - 0x7a3  :   25 - 0x19
    "00011101", -- 1956 - 0x7a4  :   29 - 0x1d
    "00001101", -- 1957 - 0x7a5  :   13 - 0xd
    "00000001", -- 1958 - 0x7a6  :    1 - 0x1
    "11111110", -- 1959 - 0x7a7  :  254 - 0xfe
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- plane 1
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11100111", -- 1963 - 0x7ab  :  231 - 0xe7
    "11100111", -- 1964 - 0x7ac  :  231 - 0xe7
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111110", -- 1967 - 0x7af  :  254 - 0xfe
    "00100000", -- 1968 - 0x7b0  :   32 - 0x20 -- Background 0x7b
    "01111000", -- 1969 - 0x7b1  :  120 - 0x78
    "01111111", -- 1970 - 0x7b2  :  127 - 0x7f
    "11111110", -- 1971 - 0x7b3  :  254 - 0xfe
    "11111110", -- 1972 - 0x7b4  :  254 - 0xfe
    "11111110", -- 1973 - 0x7b5  :  254 - 0xfe
    "11111110", -- 1974 - 0x7b6  :  254 - 0xfe
    "11111110", -- 1975 - 0x7b7  :  254 - 0xfe
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- plane 1
    "00100001", -- 1977 - 0x7b9  :   33 - 0x21
    "00100001", -- 1978 - 0x7ba  :   33 - 0x21
    "01000001", -- 1979 - 0x7bb  :   65 - 0x41
    "01000001", -- 1980 - 0x7bc  :   65 - 0x41
    "01000001", -- 1981 - 0x7bd  :   65 - 0x41
    "01000001", -- 1982 - 0x7be  :   65 - 0x41
    "01000001", -- 1983 - 0x7bf  :   65 - 0x41
    "00000100", -- 1984 - 0x7c0  :    4 - 0x4 -- Background 0x7c
    "10011010", -- 1985 - 0x7c1  :  154 - 0x9a
    "11111010", -- 1986 - 0x7c2  :  250 - 0xfa
    "11111101", -- 1987 - 0x7c3  :  253 - 0xfd
    "11111101", -- 1988 - 0x7c4  :  253 - 0xfd
    "11111101", -- 1989 - 0x7c5  :  253 - 0xfd
    "11111101", -- 1990 - 0x7c6  :  253 - 0xfd
    "11111101", -- 1991 - 0x7c7  :  253 - 0xfd
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "10000000", -- 1993 - 0x7c9  :  128 - 0x80
    "10000000", -- 1994 - 0x7ca  :  128 - 0x80
    "10000000", -- 1995 - 0x7cb  :  128 - 0x80
    "10000000", -- 1996 - 0x7cc  :  128 - 0x80
    "10000000", -- 1997 - 0x7cd  :  128 - 0x80
    "10000000", -- 1998 - 0x7ce  :  128 - 0x80
    "10000000", -- 1999 - 0x7cf  :  128 - 0x80
    "01111110", -- 2000 - 0x7d0  :  126 - 0x7e -- Background 0x7d
    "00111000", -- 2001 - 0x7d1  :   56 - 0x38
    "00100001", -- 2002 - 0x7d2  :   33 - 0x21
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000001", -- 2004 - 0x7d4  :    1 - 0x1
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000001", -- 2006 - 0x7d6  :    1 - 0x1
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00100001", -- 2008 - 0x7d8  :   33 - 0x21 -- plane 1
    "00100001", -- 2009 - 0x7d9  :   33 - 0x21
    "00000001", -- 2010 - 0x7da  :    1 - 0x1
    "00000001", -- 2011 - 0x7db  :    1 - 0x1
    "00000001", -- 2012 - 0x7dc  :    1 - 0x1
    "00000001", -- 2013 - 0x7dd  :    1 - 0x1
    "00000001", -- 2014 - 0x7de  :    1 - 0x1
    "00000001", -- 2015 - 0x7df  :    1 - 0x1
    "11111010", -- 2016 - 0x7e0  :  250 - 0xfa -- Background 0x7e
    "10001010", -- 2017 - 0x7e1  :  138 - 0x8a
    "10000100", -- 2018 - 0x7e2  :  132 - 0x84
    "10000000", -- 2019 - 0x7e3  :  128 - 0x80
    "10000000", -- 2020 - 0x7e4  :  128 - 0x80
    "10000000", -- 2021 - 0x7e5  :  128 - 0x80
    "10000000", -- 2022 - 0x7e6  :  128 - 0x80
    "10000000", -- 2023 - 0x7e7  :  128 - 0x80
    "10000000", -- 2024 - 0x7e8  :  128 - 0x80 -- plane 1
    "10000000", -- 2025 - 0x7e9  :  128 - 0x80
    "10000000", -- 2026 - 0x7ea  :  128 - 0x80
    "10000000", -- 2027 - 0x7eb  :  128 - 0x80
    "10000000", -- 2028 - 0x7ec  :  128 - 0x80
    "10000000", -- 2029 - 0x7ed  :  128 - 0x80
    "10000000", -- 2030 - 0x7ee  :  128 - 0x80
    "10000000", -- 2031 - 0x7ef  :  128 - 0x80
    "00000010", -- 2032 - 0x7f0  :    2 - 0x2 -- Background 0x7f
    "00000100", -- 2033 - 0x7f1  :    4 - 0x4
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00010000", -- 2035 - 0x7f3  :   16 - 0x10
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "01000000", -- 2037 - 0x7f5  :   64 - 0x40
    "10000000", -- 2038 - 0x7f6  :  128 - 0x80
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000001", -- 2040 - 0x7f8  :    1 - 0x1 -- plane 1
    "00000001", -- 2041 - 0x7f9  :    1 - 0x1
    "00000110", -- 2042 - 0x7fa  :    6 - 0x6
    "00001000", -- 2043 - 0x7fb  :    8 - 0x8
    "00011000", -- 2044 - 0x7fc  :   24 - 0x18
    "00100000", -- 2045 - 0x7fd  :   32 - 0x20
    "00100000", -- 2046 - 0x7fe  :   32 - 0x20
    "11000000", -- 2047 - 0x7ff  :  192 - 0xc0
    "00001011", -- 2048 - 0x800  :   11 - 0xb -- Background 0x80
    "00001011", -- 2049 - 0x801  :   11 - 0xb
    "00111011", -- 2050 - 0x802  :   59 - 0x3b
    "00001011", -- 2051 - 0x803  :   11 - 0xb
    "11111011", -- 2052 - 0x804  :  251 - 0xfb
    "00001011", -- 2053 - 0x805  :   11 - 0xb
    "00001011", -- 2054 - 0x806  :   11 - 0xb
    "00001010", -- 2055 - 0x807  :   10 - 0xa
    "00000100", -- 2056 - 0x808  :    4 - 0x4 -- plane 1
    "00000100", -- 2057 - 0x809  :    4 - 0x4
    "11000100", -- 2058 - 0x80a  :  196 - 0xc4
    "11110100", -- 2059 - 0x80b  :  244 - 0xf4
    "11110100", -- 2060 - 0x80c  :  244 - 0xf4
    "00000100", -- 2061 - 0x80d  :    4 - 0x4
    "00000100", -- 2062 - 0x80e  :    4 - 0x4
    "00000101", -- 2063 - 0x80f  :    5 - 0x5
    "10010000", -- 2064 - 0x810  :  144 - 0x90 -- Background 0x81
    "00010000", -- 2065 - 0x811  :   16 - 0x10
    "00011111", -- 2066 - 0x812  :   31 - 0x1f
    "00010000", -- 2067 - 0x813  :   16 - 0x10
    "00011111", -- 2068 - 0x814  :   31 - 0x1f
    "00010000", -- 2069 - 0x815  :   16 - 0x10
    "00010000", -- 2070 - 0x816  :   16 - 0x10
    "10010000", -- 2071 - 0x817  :  144 - 0x90
    "01110000", -- 2072 - 0x818  :  112 - 0x70 -- plane 1
    "11110000", -- 2073 - 0x819  :  240 - 0xf0
    "11110000", -- 2074 - 0x81a  :  240 - 0xf0
    "11111111", -- 2075 - 0x81b  :  255 - 0xff
    "11111111", -- 2076 - 0x81c  :  255 - 0xff
    "11110000", -- 2077 - 0x81d  :  240 - 0xf0
    "11110000", -- 2078 - 0x81e  :  240 - 0xf0
    "01110000", -- 2079 - 0x81f  :  112 - 0x70
    "00111111", -- 2080 - 0x820  :   63 - 0x3f -- Background 0x82
    "01111000", -- 2081 - 0x821  :  120 - 0x78
    "11100111", -- 2082 - 0x822  :  231 - 0xe7
    "11001111", -- 2083 - 0x823  :  207 - 0xcf
    "01011000", -- 2084 - 0x824  :   88 - 0x58
    "01011000", -- 2085 - 0x825  :   88 - 0x58
    "01010000", -- 2086 - 0x826  :   80 - 0x50
    "10010000", -- 2087 - 0x827  :  144 - 0x90
    "11000000", -- 2088 - 0x828  :  192 - 0xc0 -- plane 1
    "10000111", -- 2089 - 0x829  :  135 - 0x87
    "00011000", -- 2090 - 0x82a  :   24 - 0x18
    "10110000", -- 2091 - 0x82b  :  176 - 0xb0
    "11100111", -- 2092 - 0x82c  :  231 - 0xe7
    "11100111", -- 2093 - 0x82d  :  231 - 0xe7
    "11101111", -- 2094 - 0x82e  :  239 - 0xef
    "11101111", -- 2095 - 0x82f  :  239 - 0xef
    "10110000", -- 2096 - 0x830  :  176 - 0xb0 -- Background 0x83
    "11111100", -- 2097 - 0x831  :  252 - 0xfc
    "11100010", -- 2098 - 0x832  :  226 - 0xe2
    "11000001", -- 2099 - 0x833  :  193 - 0xc1
    "11000001", -- 2100 - 0x834  :  193 - 0xc1
    "10000011", -- 2101 - 0x835  :  131 - 0x83
    "10001111", -- 2102 - 0x836  :  143 - 0x8f
    "01111110", -- 2103 - 0x837  :  126 - 0x7e
    "01101111", -- 2104 - 0x838  :  111 - 0x6f -- plane 1
    "01000011", -- 2105 - 0x839  :   67 - 0x43
    "01011101", -- 2106 - 0x83a  :   93 - 0x5d
    "00111111", -- 2107 - 0x83b  :   63 - 0x3f
    "00111111", -- 2108 - 0x83c  :   63 - 0x3f
    "01111111", -- 2109 - 0x83d  :  127 - 0x7f
    "01111111", -- 2110 - 0x83e  :  127 - 0x7f
    "11111111", -- 2111 - 0x83f  :  255 - 0xff
    "11111110", -- 2112 - 0x840  :  254 - 0xfe -- Background 0x84
    "00000011", -- 2113 - 0x841  :    3 - 0x3
    "00001111", -- 2114 - 0x842  :   15 - 0xf
    "10010001", -- 2115 - 0x843  :  145 - 0x91
    "01110000", -- 2116 - 0x844  :  112 - 0x70
    "01100000", -- 2117 - 0x845  :   96 - 0x60
    "00100000", -- 2118 - 0x846  :   32 - 0x20
    "00110001", -- 2119 - 0x847  :   49 - 0x31
    "00000011", -- 2120 - 0x848  :    3 - 0x3 -- plane 1
    "11111111", -- 2121 - 0x849  :  255 - 0xff
    "11110001", -- 2122 - 0x84a  :  241 - 0xf1
    "01101110", -- 2123 - 0x84b  :  110 - 0x6e
    "11001111", -- 2124 - 0x84c  :  207 - 0xcf
    "11011111", -- 2125 - 0x84d  :  223 - 0xdf
    "11111111", -- 2126 - 0x84e  :  255 - 0xff
    "11111111", -- 2127 - 0x84f  :  255 - 0xff
    "00111111", -- 2128 - 0x850  :   63 - 0x3f -- Background 0x85
    "00111111", -- 2129 - 0x851  :   63 - 0x3f
    "00011101", -- 2130 - 0x852  :   29 - 0x1d
    "00111001", -- 2131 - 0x853  :   57 - 0x39
    "01111011", -- 2132 - 0x854  :  123 - 0x7b
    "11110011", -- 2133 - 0x855  :  243 - 0xf3
    "10000110", -- 2134 - 0x856  :  134 - 0x86
    "11111110", -- 2135 - 0x857  :  254 - 0xfe
    "11111101", -- 2136 - 0x858  :  253 - 0xfd -- plane 1
    "11111011", -- 2137 - 0x859  :  251 - 0xfb
    "11111011", -- 2138 - 0x85a  :  251 - 0xfb
    "11110111", -- 2139 - 0x85b  :  247 - 0xf7
    "11110111", -- 2140 - 0x85c  :  247 - 0xf7
    "00001111", -- 2141 - 0x85d  :   15 - 0xf
    "01111111", -- 2142 - 0x85e  :  127 - 0x7f
    "11111111", -- 2143 - 0x85f  :  255 - 0xff
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Background 0x86
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11111111", -- 2147 - 0x863  :  255 - 0xff
    "11111111", -- 2148 - 0x864  :  255 - 0xff
    "10000000", -- 2149 - 0x865  :  128 - 0x80
    "10000000", -- 2150 - 0x866  :  128 - 0x80
    "11111111", -- 2151 - 0x867  :  255 - 0xff
    "11111111", -- 2152 - 0x868  :  255 - 0xff -- plane 1
    "10000000", -- 2153 - 0x869  :  128 - 0x80
    "10000000", -- 2154 - 0x86a  :  128 - 0x80
    "10000000", -- 2155 - 0x86b  :  128 - 0x80
    "10000000", -- 2156 - 0x86c  :  128 - 0x80
    "11111111", -- 2157 - 0x86d  :  255 - 0xff
    "11111111", -- 2158 - 0x86e  :  255 - 0xff
    "10000000", -- 2159 - 0x86f  :  128 - 0x80
    "11111110", -- 2160 - 0x870  :  254 - 0xfe -- Background 0x87
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "00000011", -- 2165 - 0x875  :    3 - 0x3
    "00000011", -- 2166 - 0x876  :    3 - 0x3
    "11111111", -- 2167 - 0x877  :  255 - 0xff
    "11111110", -- 2168 - 0x878  :  254 - 0xfe -- plane 1
    "00000011", -- 2169 - 0x879  :    3 - 0x3
    "00000011", -- 2170 - 0x87a  :    3 - 0x3
    "00000011", -- 2171 - 0x87b  :    3 - 0x3
    "00000011", -- 2172 - 0x87c  :    3 - 0x3
    "11111111", -- 2173 - 0x87d  :  255 - 0xff
    "11111111", -- 2174 - 0x87e  :  255 - 0xff
    "00000011", -- 2175 - 0x87f  :    3 - 0x3
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Background 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "11111111", -- 2178 - 0x882  :  255 - 0xff
    "11111111", -- 2179 - 0x883  :  255 - 0xff
    "11111111", -- 2180 - 0x884  :  255 - 0xff
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "00000000", -- 2182 - 0x886  :    0 - 0x0
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "11111111", -- 2185 - 0x889  :  255 - 0xff
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "11111111", -- 2190 - 0x88e  :  255 - 0xff
    "11111111", -- 2191 - 0x88f  :  255 - 0xff
    "00111100", -- 2192 - 0x890  :   60 - 0x3c -- Background 0x89
    "11111100", -- 2193 - 0x891  :  252 - 0xfc
    "11111100", -- 2194 - 0x892  :  252 - 0xfc
    "11111100", -- 2195 - 0x893  :  252 - 0xfc
    "11111100", -- 2196 - 0x894  :  252 - 0xfc
    "11111100", -- 2197 - 0x895  :  252 - 0xfc
    "00000100", -- 2198 - 0x896  :    4 - 0x4
    "00000100", -- 2199 - 0x897  :    4 - 0x4
    "00100011", -- 2200 - 0x898  :   35 - 0x23 -- plane 1
    "11110011", -- 2201 - 0x899  :  243 - 0xf3
    "00001011", -- 2202 - 0x89a  :   11 - 0xb
    "00001011", -- 2203 - 0x89b  :   11 - 0xb
    "00001011", -- 2204 - 0x89c  :   11 - 0xb
    "00000111", -- 2205 - 0x89d  :    7 - 0x7
    "11111111", -- 2206 - 0x89e  :  255 - 0xff
    "11111111", -- 2207 - 0x89f  :  255 - 0xff
    "11111111", -- 2208 - 0x8a0  :  255 - 0xff -- Background 0x8a
    "11111111", -- 2209 - 0x8a1  :  255 - 0xff
    "11111111", -- 2210 - 0x8a2  :  255 - 0xff
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "10000000", -- 2212 - 0x8a4  :  128 - 0x80
    "11111111", -- 2213 - 0x8a5  :  255 - 0xff
    "11111111", -- 2214 - 0x8a6  :  255 - 0xff
    "11111111", -- 2215 - 0x8a7  :  255 - 0xff
    "10000000", -- 2216 - 0x8a8  :  128 - 0x80 -- plane 1
    "10000000", -- 2217 - 0x8a9  :  128 - 0x80
    "10000000", -- 2218 - 0x8aa  :  128 - 0x80
    "10000000", -- 2219 - 0x8ab  :  128 - 0x80
    "11111111", -- 2220 - 0x8ac  :  255 - 0xff
    "10000000", -- 2221 - 0x8ad  :  128 - 0x80
    "10000000", -- 2222 - 0x8ae  :  128 - 0x80
    "10000000", -- 2223 - 0x8af  :  128 - 0x80
    "11111111", -- 2224 - 0x8b0  :  255 - 0xff -- Background 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11111111", -- 2226 - 0x8b2  :  255 - 0xff
    "11111111", -- 2227 - 0x8b3  :  255 - 0xff
    "00000011", -- 2228 - 0x8b4  :    3 - 0x3
    "11111111", -- 2229 - 0x8b5  :  255 - 0xff
    "11111111", -- 2230 - 0x8b6  :  255 - 0xff
    "11111111", -- 2231 - 0x8b7  :  255 - 0xff
    "00000011", -- 2232 - 0x8b8  :    3 - 0x3 -- plane 1
    "00000011", -- 2233 - 0x8b9  :    3 - 0x3
    "00000011", -- 2234 - 0x8ba  :    3 - 0x3
    "00000011", -- 2235 - 0x8bb  :    3 - 0x3
    "11111111", -- 2236 - 0x8bc  :  255 - 0xff
    "00000011", -- 2237 - 0x8bd  :    3 - 0x3
    "00000011", -- 2238 - 0x8be  :    3 - 0x3
    "00000011", -- 2239 - 0x8bf  :    3 - 0x3
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Background 0x8c
    "11111111", -- 2241 - 0x8c1  :  255 - 0xff
    "11111111", -- 2242 - 0x8c2  :  255 - 0xff
    "11111111", -- 2243 - 0x8c3  :  255 - 0xff
    "11111111", -- 2244 - 0x8c4  :  255 - 0xff
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "11111111", -- 2246 - 0x8c6  :  255 - 0xff
    "11111111", -- 2247 - 0x8c7  :  255 - 0xff
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "11111111", -- 2253 - 0x8cd  :  255 - 0xff
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "11111100", -- 2256 - 0x8d0  :  252 - 0xfc -- Background 0x8d
    "11111100", -- 2257 - 0x8d1  :  252 - 0xfc
    "11111110", -- 2258 - 0x8d2  :  254 - 0xfe
    "11111110", -- 2259 - 0x8d3  :  254 - 0xfe
    "11111110", -- 2260 - 0x8d4  :  254 - 0xfe
    "00000010", -- 2261 - 0x8d5  :    2 - 0x2
    "11111110", -- 2262 - 0x8d6  :  254 - 0xfe
    "11111110", -- 2263 - 0x8d7  :  254 - 0xfe
    "00000111", -- 2264 - 0x8d8  :    7 - 0x7 -- plane 1
    "00000111", -- 2265 - 0x8d9  :    7 - 0x7
    "00000011", -- 2266 - 0x8da  :    3 - 0x3
    "00000011", -- 2267 - 0x8db  :    3 - 0x3
    "00000011", -- 2268 - 0x8dc  :    3 - 0x3
    "11111111", -- 2269 - 0x8dd  :  255 - 0xff
    "00000011", -- 2270 - 0x8de  :    3 - 0x3
    "00000011", -- 2271 - 0x8df  :    3 - 0x3
    "11111111", -- 2272 - 0x8e0  :  255 - 0xff -- Background 0x8e
    "10000000", -- 2273 - 0x8e1  :  128 - 0x80
    "10000000", -- 2274 - 0x8e2  :  128 - 0x80
    "10000000", -- 2275 - 0x8e3  :  128 - 0x80
    "10000000", -- 2276 - 0x8e4  :  128 - 0x80
    "10000000", -- 2277 - 0x8e5  :  128 - 0x80
    "10000000", -- 2278 - 0x8e6  :  128 - 0x80
    "10000000", -- 2279 - 0x8e7  :  128 - 0x80
    "10000000", -- 2280 - 0x8e8  :  128 - 0x80 -- plane 1
    "11111111", -- 2281 - 0x8e9  :  255 - 0xff
    "11111111", -- 2282 - 0x8ea  :  255 - 0xff
    "11111111", -- 2283 - 0x8eb  :  255 - 0xff
    "11111111", -- 2284 - 0x8ec  :  255 - 0xff
    "11111111", -- 2285 - 0x8ed  :  255 - 0xff
    "11111111", -- 2286 - 0x8ee  :  255 - 0xff
    "11111111", -- 2287 - 0x8ef  :  255 - 0xff
    "11111111", -- 2288 - 0x8f0  :  255 - 0xff -- Background 0x8f
    "00000011", -- 2289 - 0x8f1  :    3 - 0x3
    "00000011", -- 2290 - 0x8f2  :    3 - 0x3
    "00000011", -- 2291 - 0x8f3  :    3 - 0x3
    "00000011", -- 2292 - 0x8f4  :    3 - 0x3
    "00000011", -- 2293 - 0x8f5  :    3 - 0x3
    "00000011", -- 2294 - 0x8f6  :    3 - 0x3
    "00000011", -- 2295 - 0x8f7  :    3 - 0x3
    "00000011", -- 2296 - 0x8f8  :    3 - 0x3 -- plane 1
    "11111111", -- 2297 - 0x8f9  :  255 - 0xff
    "11111111", -- 2298 - 0x8fa  :  255 - 0xff
    "11111111", -- 2299 - 0x8fb  :  255 - 0xff
    "11111111", -- 2300 - 0x8fc  :  255 - 0xff
    "11111111", -- 2301 - 0x8fd  :  255 - 0xff
    "11111111", -- 2302 - 0x8fe  :  255 - 0xff
    "11111111", -- 2303 - 0x8ff  :  255 - 0xff
    "00000010", -- 2304 - 0x900  :    2 - 0x2 -- Background 0x90
    "00000010", -- 2305 - 0x901  :    2 - 0x2
    "00000010", -- 2306 - 0x902  :    2 - 0x2
    "00000010", -- 2307 - 0x903  :    2 - 0x2
    "00000010", -- 2308 - 0x904  :    2 - 0x2
    "00000010", -- 2309 - 0x905  :    2 - 0x2
    "00000100", -- 2310 - 0x906  :    4 - 0x4
    "00000100", -- 2311 - 0x907  :    4 - 0x4
    "11111111", -- 2312 - 0x908  :  255 - 0xff -- plane 1
    "11111111", -- 2313 - 0x909  :  255 - 0xff
    "11111111", -- 2314 - 0x90a  :  255 - 0xff
    "11111111", -- 2315 - 0x90b  :  255 - 0xff
    "11111111", -- 2316 - 0x90c  :  255 - 0xff
    "11111111", -- 2317 - 0x90d  :  255 - 0xff
    "11111111", -- 2318 - 0x90e  :  255 - 0xff
    "11111111", -- 2319 - 0x90f  :  255 - 0xff
    "10000000", -- 2320 - 0x910  :  128 - 0x80 -- Background 0x91
    "10000000", -- 2321 - 0x911  :  128 - 0x80
    "10101010", -- 2322 - 0x912  :  170 - 0xaa
    "11010101", -- 2323 - 0x913  :  213 - 0xd5
    "10101010", -- 2324 - 0x914  :  170 - 0xaa
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "11111111", -- 2326 - 0x916  :  255 - 0xff
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "11111111", -- 2328 - 0x918  :  255 - 0xff -- plane 1
    "11111111", -- 2329 - 0x919  :  255 - 0xff
    "11010101", -- 2330 - 0x91a  :  213 - 0xd5
    "10101010", -- 2331 - 0x91b  :  170 - 0xaa
    "11010101", -- 2332 - 0x91c  :  213 - 0xd5
    "10000000", -- 2333 - 0x91d  :  128 - 0x80
    "10000000", -- 2334 - 0x91e  :  128 - 0x80
    "11111111", -- 2335 - 0x91f  :  255 - 0xff
    "00000011", -- 2336 - 0x920  :    3 - 0x3 -- Background 0x92
    "00000011", -- 2337 - 0x921  :    3 - 0x3
    "10101011", -- 2338 - 0x922  :  171 - 0xab
    "01010111", -- 2339 - 0x923  :   87 - 0x57
    "10101011", -- 2340 - 0x924  :  171 - 0xab
    "11111111", -- 2341 - 0x925  :  255 - 0xff
    "11111111", -- 2342 - 0x926  :  255 - 0xff
    "11111110", -- 2343 - 0x927  :  254 - 0xfe
    "11111111", -- 2344 - 0x928  :  255 - 0xff -- plane 1
    "11111111", -- 2345 - 0x929  :  255 - 0xff
    "01010111", -- 2346 - 0x92a  :   87 - 0x57
    "10101011", -- 2347 - 0x92b  :  171 - 0xab
    "01010111", -- 2348 - 0x92c  :   87 - 0x57
    "00000011", -- 2349 - 0x92d  :    3 - 0x3
    "00000011", -- 2350 - 0x92e  :    3 - 0x3
    "11111110", -- 2351 - 0x92f  :  254 - 0xfe
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x93
    "01010101", -- 2353 - 0x931  :   85 - 0x55
    "10101010", -- 2354 - 0x932  :  170 - 0xaa
    "01010101", -- 2355 - 0x933  :   85 - 0x55
    "11111111", -- 2356 - 0x934  :  255 - 0xff
    "11111111", -- 2357 - 0x935  :  255 - 0xff
    "11111111", -- 2358 - 0x936  :  255 - 0xff
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "11111111", -- 2360 - 0x938  :  255 - 0xff -- plane 1
    "10101010", -- 2361 - 0x939  :  170 - 0xaa
    "01010101", -- 2362 - 0x93a  :   85 - 0x55
    "10101010", -- 2363 - 0x93b  :  170 - 0xaa
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000100", -- 2368 - 0x940  :    4 - 0x4 -- Background 0x94
    "01010100", -- 2369 - 0x941  :   84 - 0x54
    "10101100", -- 2370 - 0x942  :  172 - 0xac
    "01011100", -- 2371 - 0x943  :   92 - 0x5c
    "11111100", -- 2372 - 0x944  :  252 - 0xfc
    "11111100", -- 2373 - 0x945  :  252 - 0xfc
    "11111100", -- 2374 - 0x946  :  252 - 0xfc
    "00111100", -- 2375 - 0x947  :   60 - 0x3c
    "11111111", -- 2376 - 0x948  :  255 - 0xff -- plane 1
    "10101111", -- 2377 - 0x949  :  175 - 0xaf
    "01010111", -- 2378 - 0x94a  :   87 - 0x57
    "10101011", -- 2379 - 0x94b  :  171 - 0xab
    "00001011", -- 2380 - 0x94c  :   11 - 0xb
    "00001011", -- 2381 - 0x94d  :   11 - 0xb
    "11110011", -- 2382 - 0x94e  :  243 - 0xf3
    "00100011", -- 2383 - 0x94f  :   35 - 0x23
    "00111111", -- 2384 - 0x950  :   63 - 0x3f -- Background 0x95
    "00111111", -- 2385 - 0x951  :   63 - 0x3f
    "00111111", -- 2386 - 0x952  :   63 - 0x3f
    "00111111", -- 2387 - 0x953  :   63 - 0x3f
    "00000000", -- 2388 - 0x954  :    0 - 0x0
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "11111111", -- 2391 - 0x957  :  255 - 0xff
    "11111111", -- 2392 - 0x958  :  255 - 0xff -- plane 1
    "11111111", -- 2393 - 0x959  :  255 - 0xff
    "11111111", -- 2394 - 0x95a  :  255 - 0xff
    "11111111", -- 2395 - 0x95b  :  255 - 0xff
    "11111111", -- 2396 - 0x95c  :  255 - 0xff
    "11111111", -- 2397 - 0x95d  :  255 - 0xff
    "11111111", -- 2398 - 0x95e  :  255 - 0xff
    "11111111", -- 2399 - 0x95f  :  255 - 0xff
    "01111110", -- 2400 - 0x960  :  126 - 0x7e -- Background 0x96
    "01111100", -- 2401 - 0x961  :  124 - 0x7c
    "01111100", -- 2402 - 0x962  :  124 - 0x7c
    "01111000", -- 2403 - 0x963  :  120 - 0x78
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "11111111", -- 2407 - 0x967  :  255 - 0xff
    "11111111", -- 2408 - 0x968  :  255 - 0xff -- plane 1
    "11111111", -- 2409 - 0x969  :  255 - 0xff
    "11111111", -- 2410 - 0x96a  :  255 - 0xff
    "11111111", -- 2411 - 0x96b  :  255 - 0xff
    "11111111", -- 2412 - 0x96c  :  255 - 0xff
    "11111111", -- 2413 - 0x96d  :  255 - 0xff
    "11111111", -- 2414 - 0x96e  :  255 - 0xff
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00011111", -- 2416 - 0x970  :   31 - 0x1f -- Background 0x97
    "00001111", -- 2417 - 0x971  :   15 - 0xf
    "00001111", -- 2418 - 0x972  :   15 - 0xf
    "00000111", -- 2419 - 0x973  :    7 - 0x7
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "11111111", -- 2423 - 0x977  :  255 - 0xff
    "11111111", -- 2424 - 0x978  :  255 - 0xff -- plane 1
    "11111111", -- 2425 - 0x979  :  255 - 0xff
    "11111111", -- 2426 - 0x97a  :  255 - 0xff
    "11111111", -- 2427 - 0x97b  :  255 - 0xff
    "11111111", -- 2428 - 0x97c  :  255 - 0xff
    "11111111", -- 2429 - 0x97d  :  255 - 0xff
    "11111111", -- 2430 - 0x97e  :  255 - 0xff
    "11111111", -- 2431 - 0x97f  :  255 - 0xff
    "11111110", -- 2432 - 0x980  :  254 - 0xfe -- Background 0x98
    "11111100", -- 2433 - 0x981  :  252 - 0xfc
    "11111100", -- 2434 - 0x982  :  252 - 0xfc
    "11111000", -- 2435 - 0x983  :  248 - 0xf8
    "00000000", -- 2436 - 0x984  :    0 - 0x0
    "00000000", -- 2437 - 0x985  :    0 - 0x0
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "11111111", -- 2440 - 0x988  :  255 - 0xff -- plane 1
    "11111111", -- 2441 - 0x989  :  255 - 0xff
    "11111111", -- 2442 - 0x98a  :  255 - 0xff
    "11111111", -- 2443 - 0x98b  :  255 - 0xff
    "11111111", -- 2444 - 0x98c  :  255 - 0xff
    "11111111", -- 2445 - 0x98d  :  255 - 0xff
    "11111111", -- 2446 - 0x98e  :  255 - 0xff
    "11111111", -- 2447 - 0x98f  :  255 - 0xff
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Background 0x99
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "11111111", -- 2452 - 0x994  :  255 - 0xff
    "11111111", -- 2453 - 0x995  :  255 - 0xff
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "00000000", -- 2456 - 0x998  :    0 - 0x0 -- plane 1
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00011000", -- 2464 - 0x9a0  :   24 - 0x18 -- Background 0x9a
    "00011000", -- 2465 - 0x9a1  :   24 - 0x18
    "00011000", -- 2466 - 0x9a2  :   24 - 0x18
    "00011000", -- 2467 - 0x9a3  :   24 - 0x18
    "00011000", -- 2468 - 0x9a4  :   24 - 0x18
    "00011000", -- 2469 - 0x9a5  :   24 - 0x18
    "00011000", -- 2470 - 0x9a6  :   24 - 0x18
    "00011000", -- 2471 - 0x9a7  :   24 - 0x18
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000111", -- 2480 - 0x9b0  :    7 - 0x7 -- Background 0x9b
    "00011111", -- 2481 - 0x9b1  :   31 - 0x1f
    "00111111", -- 2482 - 0x9b2  :   63 - 0x3f
    "11111111", -- 2483 - 0x9b3  :  255 - 0xff
    "01111111", -- 2484 - 0x9b4  :  127 - 0x7f
    "01111111", -- 2485 - 0x9b5  :  127 - 0x7f
    "11111111", -- 2486 - 0x9b6  :  255 - 0xff
    "11111111", -- 2487 - 0x9b7  :  255 - 0xff
    "11111111", -- 2488 - 0x9b8  :  255 - 0xff -- plane 1
    "11111111", -- 2489 - 0x9b9  :  255 - 0xff
    "11111111", -- 2490 - 0x9ba  :  255 - 0xff
    "11111111", -- 2491 - 0x9bb  :  255 - 0xff
    "11111111", -- 2492 - 0x9bc  :  255 - 0xff
    "11111111", -- 2493 - 0x9bd  :  255 - 0xff
    "11111111", -- 2494 - 0x9be  :  255 - 0xff
    "11111111", -- 2495 - 0x9bf  :  255 - 0xff
    "11100001", -- 2496 - 0x9c0  :  225 - 0xe1 -- Background 0x9c
    "11111001", -- 2497 - 0x9c1  :  249 - 0xf9
    "11111101", -- 2498 - 0x9c2  :  253 - 0xfd
    "11111111", -- 2499 - 0x9c3  :  255 - 0xff
    "11111110", -- 2500 - 0x9c4  :  254 - 0xfe
    "11111110", -- 2501 - 0x9c5  :  254 - 0xfe
    "11111111", -- 2502 - 0x9c6  :  255 - 0xff
    "11111111", -- 2503 - 0x9c7  :  255 - 0xff
    "11111111", -- 2504 - 0x9c8  :  255 - 0xff -- plane 1
    "11111111", -- 2505 - 0x9c9  :  255 - 0xff
    "11111111", -- 2506 - 0x9ca  :  255 - 0xff
    "11111111", -- 2507 - 0x9cb  :  255 - 0xff
    "11111111", -- 2508 - 0x9cc  :  255 - 0xff
    "11111111", -- 2509 - 0x9cd  :  255 - 0xff
    "11111111", -- 2510 - 0x9ce  :  255 - 0xff
    "11111111", -- 2511 - 0x9cf  :  255 - 0xff
    "11110000", -- 2512 - 0x9d0  :  240 - 0xf0 -- Background 0x9d
    "00010000", -- 2513 - 0x9d1  :   16 - 0x10
    "00010000", -- 2514 - 0x9d2  :   16 - 0x10
    "00010000", -- 2515 - 0x9d3  :   16 - 0x10
    "00010000", -- 2516 - 0x9d4  :   16 - 0x10
    "00010000", -- 2517 - 0x9d5  :   16 - 0x10
    "00010000", -- 2518 - 0x9d6  :   16 - 0x10
    "11111111", -- 2519 - 0x9d7  :  255 - 0xff
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- plane 1
    "11100000", -- 2521 - 0x9d9  :  224 - 0xe0
    "11100000", -- 2522 - 0x9da  :  224 - 0xe0
    "11100000", -- 2523 - 0x9db  :  224 - 0xe0
    "11100000", -- 2524 - 0x9dc  :  224 - 0xe0
    "11100000", -- 2525 - 0x9dd  :  224 - 0xe0
    "11100000", -- 2526 - 0x9de  :  224 - 0xe0
    "11100000", -- 2527 - 0x9df  :  224 - 0xe0
    "00011111", -- 2528 - 0x9e0  :   31 - 0x1f -- Background 0x9e
    "00010000", -- 2529 - 0x9e1  :   16 - 0x10
    "00010000", -- 2530 - 0x9e2  :   16 - 0x10
    "00010000", -- 2531 - 0x9e3  :   16 - 0x10
    "00010000", -- 2532 - 0x9e4  :   16 - 0x10
    "00010000", -- 2533 - 0x9e5  :   16 - 0x10
    "00010000", -- 2534 - 0x9e6  :   16 - 0x10
    "11111111", -- 2535 - 0x9e7  :  255 - 0xff
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- plane 1
    "00001111", -- 2537 - 0x9e9  :   15 - 0xf
    "00001111", -- 2538 - 0x9ea  :   15 - 0xf
    "00001111", -- 2539 - 0x9eb  :   15 - 0xf
    "00001111", -- 2540 - 0x9ec  :   15 - 0xf
    "00001111", -- 2541 - 0x9ed  :   15 - 0xf
    "00001111", -- 2542 - 0x9ee  :   15 - 0xf
    "00001111", -- 2543 - 0x9ef  :   15 - 0xf
    "10010010", -- 2544 - 0x9f0  :  146 - 0x92 -- Background 0x9f
    "10010010", -- 2545 - 0x9f1  :  146 - 0x92
    "10010010", -- 2546 - 0x9f2  :  146 - 0x92
    "11111110", -- 2547 - 0x9f3  :  254 - 0xfe
    "11111110", -- 2548 - 0x9f4  :  254 - 0xfe
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "01001000", -- 2552 - 0x9f8  :   72 - 0x48 -- plane 1
    "01001000", -- 2553 - 0x9f9  :   72 - 0x48
    "01101100", -- 2554 - 0x9fa  :  108 - 0x6c
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "11111110", -- 2558 - 0x9fe  :  254 - 0xfe
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00001010", -- 2560 - 0xa00  :   10 - 0xa -- Background 0xa0
    "00001010", -- 2561 - 0xa01  :   10 - 0xa
    "00111010", -- 2562 - 0xa02  :   58 - 0x3a
    "00001010", -- 2563 - 0xa03  :   10 - 0xa
    "11111011", -- 2564 - 0xa04  :  251 - 0xfb
    "00001011", -- 2565 - 0xa05  :   11 - 0xb
    "00001011", -- 2566 - 0xa06  :   11 - 0xb
    "00001011", -- 2567 - 0xa07  :   11 - 0xb
    "00000101", -- 2568 - 0xa08  :    5 - 0x5 -- plane 1
    "00000101", -- 2569 - 0xa09  :    5 - 0x5
    "11000101", -- 2570 - 0xa0a  :  197 - 0xc5
    "11110101", -- 2571 - 0xa0b  :  245 - 0xf5
    "11110100", -- 2572 - 0xa0c  :  244 - 0xf4
    "00000100", -- 2573 - 0xa0d  :    4 - 0x4
    "00000100", -- 2574 - 0xa0e  :    4 - 0x4
    "00000100", -- 2575 - 0xa0f  :    4 - 0x4
    "10010000", -- 2576 - 0xa10  :  144 - 0x90 -- Background 0xa1
    "10010000", -- 2577 - 0xa11  :  144 - 0x90
    "10011111", -- 2578 - 0xa12  :  159 - 0x9f
    "10010000", -- 2579 - 0xa13  :  144 - 0x90
    "10011111", -- 2580 - 0xa14  :  159 - 0x9f
    "10010000", -- 2581 - 0xa15  :  144 - 0x90
    "10010000", -- 2582 - 0xa16  :  144 - 0x90
    "10010000", -- 2583 - 0xa17  :  144 - 0x90
    "01110000", -- 2584 - 0xa18  :  112 - 0x70 -- plane 1
    "01110000", -- 2585 - 0xa19  :  112 - 0x70
    "01110000", -- 2586 - 0xa1a  :  112 - 0x70
    "01111111", -- 2587 - 0xa1b  :  127 - 0x7f
    "01111111", -- 2588 - 0xa1c  :  127 - 0x7f
    "01110000", -- 2589 - 0xa1d  :  112 - 0x70
    "01110000", -- 2590 - 0xa1e  :  112 - 0x70
    "01110000", -- 2591 - 0xa1f  :  112 - 0x70
    "00000001", -- 2592 - 0xa20  :    1 - 0x1 -- Background 0xa2
    "00000001", -- 2593 - 0xa21  :    1 - 0x1
    "00000001", -- 2594 - 0xa22  :    1 - 0x1
    "00000001", -- 2595 - 0xa23  :    1 - 0x1
    "00000001", -- 2596 - 0xa24  :    1 - 0x1
    "00000001", -- 2597 - 0xa25  :    1 - 0x1
    "00000001", -- 2598 - 0xa26  :    1 - 0x1
    "00000001", -- 2599 - 0xa27  :    1 - 0x1
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- plane 1
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "10000000", -- 2608 - 0xa30  :  128 - 0x80 -- Background 0xa3
    "10000000", -- 2609 - 0xa31  :  128 - 0x80
    "10000000", -- 2610 - 0xa32  :  128 - 0x80
    "10000000", -- 2611 - 0xa33  :  128 - 0x80
    "10000000", -- 2612 - 0xa34  :  128 - 0x80
    "10000000", -- 2613 - 0xa35  :  128 - 0x80
    "10000000", -- 2614 - 0xa36  :  128 - 0x80
    "10000000", -- 2615 - 0xa37  :  128 - 0x80
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- plane 1
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00001000", -- 2624 - 0xa40  :    8 - 0x8 -- Background 0xa4
    "10001000", -- 2625 - 0xa41  :  136 - 0x88
    "10010001", -- 2626 - 0xa42  :  145 - 0x91
    "11010001", -- 2627 - 0xa43  :  209 - 0xd1
    "01010011", -- 2628 - 0xa44  :   83 - 0x53
    "01010011", -- 2629 - 0xa45  :   83 - 0x53
    "01110011", -- 2630 - 0xa46  :  115 - 0x73
    "00111111", -- 2631 - 0xa47  :   63 - 0x3f
    "11111111", -- 2632 - 0xa48  :  255 - 0xff -- plane 1
    "11111111", -- 2633 - 0xa49  :  255 - 0xff
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11111111", -- 2635 - 0xa4b  :  255 - 0xff
    "11111111", -- 2636 - 0xa4c  :  255 - 0xff
    "11111110", -- 2637 - 0xa4d  :  254 - 0xfe
    "10111110", -- 2638 - 0xa4e  :  190 - 0xbe
    "11001110", -- 2639 - 0xa4f  :  206 - 0xce
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000111", -- 2642 - 0xa52  :    7 - 0x7
    "00001111", -- 2643 - 0xa53  :   15 - 0xf
    "00001100", -- 2644 - 0xa54  :   12 - 0xc
    "00011011", -- 2645 - 0xa55  :   27 - 0x1b
    "00011011", -- 2646 - 0xa56  :   27 - 0x1b
    "00011011", -- 2647 - 0xa57  :   27 - 0x1b
    "00000000", -- 2648 - 0xa58  :    0 - 0x0 -- plane 1
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000011", -- 2652 - 0xa5c  :    3 - 0x3
    "00000100", -- 2653 - 0xa5d  :    4 - 0x4
    "00000100", -- 2654 - 0xa5e  :    4 - 0x4
    "00000100", -- 2655 - 0xa5f  :    4 - 0x4
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "11100000", -- 2658 - 0xa62  :  224 - 0xe0
    "11110000", -- 2659 - 0xa63  :  240 - 0xf0
    "11110000", -- 2660 - 0xa64  :  240 - 0xf0
    "11111000", -- 2661 - 0xa65  :  248 - 0xf8
    "11111000", -- 2662 - 0xa66  :  248 - 0xf8
    "11111000", -- 2663 - 0xa67  :  248 - 0xf8
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- plane 1
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "01100000", -- 2666 - 0xa6a  :   96 - 0x60
    "00110000", -- 2667 - 0xa6b  :   48 - 0x30
    "00110000", -- 2668 - 0xa6c  :   48 - 0x30
    "10011000", -- 2669 - 0xa6d  :  152 - 0x98
    "10011000", -- 2670 - 0xa6e  :  152 - 0x98
    "10011000", -- 2671 - 0xa6f  :  152 - 0x98
    "00011011", -- 2672 - 0xa70  :   27 - 0x1b -- Background 0xa7
    "00011011", -- 2673 - 0xa71  :   27 - 0x1b
    "00011011", -- 2674 - 0xa72  :   27 - 0x1b
    "00011011", -- 2675 - 0xa73  :   27 - 0x1b
    "00011011", -- 2676 - 0xa74  :   27 - 0x1b
    "00001111", -- 2677 - 0xa75  :   15 - 0xf
    "00001111", -- 2678 - 0xa76  :   15 - 0xf
    "00000111", -- 2679 - 0xa77  :    7 - 0x7
    "00000100", -- 2680 - 0xa78  :    4 - 0x4 -- plane 1
    "00000100", -- 2681 - 0xa79  :    4 - 0x4
    "00000100", -- 2682 - 0xa7a  :    4 - 0x4
    "00000100", -- 2683 - 0xa7b  :    4 - 0x4
    "00000100", -- 2684 - 0xa7c  :    4 - 0x4
    "00000011", -- 2685 - 0xa7d  :    3 - 0x3
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "11111000", -- 2688 - 0xa80  :  248 - 0xf8 -- Background 0xa8
    "11111000", -- 2689 - 0xa81  :  248 - 0xf8
    "11111000", -- 2690 - 0xa82  :  248 - 0xf8
    "11111000", -- 2691 - 0xa83  :  248 - 0xf8
    "11111000", -- 2692 - 0xa84  :  248 - 0xf8
    "11110000", -- 2693 - 0xa85  :  240 - 0xf0
    "11110000", -- 2694 - 0xa86  :  240 - 0xf0
    "11100000", -- 2695 - 0xa87  :  224 - 0xe0
    "10011000", -- 2696 - 0xa88  :  152 - 0x98 -- plane 1
    "10011000", -- 2697 - 0xa89  :  152 - 0x98
    "10011000", -- 2698 - 0xa8a  :  152 - 0x98
    "10011000", -- 2699 - 0xa8b  :  152 - 0x98
    "10011000", -- 2700 - 0xa8c  :  152 - 0x98
    "00110000", -- 2701 - 0xa8d  :   48 - 0x30
    "00110000", -- 2702 - 0xa8e  :   48 - 0x30
    "01100000", -- 2703 - 0xa8f  :   96 - 0x60
    "11110001", -- 2704 - 0xa90  :  241 - 0xf1 -- Background 0xa9
    "00010001", -- 2705 - 0xa91  :   17 - 0x11
    "00010001", -- 2706 - 0xa92  :   17 - 0x11
    "00011111", -- 2707 - 0xa93  :   31 - 0x1f
    "00010000", -- 2708 - 0xa94  :   16 - 0x10
    "00010000", -- 2709 - 0xa95  :   16 - 0x10
    "00010000", -- 2710 - 0xa96  :   16 - 0x10
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "00001111", -- 2712 - 0xa98  :   15 - 0xf -- plane 1
    "11101111", -- 2713 - 0xa99  :  239 - 0xef
    "11101111", -- 2714 - 0xa9a  :  239 - 0xef
    "11101111", -- 2715 - 0xa9b  :  239 - 0xef
    "11101111", -- 2716 - 0xa9c  :  239 - 0xef
    "11101111", -- 2717 - 0xa9d  :  239 - 0xef
    "11101111", -- 2718 - 0xa9e  :  239 - 0xef
    "11100000", -- 2719 - 0xa9f  :  224 - 0xe0
    "00011111", -- 2720 - 0xaa0  :   31 - 0x1f -- Background 0xaa
    "00010000", -- 2721 - 0xaa1  :   16 - 0x10
    "00010000", -- 2722 - 0xaa2  :   16 - 0x10
    "11110000", -- 2723 - 0xaa3  :  240 - 0xf0
    "00010000", -- 2724 - 0xaa4  :   16 - 0x10
    "00010000", -- 2725 - 0xaa5  :   16 - 0x10
    "00010000", -- 2726 - 0xaa6  :   16 - 0x10
    "11111111", -- 2727 - 0xaa7  :  255 - 0xff
    "11100000", -- 2728 - 0xaa8  :  224 - 0xe0 -- plane 1
    "11101111", -- 2729 - 0xaa9  :  239 - 0xef
    "11101111", -- 2730 - 0xaaa  :  239 - 0xef
    "11101111", -- 2731 - 0xaab  :  239 - 0xef
    "11101111", -- 2732 - 0xaac  :  239 - 0xef
    "11101111", -- 2733 - 0xaad  :  239 - 0xef
    "11101111", -- 2734 - 0xaae  :  239 - 0xef
    "00001111", -- 2735 - 0xaaf  :   15 - 0xf
    "01111111", -- 2736 - 0xab0  :  127 - 0x7f -- Background 0xab
    "10111111", -- 2737 - 0xab1  :  191 - 0xbf
    "11011111", -- 2738 - 0xab2  :  223 - 0xdf
    "11101111", -- 2739 - 0xab3  :  239 - 0xef
    "11110000", -- 2740 - 0xab4  :  240 - 0xf0
    "11110000", -- 2741 - 0xab5  :  240 - 0xf0
    "11110000", -- 2742 - 0xab6  :  240 - 0xf0
    "11110000", -- 2743 - 0xab7  :  240 - 0xf0
    "10000000", -- 2744 - 0xab8  :  128 - 0x80 -- plane 1
    "01000000", -- 2745 - 0xab9  :   64 - 0x40
    "00100000", -- 2746 - 0xaba  :   32 - 0x20
    "00010000", -- 2747 - 0xabb  :   16 - 0x10
    "00001111", -- 2748 - 0xabc  :   15 - 0xf
    "00001111", -- 2749 - 0xabd  :   15 - 0xf
    "00001111", -- 2750 - 0xabe  :   15 - 0xf
    "00001111", -- 2751 - 0xabf  :   15 - 0xf
    "11110000", -- 2752 - 0xac0  :  240 - 0xf0 -- Background 0xac
    "11110000", -- 2753 - 0xac1  :  240 - 0xf0
    "11110000", -- 2754 - 0xac2  :  240 - 0xf0
    "11110000", -- 2755 - 0xac3  :  240 - 0xf0
    "11111111", -- 2756 - 0xac4  :  255 - 0xff
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "11111111", -- 2758 - 0xac6  :  255 - 0xff
    "11111111", -- 2759 - 0xac7  :  255 - 0xff
    "00001111", -- 2760 - 0xac8  :   15 - 0xf -- plane 1
    "00001111", -- 2761 - 0xac9  :   15 - 0xf
    "00001111", -- 2762 - 0xaca  :   15 - 0xf
    "00001111", -- 2763 - 0xacb  :   15 - 0xf
    "00011111", -- 2764 - 0xacc  :   31 - 0x1f
    "00111111", -- 2765 - 0xacd  :   63 - 0x3f
    "01111111", -- 2766 - 0xace  :  127 - 0x7f
    "11111111", -- 2767 - 0xacf  :  255 - 0xff
    "11111111", -- 2768 - 0xad0  :  255 - 0xff -- Background 0xad
    "11111111", -- 2769 - 0xad1  :  255 - 0xff
    "11111111", -- 2770 - 0xad2  :  255 - 0xff
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "00001111", -- 2772 - 0xad4  :   15 - 0xf
    "00001111", -- 2773 - 0xad5  :   15 - 0xf
    "00001111", -- 2774 - 0xad6  :   15 - 0xf
    "00001111", -- 2775 - 0xad7  :   15 - 0xf
    "00000001", -- 2776 - 0xad8  :    1 - 0x1 -- plane 1
    "00000011", -- 2777 - 0xad9  :    3 - 0x3
    "00000111", -- 2778 - 0xada  :    7 - 0x7
    "00001111", -- 2779 - 0xadb  :   15 - 0xf
    "11111111", -- 2780 - 0xadc  :  255 - 0xff
    "11111111", -- 2781 - 0xadd  :  255 - 0xff
    "11111111", -- 2782 - 0xade  :  255 - 0xff
    "11111111", -- 2783 - 0xadf  :  255 - 0xff
    "00001111", -- 2784 - 0xae0  :   15 - 0xf -- Background 0xae
    "00001111", -- 2785 - 0xae1  :   15 - 0xf
    "00001111", -- 2786 - 0xae2  :   15 - 0xf
    "00001111", -- 2787 - 0xae3  :   15 - 0xf
    "11110111", -- 2788 - 0xae4  :  247 - 0xf7
    "11111011", -- 2789 - 0xae5  :  251 - 0xfb
    "11111101", -- 2790 - 0xae6  :  253 - 0xfd
    "11111110", -- 2791 - 0xae7  :  254 - 0xfe
    "11111111", -- 2792 - 0xae8  :  255 - 0xff -- plane 1
    "11111111", -- 2793 - 0xae9  :  255 - 0xff
    "11111111", -- 2794 - 0xaea  :  255 - 0xff
    "11111111", -- 2795 - 0xaeb  :  255 - 0xff
    "11111111", -- 2796 - 0xaec  :  255 - 0xff
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "11111111", -- 2798 - 0xaee  :  255 - 0xff
    "11111111", -- 2799 - 0xaef  :  255 - 0xff
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "00000000", -- 2802 - 0xaf2  :    0 - 0x0
    "00000000", -- 2803 - 0xaf3  :    0 - 0x0
    "00000000", -- 2804 - 0xaf4  :    0 - 0x0
    "00000000", -- 2805 - 0xaf5  :    0 - 0x0
    "00011000", -- 2806 - 0xaf6  :   24 - 0x18
    "00011000", -- 2807 - 0xaf7  :   24 - 0x18
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- plane 1
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00011111", -- 2816 - 0xb00  :   31 - 0x1f -- Background 0xb0
    "00111111", -- 2817 - 0xb01  :   63 - 0x3f
    "01111111", -- 2818 - 0xb02  :  127 - 0x7f
    "01111111", -- 2819 - 0xb03  :  127 - 0x7f
    "01111111", -- 2820 - 0xb04  :  127 - 0x7f
    "11111111", -- 2821 - 0xb05  :  255 - 0xff
    "11111111", -- 2822 - 0xb06  :  255 - 0xff
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "00011111", -- 2824 - 0xb08  :   31 - 0x1f -- plane 1
    "00100000", -- 2825 - 0xb09  :   32 - 0x20
    "01000000", -- 2826 - 0xb0a  :   64 - 0x40
    "01000000", -- 2827 - 0xb0b  :   64 - 0x40
    "01000000", -- 2828 - 0xb0c  :   64 - 0x40
    "10000000", -- 2829 - 0xb0d  :  128 - 0x80
    "10000010", -- 2830 - 0xb0e  :  130 - 0x82
    "10000010", -- 2831 - 0xb0f  :  130 - 0x82
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Background 0xb1
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "11111111", -- 2834 - 0xb12  :  255 - 0xff
    "01111111", -- 2835 - 0xb13  :  127 - 0x7f
    "01111111", -- 2836 - 0xb14  :  127 - 0x7f
    "01111111", -- 2837 - 0xb15  :  127 - 0x7f
    "00111111", -- 2838 - 0xb16  :   63 - 0x3f
    "00011110", -- 2839 - 0xb17  :   30 - 0x1e
    "10000010", -- 2840 - 0xb18  :  130 - 0x82 -- plane 1
    "10000000", -- 2841 - 0xb19  :  128 - 0x80
    "10100000", -- 2842 - 0xb1a  :  160 - 0xa0
    "01000100", -- 2843 - 0xb1b  :   68 - 0x44
    "01000011", -- 2844 - 0xb1c  :   67 - 0x43
    "01000000", -- 2845 - 0xb1d  :   64 - 0x40
    "00100001", -- 2846 - 0xb1e  :   33 - 0x21
    "00011110", -- 2847 - 0xb1f  :   30 - 0x1e
    "11111000", -- 2848 - 0xb20  :  248 - 0xf8 -- Background 0xb2
    "11111100", -- 2849 - 0xb21  :  252 - 0xfc
    "11111110", -- 2850 - 0xb22  :  254 - 0xfe
    "11111110", -- 2851 - 0xb23  :  254 - 0xfe
    "11111110", -- 2852 - 0xb24  :  254 - 0xfe
    "11111111", -- 2853 - 0xb25  :  255 - 0xff
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "11111111", -- 2855 - 0xb27  :  255 - 0xff
    "11111000", -- 2856 - 0xb28  :  248 - 0xf8 -- plane 1
    "00000100", -- 2857 - 0xb29  :    4 - 0x4
    "00000010", -- 2858 - 0xb2a  :    2 - 0x2
    "00000010", -- 2859 - 0xb2b  :    2 - 0x2
    "00000010", -- 2860 - 0xb2c  :    2 - 0x2
    "00000001", -- 2861 - 0xb2d  :    1 - 0x1
    "01000001", -- 2862 - 0xb2e  :   65 - 0x41
    "01000001", -- 2863 - 0xb2f  :   65 - 0x41
    "11111111", -- 2864 - 0xb30  :  255 - 0xff -- Background 0xb3
    "11111111", -- 2865 - 0xb31  :  255 - 0xff
    "11111111", -- 2866 - 0xb32  :  255 - 0xff
    "11111110", -- 2867 - 0xb33  :  254 - 0xfe
    "11111110", -- 2868 - 0xb34  :  254 - 0xfe
    "11111110", -- 2869 - 0xb35  :  254 - 0xfe
    "11111100", -- 2870 - 0xb36  :  252 - 0xfc
    "01111000", -- 2871 - 0xb37  :  120 - 0x78
    "01000001", -- 2872 - 0xb38  :   65 - 0x41 -- plane 1
    "00000001", -- 2873 - 0xb39  :    1 - 0x1
    "00000101", -- 2874 - 0xb3a  :    5 - 0x5
    "00100010", -- 2875 - 0xb3b  :   34 - 0x22
    "11000010", -- 2876 - 0xb3c  :  194 - 0xc2
    "00000010", -- 2877 - 0xb3d  :    2 - 0x2
    "10000100", -- 2878 - 0xb3e  :  132 - 0x84
    "01111000", -- 2879 - 0xb3f  :  120 - 0x78
    "01111111", -- 2880 - 0xb40  :  127 - 0x7f -- Background 0xb4
    "10000000", -- 2881 - 0xb41  :  128 - 0x80
    "10000000", -- 2882 - 0xb42  :  128 - 0x80
    "10000000", -- 2883 - 0xb43  :  128 - 0x80
    "10000000", -- 2884 - 0xb44  :  128 - 0x80
    "10000000", -- 2885 - 0xb45  :  128 - 0x80
    "10000000", -- 2886 - 0xb46  :  128 - 0x80
    "10000000", -- 2887 - 0xb47  :  128 - 0x80
    "10000000", -- 2888 - 0xb48  :  128 - 0x80 -- plane 1
    "01111111", -- 2889 - 0xb49  :  127 - 0x7f
    "01111111", -- 2890 - 0xb4a  :  127 - 0x7f
    "01111111", -- 2891 - 0xb4b  :  127 - 0x7f
    "01111111", -- 2892 - 0xb4c  :  127 - 0x7f
    "01111111", -- 2893 - 0xb4d  :  127 - 0x7f
    "01111111", -- 2894 - 0xb4e  :  127 - 0x7f
    "01111111", -- 2895 - 0xb4f  :  127 - 0x7f
    "11011110", -- 2896 - 0xb50  :  222 - 0xde -- Background 0xb5
    "01100001", -- 2897 - 0xb51  :   97 - 0x61
    "01100001", -- 2898 - 0xb52  :   97 - 0x61
    "01100001", -- 2899 - 0xb53  :   97 - 0x61
    "01110001", -- 2900 - 0xb54  :  113 - 0x71
    "01011110", -- 2901 - 0xb55  :   94 - 0x5e
    "01111111", -- 2902 - 0xb56  :  127 - 0x7f
    "01100001", -- 2903 - 0xb57  :   97 - 0x61
    "01100001", -- 2904 - 0xb58  :   97 - 0x61 -- plane 1
    "11011111", -- 2905 - 0xb59  :  223 - 0xdf
    "11011111", -- 2906 - 0xb5a  :  223 - 0xdf
    "11011111", -- 2907 - 0xb5b  :  223 - 0xdf
    "11011111", -- 2908 - 0xb5c  :  223 - 0xdf
    "11111111", -- 2909 - 0xb5d  :  255 - 0xff
    "11000001", -- 2910 - 0xb5e  :  193 - 0xc1
    "11011111", -- 2911 - 0xb5f  :  223 - 0xdf
    "10000000", -- 2912 - 0xb60  :  128 - 0x80 -- Background 0xb6
    "10000000", -- 2913 - 0xb61  :  128 - 0x80
    "11000000", -- 2914 - 0xb62  :  192 - 0xc0
    "11110000", -- 2915 - 0xb63  :  240 - 0xf0
    "10111111", -- 2916 - 0xb64  :  191 - 0xbf
    "10001111", -- 2917 - 0xb65  :  143 - 0x8f
    "10000001", -- 2918 - 0xb66  :  129 - 0x81
    "01111110", -- 2919 - 0xb67  :  126 - 0x7e
    "01111111", -- 2920 - 0xb68  :  127 - 0x7f -- plane 1
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "11111111", -- 2922 - 0xb6a  :  255 - 0xff
    "00111111", -- 2923 - 0xb6b  :   63 - 0x3f
    "01001111", -- 2924 - 0xb6c  :   79 - 0x4f
    "01110001", -- 2925 - 0xb6d  :  113 - 0x71
    "01111111", -- 2926 - 0xb6e  :  127 - 0x7f
    "11111111", -- 2927 - 0xb6f  :  255 - 0xff
    "01100001", -- 2928 - 0xb70  :   97 - 0x61 -- Background 0xb7
    "01100001", -- 2929 - 0xb71  :   97 - 0x61
    "11000001", -- 2930 - 0xb72  :  193 - 0xc1
    "11000001", -- 2931 - 0xb73  :  193 - 0xc1
    "10000001", -- 2932 - 0xb74  :  129 - 0x81
    "10000001", -- 2933 - 0xb75  :  129 - 0x81
    "10000011", -- 2934 - 0xb76  :  131 - 0x83
    "11111110", -- 2935 - 0xb77  :  254 - 0xfe
    "11011111", -- 2936 - 0xb78  :  223 - 0xdf -- plane 1
    "11011111", -- 2937 - 0xb79  :  223 - 0xdf
    "10111111", -- 2938 - 0xb7a  :  191 - 0xbf
    "10111111", -- 2939 - 0xb7b  :  191 - 0xbf
    "01111111", -- 2940 - 0xb7c  :  127 - 0x7f
    "01111111", -- 2941 - 0xb7d  :  127 - 0x7f
    "01111111", -- 2942 - 0xb7e  :  127 - 0x7f
    "01111111", -- 2943 - 0xb7f  :  127 - 0x7f
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000011", -- 2946 - 0xb82  :    3 - 0x3
    "00001111", -- 2947 - 0xb83  :   15 - 0xf
    "00011111", -- 2948 - 0xb84  :   31 - 0x1f
    "00111111", -- 2949 - 0xb85  :   63 - 0x3f
    "01111111", -- 2950 - 0xb86  :  127 - 0x7f
    "01111111", -- 2951 - 0xb87  :  127 - 0x7f
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- plane 1
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000011", -- 2954 - 0xb8a  :    3 - 0x3
    "00001100", -- 2955 - 0xb8b  :   12 - 0xc
    "00010000", -- 2956 - 0xb8c  :   16 - 0x10
    "00100000", -- 2957 - 0xb8d  :   32 - 0x20
    "01000000", -- 2958 - 0xb8e  :   64 - 0x40
    "01000000", -- 2959 - 0xb8f  :   64 - 0x40
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Background 0xb9
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "11000000", -- 2962 - 0xb92  :  192 - 0xc0
    "11110000", -- 2963 - 0xb93  :  240 - 0xf0
    "11111000", -- 2964 - 0xb94  :  248 - 0xf8
    "11111100", -- 2965 - 0xb95  :  252 - 0xfc
    "11111110", -- 2966 - 0xb96  :  254 - 0xfe
    "11111110", -- 2967 - 0xb97  :  254 - 0xfe
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- plane 1
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "11000000", -- 2970 - 0xb9a  :  192 - 0xc0
    "00110000", -- 2971 - 0xb9b  :   48 - 0x30
    "00001000", -- 2972 - 0xb9c  :    8 - 0x8
    "00000100", -- 2973 - 0xb9d  :    4 - 0x4
    "00000010", -- 2974 - 0xb9e  :    2 - 0x2
    "00000010", -- 2975 - 0xb9f  :    2 - 0x2
    "11111111", -- 2976 - 0xba0  :  255 - 0xff -- Background 0xba
    "11111111", -- 2977 - 0xba1  :  255 - 0xff
    "11111111", -- 2978 - 0xba2  :  255 - 0xff
    "11111111", -- 2979 - 0xba3  :  255 - 0xff
    "11111111", -- 2980 - 0xba4  :  255 - 0xff
    "11111111", -- 2981 - 0xba5  :  255 - 0xff
    "11111111", -- 2982 - 0xba6  :  255 - 0xff
    "11111111", -- 2983 - 0xba7  :  255 - 0xff
    "10000000", -- 2984 - 0xba8  :  128 - 0x80 -- plane 1
    "10000000", -- 2985 - 0xba9  :  128 - 0x80
    "10000000", -- 2986 - 0xbaa  :  128 - 0x80
    "10000000", -- 2987 - 0xbab  :  128 - 0x80
    "10000000", -- 2988 - 0xbac  :  128 - 0x80
    "10000000", -- 2989 - 0xbad  :  128 - 0x80
    "10000000", -- 2990 - 0xbae  :  128 - 0x80
    "10000000", -- 2991 - 0xbaf  :  128 - 0x80
    "11111111", -- 2992 - 0xbb0  :  255 - 0xff -- Background 0xbb
    "11111111", -- 2993 - 0xbb1  :  255 - 0xff
    "11111111", -- 2994 - 0xbb2  :  255 - 0xff
    "11111111", -- 2995 - 0xbb3  :  255 - 0xff
    "11111111", -- 2996 - 0xbb4  :  255 - 0xff
    "11111111", -- 2997 - 0xbb5  :  255 - 0xff
    "11111111", -- 2998 - 0xbb6  :  255 - 0xff
    "11111111", -- 2999 - 0xbb7  :  255 - 0xff
    "00000001", -- 3000 - 0xbb8  :    1 - 0x1 -- plane 1
    "00000001", -- 3001 - 0xbb9  :    1 - 0x1
    "00000001", -- 3002 - 0xbba  :    1 - 0x1
    "00000001", -- 3003 - 0xbbb  :    1 - 0x1
    "00000001", -- 3004 - 0xbbc  :    1 - 0x1
    "00000001", -- 3005 - 0xbbd  :    1 - 0x1
    "00000001", -- 3006 - 0xbbe  :    1 - 0x1
    "00000001", -- 3007 - 0xbbf  :    1 - 0x1
    "01111111", -- 3008 - 0xbc0  :  127 - 0x7f -- Background 0xbc
    "01111111", -- 3009 - 0xbc1  :  127 - 0x7f
    "01111111", -- 3010 - 0xbc2  :  127 - 0x7f
    "00111111", -- 3011 - 0xbc3  :   63 - 0x3f
    "00111111", -- 3012 - 0xbc4  :   63 - 0x3f
    "00011111", -- 3013 - 0xbc5  :   31 - 0x1f
    "00001111", -- 3014 - 0xbc6  :   15 - 0xf
    "00000111", -- 3015 - 0xbc7  :    7 - 0x7
    "01000000", -- 3016 - 0xbc8  :   64 - 0x40 -- plane 1
    "01000000", -- 3017 - 0xbc9  :   64 - 0x40
    "01000000", -- 3018 - 0xbca  :   64 - 0x40
    "00100000", -- 3019 - 0xbcb  :   32 - 0x20
    "00110000", -- 3020 - 0xbcc  :   48 - 0x30
    "00011100", -- 3021 - 0xbcd  :   28 - 0x1c
    "00001111", -- 3022 - 0xbce  :   15 - 0xf
    "00000111", -- 3023 - 0xbcf  :    7 - 0x7
    "11111110", -- 3024 - 0xbd0  :  254 - 0xfe -- Background 0xbd
    "11111110", -- 3025 - 0xbd1  :  254 - 0xfe
    "11111110", -- 3026 - 0xbd2  :  254 - 0xfe
    "11111100", -- 3027 - 0xbd3  :  252 - 0xfc
    "11111100", -- 3028 - 0xbd4  :  252 - 0xfc
    "11111000", -- 3029 - 0xbd5  :  248 - 0xf8
    "11110000", -- 3030 - 0xbd6  :  240 - 0xf0
    "11110000", -- 3031 - 0xbd7  :  240 - 0xf0
    "00000010", -- 3032 - 0xbd8  :    2 - 0x2 -- plane 1
    "00000010", -- 3033 - 0xbd9  :    2 - 0x2
    "00000010", -- 3034 - 0xbda  :    2 - 0x2
    "00000100", -- 3035 - 0xbdb  :    4 - 0x4
    "00001100", -- 3036 - 0xbdc  :   12 - 0xc
    "00111000", -- 3037 - 0xbdd  :   56 - 0x38
    "11110000", -- 3038 - 0xbde  :  240 - 0xf0
    "11110000", -- 3039 - 0xbdf  :  240 - 0xf0
    "00001111", -- 3040 - 0xbe0  :   15 - 0xf -- Background 0xbe
    "00001111", -- 3041 - 0xbe1  :   15 - 0xf
    "00001111", -- 3042 - 0xbe2  :   15 - 0xf
    "00001111", -- 3043 - 0xbe3  :   15 - 0xf
    "00001111", -- 3044 - 0xbe4  :   15 - 0xf
    "00001111", -- 3045 - 0xbe5  :   15 - 0xf
    "00000111", -- 3046 - 0xbe6  :    7 - 0x7
    "00001111", -- 3047 - 0xbe7  :   15 - 0xf
    "00001000", -- 3048 - 0xbe8  :    8 - 0x8 -- plane 1
    "00001000", -- 3049 - 0xbe9  :    8 - 0x8
    "00001000", -- 3050 - 0xbea  :    8 - 0x8
    "00001000", -- 3051 - 0xbeb  :    8 - 0x8
    "00001000", -- 3052 - 0xbec  :    8 - 0x8
    "00001100", -- 3053 - 0xbed  :   12 - 0xc
    "00000101", -- 3054 - 0xbee  :    5 - 0x5
    "00001010", -- 3055 - 0xbef  :   10 - 0xa
    "11110000", -- 3056 - 0xbf0  :  240 - 0xf0 -- Background 0xbf
    "11110000", -- 3057 - 0xbf1  :  240 - 0xf0
    "11110000", -- 3058 - 0xbf2  :  240 - 0xf0
    "11110000", -- 3059 - 0xbf3  :  240 - 0xf0
    "11110000", -- 3060 - 0xbf4  :  240 - 0xf0
    "11110000", -- 3061 - 0xbf5  :  240 - 0xf0
    "11100000", -- 3062 - 0xbf6  :  224 - 0xe0
    "11110000", -- 3063 - 0xbf7  :  240 - 0xf0
    "00010000", -- 3064 - 0xbf8  :   16 - 0x10 -- plane 1
    "01010000", -- 3065 - 0xbf9  :   80 - 0x50
    "01010000", -- 3066 - 0xbfa  :   80 - 0x50
    "01010000", -- 3067 - 0xbfb  :   80 - 0x50
    "01010000", -- 3068 - 0xbfc  :   80 - 0x50
    "00110000", -- 3069 - 0xbfd  :   48 - 0x30
    "10100000", -- 3070 - 0xbfe  :  160 - 0xa0
    "01010000", -- 3071 - 0xbff  :   80 - 0x50
    "10000001", -- 3072 - 0xc00  :  129 - 0x81 -- Background 0xc0
    "11000001", -- 3073 - 0xc01  :  193 - 0xc1
    "10100011", -- 3074 - 0xc02  :  163 - 0xa3
    "10100011", -- 3075 - 0xc03  :  163 - 0xa3
    "10011101", -- 3076 - 0xc04  :  157 - 0x9d
    "10000001", -- 3077 - 0xc05  :  129 - 0x81
    "10000001", -- 3078 - 0xc06  :  129 - 0x81
    "10000001", -- 3079 - 0xc07  :  129 - 0x81
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- plane 1
    "01000001", -- 3081 - 0xc09  :   65 - 0x41
    "00100010", -- 3082 - 0xc0a  :   34 - 0x22
    "00100010", -- 3083 - 0xc0b  :   34 - 0x22
    "00011100", -- 3084 - 0xc0c  :   28 - 0x1c
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "11100011", -- 3088 - 0xc10  :  227 - 0xe3 -- Background 0xc1
    "11110111", -- 3089 - 0xc11  :  247 - 0xf7
    "11000001", -- 3090 - 0xc12  :  193 - 0xc1
    "11000001", -- 3091 - 0xc13  :  193 - 0xc1
    "11000001", -- 3092 - 0xc14  :  193 - 0xc1
    "11000001", -- 3093 - 0xc15  :  193 - 0xc1
    "11110111", -- 3094 - 0xc16  :  247 - 0xf7
    "11100011", -- 3095 - 0xc17  :  227 - 0xe3
    "11100011", -- 3096 - 0xc18  :  227 - 0xe3 -- plane 1
    "00010100", -- 3097 - 0xc19  :   20 - 0x14
    "00111110", -- 3098 - 0xc1a  :   62 - 0x3e
    "00111110", -- 3099 - 0xc1b  :   62 - 0x3e
    "00111110", -- 3100 - 0xc1c  :   62 - 0x3e
    "00111110", -- 3101 - 0xc1d  :   62 - 0x3e
    "00010100", -- 3102 - 0xc1e  :   20 - 0x14
    "11100011", -- 3103 - 0xc1f  :  227 - 0xe3
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000111", -- 3106 - 0xc22  :    7 - 0x7
    "00001111", -- 3107 - 0xc23  :   15 - 0xf
    "00001100", -- 3108 - 0xc24  :   12 - 0xc
    "00011011", -- 3109 - 0xc25  :   27 - 0x1b
    "00011011", -- 3110 - 0xc26  :   27 - 0x1b
    "00011011", -- 3111 - 0xc27  :   27 - 0x1b
    "11111111", -- 3112 - 0xc28  :  255 - 0xff -- plane 1
    "11111111", -- 3113 - 0xc29  :  255 - 0xff
    "11111000", -- 3114 - 0xc2a  :  248 - 0xf8
    "11110000", -- 3115 - 0xc2b  :  240 - 0xf0
    "11110000", -- 3116 - 0xc2c  :  240 - 0xf0
    "11100000", -- 3117 - 0xc2d  :  224 - 0xe0
    "11100000", -- 3118 - 0xc2e  :  224 - 0xe0
    "11100000", -- 3119 - 0xc2f  :  224 - 0xe0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "11100000", -- 3122 - 0xc32  :  224 - 0xe0
    "11110000", -- 3123 - 0xc33  :  240 - 0xf0
    "11110000", -- 3124 - 0xc34  :  240 - 0xf0
    "11111000", -- 3125 - 0xc35  :  248 - 0xf8
    "11111000", -- 3126 - 0xc36  :  248 - 0xf8
    "11111000", -- 3127 - 0xc37  :  248 - 0xf8
    "11111111", -- 3128 - 0xc38  :  255 - 0xff -- plane 1
    "11111111", -- 3129 - 0xc39  :  255 - 0xff
    "01111111", -- 3130 - 0xc3a  :  127 - 0x7f
    "00111111", -- 3131 - 0xc3b  :   63 - 0x3f
    "00111111", -- 3132 - 0xc3c  :   63 - 0x3f
    "10011111", -- 3133 - 0xc3d  :  159 - 0x9f
    "10011111", -- 3134 - 0xc3e  :  159 - 0x9f
    "10011111", -- 3135 - 0xc3f  :  159 - 0x9f
    "00011011", -- 3136 - 0xc40  :   27 - 0x1b -- Background 0xc4
    "00011011", -- 3137 - 0xc41  :   27 - 0x1b
    "00011011", -- 3138 - 0xc42  :   27 - 0x1b
    "00011011", -- 3139 - 0xc43  :   27 - 0x1b
    "00011011", -- 3140 - 0xc44  :   27 - 0x1b
    "00001111", -- 3141 - 0xc45  :   15 - 0xf
    "00001111", -- 3142 - 0xc46  :   15 - 0xf
    "00000111", -- 3143 - 0xc47  :    7 - 0x7
    "11100000", -- 3144 - 0xc48  :  224 - 0xe0 -- plane 1
    "11100000", -- 3145 - 0xc49  :  224 - 0xe0
    "11100000", -- 3146 - 0xc4a  :  224 - 0xe0
    "11100000", -- 3147 - 0xc4b  :  224 - 0xe0
    "11100000", -- 3148 - 0xc4c  :  224 - 0xe0
    "11110011", -- 3149 - 0xc4d  :  243 - 0xf3
    "11110000", -- 3150 - 0xc4e  :  240 - 0xf0
    "11111000", -- 3151 - 0xc4f  :  248 - 0xf8
    "11111000", -- 3152 - 0xc50  :  248 - 0xf8 -- Background 0xc5
    "11111000", -- 3153 - 0xc51  :  248 - 0xf8
    "11111000", -- 3154 - 0xc52  :  248 - 0xf8
    "11111000", -- 3155 - 0xc53  :  248 - 0xf8
    "11111000", -- 3156 - 0xc54  :  248 - 0xf8
    "11110000", -- 3157 - 0xc55  :  240 - 0xf0
    "11110000", -- 3158 - 0xc56  :  240 - 0xf0
    "11100000", -- 3159 - 0xc57  :  224 - 0xe0
    "10011111", -- 3160 - 0xc58  :  159 - 0x9f -- plane 1
    "10011111", -- 3161 - 0xc59  :  159 - 0x9f
    "10011111", -- 3162 - 0xc5a  :  159 - 0x9f
    "10011111", -- 3163 - 0xc5b  :  159 - 0x9f
    "10011111", -- 3164 - 0xc5c  :  159 - 0x9f
    "00111111", -- 3165 - 0xc5d  :   63 - 0x3f
    "00111111", -- 3166 - 0xc5e  :   63 - 0x3f
    "01111111", -- 3167 - 0xc5f  :  127 - 0x7f
    "11100000", -- 3168 - 0xc60  :  224 - 0xe0 -- Background 0xc6
    "11111111", -- 3169 - 0xc61  :  255 - 0xff
    "11111111", -- 3170 - 0xc62  :  255 - 0xff
    "11111111", -- 3171 - 0xc63  :  255 - 0xff
    "11111111", -- 3172 - 0xc64  :  255 - 0xff
    "11111111", -- 3173 - 0xc65  :  255 - 0xff
    "11111111", -- 3174 - 0xc66  :  255 - 0xff
    "11111111", -- 3175 - 0xc67  :  255 - 0xff
    "00000000", -- 3176 - 0xc68  :    0 - 0x0 -- plane 1
    "01110000", -- 3177 - 0xc69  :  112 - 0x70
    "00011111", -- 3178 - 0xc6a  :   31 - 0x1f
    "00010000", -- 3179 - 0xc6b  :   16 - 0x10
    "01110000", -- 3180 - 0xc6c  :  112 - 0x70
    "01111111", -- 3181 - 0xc6d  :  127 - 0x7f
    "01111111", -- 3182 - 0xc6e  :  127 - 0x7f
    "01111111", -- 3183 - 0xc6f  :  127 - 0x7f
    "00000111", -- 3184 - 0xc70  :    7 - 0x7 -- Background 0xc7
    "11111111", -- 3185 - 0xc71  :  255 - 0xff
    "11111111", -- 3186 - 0xc72  :  255 - 0xff
    "11111111", -- 3187 - 0xc73  :  255 - 0xff
    "11111111", -- 3188 - 0xc74  :  255 - 0xff
    "11111111", -- 3189 - 0xc75  :  255 - 0xff
    "11111111", -- 3190 - 0xc76  :  255 - 0xff
    "11111111", -- 3191 - 0xc77  :  255 - 0xff
    "00000000", -- 3192 - 0xc78  :    0 - 0x0 -- plane 1
    "00000011", -- 3193 - 0xc79  :    3 - 0x3
    "11111000", -- 3194 - 0xc7a  :  248 - 0xf8
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000011", -- 3196 - 0xc7c  :    3 - 0x3
    "11111011", -- 3197 - 0xc7d  :  251 - 0xfb
    "11111011", -- 3198 - 0xc7e  :  251 - 0xfb
    "11111011", -- 3199 - 0xc7f  :  251 - 0xfb
    "11111111", -- 3200 - 0xc80  :  255 - 0xff -- Background 0xc8
    "11111111", -- 3201 - 0xc81  :  255 - 0xff
    "11111111", -- 3202 - 0xc82  :  255 - 0xff
    "11111111", -- 3203 - 0xc83  :  255 - 0xff
    "11111111", -- 3204 - 0xc84  :  255 - 0xff
    "11111110", -- 3205 - 0xc85  :  254 - 0xfe
    "11111111", -- 3206 - 0xc86  :  255 - 0xff
    "11101111", -- 3207 - 0xc87  :  239 - 0xef
    "01111100", -- 3208 - 0xc88  :  124 - 0x7c -- plane 1
    "01111011", -- 3209 - 0xc89  :  123 - 0x7b
    "01110110", -- 3210 - 0xc8a  :  118 - 0x76
    "01110101", -- 3211 - 0xc8b  :  117 - 0x75
    "01110101", -- 3212 - 0xc8c  :  117 - 0x75
    "01110111", -- 3213 - 0xc8d  :  119 - 0x77
    "00010111", -- 3214 - 0xc8e  :   23 - 0x17
    "01100111", -- 3215 - 0xc8f  :  103 - 0x67
    "11111111", -- 3216 - 0xc90  :  255 - 0xff -- Background 0xc9
    "11011111", -- 3217 - 0xc91  :  223 - 0xdf
    "11101111", -- 3218 - 0xc92  :  239 - 0xef
    "10101111", -- 3219 - 0xc93  :  175 - 0xaf
    "10101111", -- 3220 - 0xc94  :  175 - 0xaf
    "01101111", -- 3221 - 0xc95  :  111 - 0x6f
    "11101111", -- 3222 - 0xc96  :  239 - 0xef
    "11100111", -- 3223 - 0xc97  :  231 - 0xe7
    "00111011", -- 3224 - 0xc98  :   59 - 0x3b -- plane 1
    "11111011", -- 3225 - 0xc99  :  251 - 0xfb
    "01111011", -- 3226 - 0xc9a  :  123 - 0x7b
    "11111011", -- 3227 - 0xc9b  :  251 - 0xfb
    "11111011", -- 3228 - 0xc9c  :  251 - 0xfb
    "11110011", -- 3229 - 0xc9d  :  243 - 0xf3
    "11111000", -- 3230 - 0xc9e  :  248 - 0xf8
    "11110011", -- 3231 - 0xc9f  :  243 - 0xf3
    "00011111", -- 3232 - 0xca0  :   31 - 0x1f -- Background 0xca
    "00011111", -- 3233 - 0xca1  :   31 - 0x1f
    "00111111", -- 3234 - 0xca2  :   63 - 0x3f
    "00111111", -- 3235 - 0xca3  :   63 - 0x3f
    "01110000", -- 3236 - 0xca4  :  112 - 0x70
    "01100011", -- 3237 - 0xca5  :   99 - 0x63
    "11100111", -- 3238 - 0xca6  :  231 - 0xe7
    "11100101", -- 3239 - 0xca7  :  229 - 0xe5
    "00001111", -- 3240 - 0xca8  :   15 - 0xf -- plane 1
    "00001111", -- 3241 - 0xca9  :   15 - 0xf
    "00011111", -- 3242 - 0xcaa  :   31 - 0x1f
    "00011111", -- 3243 - 0xcab  :   31 - 0x1f
    "00111111", -- 3244 - 0xcac  :   63 - 0x3f
    "00111100", -- 3245 - 0xcad  :   60 - 0x3c
    "01111000", -- 3246 - 0xcae  :  120 - 0x78
    "01111010", -- 3247 - 0xcaf  :  122 - 0x7a
    "11110000", -- 3248 - 0xcb0  :  240 - 0xf0 -- Background 0xcb
    "11110000", -- 3249 - 0xcb1  :  240 - 0xf0
    "11111000", -- 3250 - 0xcb2  :  248 - 0xf8
    "11111000", -- 3251 - 0xcb3  :  248 - 0xf8
    "00001100", -- 3252 - 0xcb4  :   12 - 0xc
    "11000100", -- 3253 - 0xcb5  :  196 - 0xc4
    "11100100", -- 3254 - 0xcb6  :  228 - 0xe4
    "10100110", -- 3255 - 0xcb7  :  166 - 0xa6
    "11111000", -- 3256 - 0xcb8  :  248 - 0xf8 -- plane 1
    "11111000", -- 3257 - 0xcb9  :  248 - 0xf8
    "11111100", -- 3258 - 0xcba  :  252 - 0xfc
    "11111100", -- 3259 - 0xcbb  :  252 - 0xfc
    "11111110", -- 3260 - 0xcbc  :  254 - 0xfe
    "00111110", -- 3261 - 0xcbd  :   62 - 0x3e
    "00011110", -- 3262 - 0xcbe  :   30 - 0x1e
    "01011111", -- 3263 - 0xcbf  :   95 - 0x5f
    "11101001", -- 3264 - 0xcc0  :  233 - 0xe9 -- Background 0xcc
    "11101001", -- 3265 - 0xcc1  :  233 - 0xe9
    "11101001", -- 3266 - 0xcc2  :  233 - 0xe9
    "11101111", -- 3267 - 0xcc3  :  239 - 0xef
    "11100010", -- 3268 - 0xcc4  :  226 - 0xe2
    "11100011", -- 3269 - 0xcc5  :  227 - 0xe3
    "11110000", -- 3270 - 0xcc6  :  240 - 0xf0
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "01110110", -- 3272 - 0xcc8  :  118 - 0x76 -- plane 1
    "01110110", -- 3273 - 0xcc9  :  118 - 0x76
    "01110110", -- 3274 - 0xcca  :  118 - 0x76
    "01110000", -- 3275 - 0xccb  :  112 - 0x70
    "01111101", -- 3276 - 0xccc  :  125 - 0x7d
    "01111100", -- 3277 - 0xccd  :  124 - 0x7c
    "01111111", -- 3278 - 0xcce  :  127 - 0x7f
    "01111111", -- 3279 - 0xccf  :  127 - 0x7f
    "10010110", -- 3280 - 0xcd0  :  150 - 0x96 -- Background 0xcd
    "10010110", -- 3281 - 0xcd1  :  150 - 0x96
    "10010110", -- 3282 - 0xcd2  :  150 - 0x96
    "11110110", -- 3283 - 0xcd3  :  246 - 0xf6
    "01000110", -- 3284 - 0xcd4  :   70 - 0x46
    "11000110", -- 3285 - 0xcd5  :  198 - 0xc6
    "00001110", -- 3286 - 0xcd6  :   14 - 0xe
    "11111110", -- 3287 - 0xcd7  :  254 - 0xfe
    "01101111", -- 3288 - 0xcd8  :  111 - 0x6f -- plane 1
    "01101111", -- 3289 - 0xcd9  :  111 - 0x6f
    "01101111", -- 3290 - 0xcda  :  111 - 0x6f
    "00001111", -- 3291 - 0xcdb  :   15 - 0xf
    "10111111", -- 3292 - 0xcdc  :  191 - 0xbf
    "00111111", -- 3293 - 0xcdd  :   63 - 0x3f
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "01111110", -- 3302 - 0xce6  :  126 - 0x7e
    "00111100", -- 3303 - 0xce7  :   60 - 0x3c
    "00111100", -- 3304 - 0xce8  :   60 - 0x3c -- plane 1
    "01111110", -- 3305 - 0xce9  :  126 - 0x7e
    "01111110", -- 3306 - 0xcea  :  126 - 0x7e
    "11111111", -- 3307 - 0xceb  :  255 - 0xff
    "11111111", -- 3308 - 0xcec  :  255 - 0xff
    "11111111", -- 3309 - 0xced  :  255 - 0xff
    "01000010", -- 3310 - 0xcee  :   66 - 0x42
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00111100", -- 3312 - 0xcf0  :   60 - 0x3c -- Background 0xcf
    "01000010", -- 3313 - 0xcf1  :   66 - 0x42
    "10011001", -- 3314 - 0xcf2  :  153 - 0x99
    "10100001", -- 3315 - 0xcf3  :  161 - 0xa1
    "10100001", -- 3316 - 0xcf4  :  161 - 0xa1
    "10011001", -- 3317 - 0xcf5  :  153 - 0x99
    "01000010", -- 3318 - 0xcf6  :   66 - 0x42
    "00111100", -- 3319 - 0xcf7  :   60 - 0x3c
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00001111", -- 3328 - 0xd00  :   15 - 0xf -- Background 0xd0
    "00011111", -- 3329 - 0xd01  :   31 - 0x1f
    "00011111", -- 3330 - 0xd02  :   31 - 0x1f
    "00111111", -- 3331 - 0xd03  :   63 - 0x3f
    "00111111", -- 3332 - 0xd04  :   63 - 0x3f
    "01111111", -- 3333 - 0xd05  :  127 - 0x7f
    "01111111", -- 3334 - 0xd06  :  127 - 0x7f
    "01111111", -- 3335 - 0xd07  :  127 - 0x7f
    "11110000", -- 3336 - 0xd08  :  240 - 0xf0 -- plane 1
    "11100000", -- 3337 - 0xd09  :  224 - 0xe0
    "11100000", -- 3338 - 0xd0a  :  224 - 0xe0
    "11000000", -- 3339 - 0xd0b  :  192 - 0xc0
    "11000000", -- 3340 - 0xd0c  :  192 - 0xc0
    "10000000", -- 3341 - 0xd0d  :  128 - 0x80
    "10000000", -- 3342 - 0xd0e  :  128 - 0x80
    "10000000", -- 3343 - 0xd0f  :  128 - 0x80
    "11110000", -- 3344 - 0xd10  :  240 - 0xf0 -- Background 0xd1
    "11111000", -- 3345 - 0xd11  :  248 - 0xf8
    "11111000", -- 3346 - 0xd12  :  248 - 0xf8
    "11111100", -- 3347 - 0xd13  :  252 - 0xfc
    "11111100", -- 3348 - 0xd14  :  252 - 0xfc
    "11111110", -- 3349 - 0xd15  :  254 - 0xfe
    "11111110", -- 3350 - 0xd16  :  254 - 0xfe
    "11111110", -- 3351 - 0xd17  :  254 - 0xfe
    "00001111", -- 3352 - 0xd18  :   15 - 0xf -- plane 1
    "00000111", -- 3353 - 0xd19  :    7 - 0x7
    "00000111", -- 3354 - 0xd1a  :    7 - 0x7
    "00000011", -- 3355 - 0xd1b  :    3 - 0x3
    "00000011", -- 3356 - 0xd1c  :    3 - 0x3
    "00000001", -- 3357 - 0xd1d  :    1 - 0x1
    "00000001", -- 3358 - 0xd1e  :    1 - 0x1
    "00000001", -- 3359 - 0xd1f  :    1 - 0x1
    "01111111", -- 3360 - 0xd20  :  127 - 0x7f -- Background 0xd2
    "01111111", -- 3361 - 0xd21  :  127 - 0x7f
    "00111111", -- 3362 - 0xd22  :   63 - 0x3f
    "00111111", -- 3363 - 0xd23  :   63 - 0x3f
    "00111111", -- 3364 - 0xd24  :   63 - 0x3f
    "00111111", -- 3365 - 0xd25  :   63 - 0x3f
    "00011111", -- 3366 - 0xd26  :   31 - 0x1f
    "00011111", -- 3367 - 0xd27  :   31 - 0x1f
    "10000000", -- 3368 - 0xd28  :  128 - 0x80 -- plane 1
    "10000000", -- 3369 - 0xd29  :  128 - 0x80
    "11000000", -- 3370 - 0xd2a  :  192 - 0xc0
    "11000000", -- 3371 - 0xd2b  :  192 - 0xc0
    "11100000", -- 3372 - 0xd2c  :  224 - 0xe0
    "11111000", -- 3373 - 0xd2d  :  248 - 0xf8
    "11111110", -- 3374 - 0xd2e  :  254 - 0xfe
    "11111111", -- 3375 - 0xd2f  :  255 - 0xff
    "11111110", -- 3376 - 0xd30  :  254 - 0xfe -- Background 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11111100", -- 3380 - 0xd34  :  252 - 0xfc
    "11111100", -- 3381 - 0xd35  :  252 - 0xfc
    "11111110", -- 3382 - 0xd36  :  254 - 0xfe
    "11111110", -- 3383 - 0xd37  :  254 - 0xfe
    "11111111", -- 3384 - 0xd38  :  255 - 0xff -- plane 1
    "01111111", -- 3385 - 0xd39  :  127 - 0x7f
    "00011111", -- 3386 - 0xd3a  :   31 - 0x1f
    "00000111", -- 3387 - 0xd3b  :    7 - 0x7
    "00000011", -- 3388 - 0xd3c  :    3 - 0x3
    "00000011", -- 3389 - 0xd3d  :    3 - 0x3
    "00000001", -- 3390 - 0xd3e  :    1 - 0x1
    "10000001", -- 3391 - 0xd3f  :  129 - 0x81
    "01111111", -- 3392 - 0xd40  :  127 - 0x7f -- Background 0xd4
    "01111111", -- 3393 - 0xd41  :  127 - 0x7f
    "01111111", -- 3394 - 0xd42  :  127 - 0x7f
    "00111111", -- 3395 - 0xd43  :   63 - 0x3f
    "00111111", -- 3396 - 0xd44  :   63 - 0x3f
    "00111111", -- 3397 - 0xd45  :   63 - 0x3f
    "00111111", -- 3398 - 0xd46  :   63 - 0x3f
    "00011111", -- 3399 - 0xd47  :   31 - 0x1f
    "10000000", -- 3400 - 0xd48  :  128 - 0x80 -- plane 1
    "10000000", -- 3401 - 0xd49  :  128 - 0x80
    "10000000", -- 3402 - 0xd4a  :  128 - 0x80
    "11000000", -- 3403 - 0xd4b  :  192 - 0xc0
    "11000000", -- 3404 - 0xd4c  :  192 - 0xc0
    "11100000", -- 3405 - 0xd4d  :  224 - 0xe0
    "11100000", -- 3406 - 0xd4e  :  224 - 0xe0
    "11110000", -- 3407 - 0xd4f  :  240 - 0xf0
    "11111110", -- 3408 - 0xd50  :  254 - 0xfe -- Background 0xd5
    "11111110", -- 3409 - 0xd51  :  254 - 0xfe
    "11111111", -- 3410 - 0xd52  :  255 - 0xff
    "11111111", -- 3411 - 0xd53  :  255 - 0xff
    "11111111", -- 3412 - 0xd54  :  255 - 0xff
    "11111111", -- 3413 - 0xd55  :  255 - 0xff
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111110", -- 3415 - 0xd57  :  254 - 0xfe
    "00000001", -- 3416 - 0xd58  :    1 - 0x1 -- plane 1
    "00000001", -- 3417 - 0xd59  :    1 - 0x1
    "00000001", -- 3418 - 0xd5a  :    1 - 0x1
    "00000011", -- 3419 - 0xd5b  :    3 - 0x3
    "00000011", -- 3420 - 0xd5c  :    3 - 0x3
    "00000111", -- 3421 - 0xd5d  :    7 - 0x7
    "00000111", -- 3422 - 0xd5e  :    7 - 0x7
    "00001111", -- 3423 - 0xd5f  :   15 - 0xf
    "00011111", -- 3424 - 0xd60  :   31 - 0x1f -- Background 0xd6
    "00001111", -- 3425 - 0xd61  :   15 - 0xf
    "00001111", -- 3426 - 0xd62  :   15 - 0xf
    "00000111", -- 3427 - 0xd63  :    7 - 0x7
    "00000000", -- 3428 - 0xd64  :    0 - 0x0
    "00000000", -- 3429 - 0xd65  :    0 - 0x0
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "00000000", -- 3431 - 0xd67  :    0 - 0x0
    "11111111", -- 3432 - 0xd68  :  255 - 0xff -- plane 1
    "11111111", -- 3433 - 0xd69  :  255 - 0xff
    "11111111", -- 3434 - 0xd6a  :  255 - 0xff
    "11111111", -- 3435 - 0xd6b  :  255 - 0xff
    "11111111", -- 3436 - 0xd6c  :  255 - 0xff
    "11111111", -- 3437 - 0xd6d  :  255 - 0xff
    "11111111", -- 3438 - 0xd6e  :  255 - 0xff
    "11111111", -- 3439 - 0xd6f  :  255 - 0xff
    "11111110", -- 3440 - 0xd70  :  254 - 0xfe -- Background 0xd7
    "11111100", -- 3441 - 0xd71  :  252 - 0xfc
    "11111100", -- 3442 - 0xd72  :  252 - 0xfc
    "11111000", -- 3443 - 0xd73  :  248 - 0xf8
    "00000000", -- 3444 - 0xd74  :    0 - 0x0
    "00000000", -- 3445 - 0xd75  :    0 - 0x0
    "00000000", -- 3446 - 0xd76  :    0 - 0x0
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "11111111", -- 3448 - 0xd78  :  255 - 0xff -- plane 1
    "11111111", -- 3449 - 0xd79  :  255 - 0xff
    "11111111", -- 3450 - 0xd7a  :  255 - 0xff
    "11111111", -- 3451 - 0xd7b  :  255 - 0xff
    "11111111", -- 3452 - 0xd7c  :  255 - 0xff
    "11111111", -- 3453 - 0xd7d  :  255 - 0xff
    "11111111", -- 3454 - 0xd7e  :  255 - 0xff
    "11111111", -- 3455 - 0xd7f  :  255 - 0xff
    "01111110", -- 3456 - 0xd80  :  126 - 0x7e -- Background 0xd8
    "01111110", -- 3457 - 0xd81  :  126 - 0x7e
    "01111110", -- 3458 - 0xd82  :  126 - 0x7e
    "01111110", -- 3459 - 0xd83  :  126 - 0x7e
    "01111111", -- 3460 - 0xd84  :  127 - 0x7f
    "01111111", -- 3461 - 0xd85  :  127 - 0x7f
    "01111111", -- 3462 - 0xd86  :  127 - 0x7f
    "01111111", -- 3463 - 0xd87  :  127 - 0x7f
    "10000001", -- 3464 - 0xd88  :  129 - 0x81 -- plane 1
    "10000001", -- 3465 - 0xd89  :  129 - 0x81
    "10000001", -- 3466 - 0xd8a  :  129 - 0x81
    "10000001", -- 3467 - 0xd8b  :  129 - 0x81
    "10000001", -- 3468 - 0xd8c  :  129 - 0x81
    "10000001", -- 3469 - 0xd8d  :  129 - 0x81
    "10000001", -- 3470 - 0xd8e  :  129 - 0x81
    "10000001", -- 3471 - 0xd8f  :  129 - 0x81
    "11111111", -- 3472 - 0xd90  :  255 - 0xff -- Background 0xd9
    "11111111", -- 3473 - 0xd91  :  255 - 0xff
    "11111111", -- 3474 - 0xd92  :  255 - 0xff
    "11111111", -- 3475 - 0xd93  :  255 - 0xff
    "11111111", -- 3476 - 0xd94  :  255 - 0xff
    "11111111", -- 3477 - 0xd95  :  255 - 0xff
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111110", -- 3479 - 0xd97  :  254 - 0xfe
    "00000001", -- 3480 - 0xd98  :    1 - 0x1 -- plane 1
    "00000001", -- 3481 - 0xd99  :    1 - 0x1
    "00000001", -- 3482 - 0xd9a  :    1 - 0x1
    "00000011", -- 3483 - 0xd9b  :    3 - 0x3
    "00000011", -- 3484 - 0xd9c  :    3 - 0x3
    "00000111", -- 3485 - 0xd9d  :    7 - 0x7
    "00000111", -- 3486 - 0xd9e  :    7 - 0x7
    "00001111", -- 3487 - 0xd9f  :   15 - 0xf
    "11111110", -- 3488 - 0xda0  :  254 - 0xfe -- Background 0xda
    "11111110", -- 3489 - 0xda1  :  254 - 0xfe
    "11111110", -- 3490 - 0xda2  :  254 - 0xfe
    "11111110", -- 3491 - 0xda3  :  254 - 0xfe
    "11111111", -- 3492 - 0xda4  :  255 - 0xff
    "11111111", -- 3493 - 0xda5  :  255 - 0xff
    "11111111", -- 3494 - 0xda6  :  255 - 0xff
    "11111111", -- 3495 - 0xda7  :  255 - 0xff
    "00000001", -- 3496 - 0xda8  :    1 - 0x1 -- plane 1
    "00000001", -- 3497 - 0xda9  :    1 - 0x1
    "00000001", -- 3498 - 0xdaa  :    1 - 0x1
    "00000001", -- 3499 - 0xdab  :    1 - 0x1
    "00000001", -- 3500 - 0xdac  :    1 - 0x1
    "00000001", -- 3501 - 0xdad  :    1 - 0x1
    "00000001", -- 3502 - 0xdae  :    1 - 0x1
    "00000001", -- 3503 - 0xdaf  :    1 - 0x1
    "01111111", -- 3504 - 0xdb0  :  127 - 0x7f -- Background 0xdb
    "01111111", -- 3505 - 0xdb1  :  127 - 0x7f
    "01111111", -- 3506 - 0xdb2  :  127 - 0x7f
    "01111111", -- 3507 - 0xdb3  :  127 - 0x7f
    "01111111", -- 3508 - 0xdb4  :  127 - 0x7f
    "01111111", -- 3509 - 0xdb5  :  127 - 0x7f
    "01111111", -- 3510 - 0xdb6  :  127 - 0x7f
    "01111111", -- 3511 - 0xdb7  :  127 - 0x7f
    "10000001", -- 3512 - 0xdb8  :  129 - 0x81 -- plane 1
    "10000001", -- 3513 - 0xdb9  :  129 - 0x81
    "10000001", -- 3514 - 0xdba  :  129 - 0x81
    "10000001", -- 3515 - 0xdbb  :  129 - 0x81
    "10000001", -- 3516 - 0xdbc  :  129 - 0x81
    "10000001", -- 3517 - 0xdbd  :  129 - 0x81
    "10000001", -- 3518 - 0xdbe  :  129 - 0x81
    "10000001", -- 3519 - 0xdbf  :  129 - 0x81
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Background 0xdc
    "11111111", -- 3521 - 0xdc1  :  255 - 0xff
    "11111111", -- 3522 - 0xdc2  :  255 - 0xff
    "11111111", -- 3523 - 0xdc3  :  255 - 0xff
    "11111100", -- 3524 - 0xdc4  :  252 - 0xfc
    "11111110", -- 3525 - 0xdc5  :  254 - 0xfe
    "11111110", -- 3526 - 0xdc6  :  254 - 0xfe
    "01111110", -- 3527 - 0xdc7  :  126 - 0x7e
    "11111111", -- 3528 - 0xdc8  :  255 - 0xff -- plane 1
    "00000011", -- 3529 - 0xdc9  :    3 - 0x3
    "00000011", -- 3530 - 0xdca  :    3 - 0x3
    "00000011", -- 3531 - 0xdcb  :    3 - 0x3
    "00000011", -- 3532 - 0xdcc  :    3 - 0x3
    "00000011", -- 3533 - 0xdcd  :    3 - 0x3
    "00000011", -- 3534 - 0xdce  :    3 - 0x3
    "11111111", -- 3535 - 0xdcf  :  255 - 0xff
    "11111111", -- 3536 - 0xdd0  :  255 - 0xff -- Background 0xdd
    "11111111", -- 3537 - 0xdd1  :  255 - 0xff
    "11111111", -- 3538 - 0xdd2  :  255 - 0xff
    "11111111", -- 3539 - 0xdd3  :  255 - 0xff
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "00000000", -- 3541 - 0xdd5  :    0 - 0x0
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "11111111", -- 3544 - 0xdd8  :  255 - 0xff -- plane 1
    "11111111", -- 3545 - 0xdd9  :  255 - 0xff
    "11111111", -- 3546 - 0xdda  :  255 - 0xff
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "11111111", -- 3548 - 0xddc  :  255 - 0xff
    "11111111", -- 3549 - 0xddd  :  255 - 0xff
    "11111111", -- 3550 - 0xdde  :  255 - 0xff
    "11111111", -- 3551 - 0xddf  :  255 - 0xff
    "01111111", -- 3552 - 0xde0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 3553 - 0xde1  :  127 - 0x7f
    "01111111", -- 3554 - 0xde2  :  127 - 0x7f
    "01111111", -- 3555 - 0xde3  :  127 - 0x7f
    "01111111", -- 3556 - 0xde4  :  127 - 0x7f
    "01111111", -- 3557 - 0xde5  :  127 - 0x7f
    "01111111", -- 3558 - 0xde6  :  127 - 0x7f
    "01111111", -- 3559 - 0xde7  :  127 - 0x7f
    "10000000", -- 3560 - 0xde8  :  128 - 0x80 -- plane 1
    "10000000", -- 3561 - 0xde9  :  128 - 0x80
    "10000000", -- 3562 - 0xdea  :  128 - 0x80
    "10000000", -- 3563 - 0xdeb  :  128 - 0x80
    "10000000", -- 3564 - 0xdec  :  128 - 0x80
    "10000000", -- 3565 - 0xded  :  128 - 0x80
    "10000000", -- 3566 - 0xdee  :  128 - 0x80
    "10000000", -- 3567 - 0xdef  :  128 - 0x80
    "11111111", -- 3568 - 0xdf0  :  255 - 0xff -- Background 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "11111111", -- 3570 - 0xdf2  :  255 - 0xff
    "11111111", -- 3571 - 0xdf3  :  255 - 0xff
    "11111111", -- 3572 - 0xdf4  :  255 - 0xff
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111110", -- 3575 - 0xdf7  :  254 - 0xfe
    "00000001", -- 3576 - 0xdf8  :    1 - 0x1 -- plane 1
    "00000001", -- 3577 - 0xdf9  :    1 - 0x1
    "00000001", -- 3578 - 0xdfa  :    1 - 0x1
    "00000011", -- 3579 - 0xdfb  :    3 - 0x3
    "00000111", -- 3580 - 0xdfc  :    7 - 0x7
    "00000011", -- 3581 - 0xdfd  :    3 - 0x3
    "00000001", -- 3582 - 0xdfe  :    1 - 0x1
    "00000001", -- 3583 - 0xdff  :    1 - 0x1
    "01111110", -- 3584 - 0xe00  :  126 - 0x7e -- Background 0xe0
    "01111110", -- 3585 - 0xe01  :  126 - 0x7e
    "01111111", -- 3586 - 0xe02  :  127 - 0x7f
    "01111111", -- 3587 - 0xe03  :  127 - 0x7f
    "01111111", -- 3588 - 0xe04  :  127 - 0x7f
    "01111111", -- 3589 - 0xe05  :  127 - 0x7f
    "01111111", -- 3590 - 0xe06  :  127 - 0x7f
    "01111111", -- 3591 - 0xe07  :  127 - 0x7f
    "10000001", -- 3592 - 0xe08  :  129 - 0x81 -- plane 1
    "10000001", -- 3593 - 0xe09  :  129 - 0x81
    "10000001", -- 3594 - 0xe0a  :  129 - 0x81
    "10000001", -- 3595 - 0xe0b  :  129 - 0x81
    "10000001", -- 3596 - 0xe0c  :  129 - 0x81
    "10000001", -- 3597 - 0xe0d  :  129 - 0x81
    "10000001", -- 3598 - 0xe0e  :  129 - 0x81
    "10000001", -- 3599 - 0xe0f  :  129 - 0x81
    "00111111", -- 3600 - 0xe10  :   63 - 0x3f -- Background 0xe1
    "00111111", -- 3601 - 0xe11  :   63 - 0x3f
    "00111111", -- 3602 - 0xe12  :   63 - 0x3f
    "00111111", -- 3603 - 0xe13  :   63 - 0x3f
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "11111111", -- 3608 - 0xe18  :  255 - 0xff -- plane 1
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "11111111", -- 3610 - 0xe1a  :  255 - 0xff
    "11111111", -- 3611 - 0xe1b  :  255 - 0xff
    "11111111", -- 3612 - 0xe1c  :  255 - 0xff
    "11111111", -- 3613 - 0xe1d  :  255 - 0xff
    "11111111", -- 3614 - 0xe1e  :  255 - 0xff
    "11111111", -- 3615 - 0xe1f  :  255 - 0xff
    "01111110", -- 3616 - 0xe20  :  126 - 0x7e -- Background 0xe2
    "01111100", -- 3617 - 0xe21  :  124 - 0x7c
    "01111100", -- 3618 - 0xe22  :  124 - 0x7c
    "01111000", -- 3619 - 0xe23  :  120 - 0x78
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "11111111", -- 3624 - 0xe28  :  255 - 0xff -- plane 1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "11111111", -- 3631 - 0xe2f  :  255 - 0xff
    "11111110", -- 3632 - 0xe30  :  254 - 0xfe -- Background 0xe3
    "11111110", -- 3633 - 0xe31  :  254 - 0xfe
    "11111111", -- 3634 - 0xe32  :  255 - 0xff
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "01111111", -- 3636 - 0xe34  :  127 - 0x7f
    "01111111", -- 3637 - 0xe35  :  127 - 0x7f
    "01111111", -- 3638 - 0xe36  :  127 - 0x7f
    "01111111", -- 3639 - 0xe37  :  127 - 0x7f
    "10000001", -- 3640 - 0xe38  :  129 - 0x81 -- plane 1
    "10000001", -- 3641 - 0xe39  :  129 - 0x81
    "10000001", -- 3642 - 0xe3a  :  129 - 0x81
    "10000001", -- 3643 - 0xe3b  :  129 - 0x81
    "10000001", -- 3644 - 0xe3c  :  129 - 0x81
    "10000001", -- 3645 - 0xe3d  :  129 - 0x81
    "10000001", -- 3646 - 0xe3e  :  129 - 0x81
    "10000001", -- 3647 - 0xe3f  :  129 - 0x81
    "01111111", -- 3648 - 0xe40  :  127 - 0x7f -- Background 0xe4
    "01111111", -- 3649 - 0xe41  :  127 - 0x7f
    "00111111", -- 3650 - 0xe42  :   63 - 0x3f
    "00111111", -- 3651 - 0xe43  :   63 - 0x3f
    "00111111", -- 3652 - 0xe44  :   63 - 0x3f
    "00111111", -- 3653 - 0xe45  :   63 - 0x3f
    "00011111", -- 3654 - 0xe46  :   31 - 0x1f
    "00011111", -- 3655 - 0xe47  :   31 - 0x1f
    "10000000", -- 3656 - 0xe48  :  128 - 0x80 -- plane 1
    "10000000", -- 3657 - 0xe49  :  128 - 0x80
    "11000000", -- 3658 - 0xe4a  :  192 - 0xc0
    "11000000", -- 3659 - 0xe4b  :  192 - 0xc0
    "11100000", -- 3660 - 0xe4c  :  224 - 0xe0
    "11111000", -- 3661 - 0xe4d  :  248 - 0xf8
    "11111110", -- 3662 - 0xe4e  :  254 - 0xfe
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "00111111", -- 3664 - 0xe50  :   63 - 0x3f -- Background 0xe5
    "10111111", -- 3665 - 0xe51  :  191 - 0xbf
    "11111111", -- 3666 - 0xe52  :  255 - 0xff
    "11111111", -- 3667 - 0xe53  :  255 - 0xff
    "11111100", -- 3668 - 0xe54  :  252 - 0xfc
    "11111100", -- 3669 - 0xe55  :  252 - 0xfc
    "11111110", -- 3670 - 0xe56  :  254 - 0xfe
    "11111110", -- 3671 - 0xe57  :  254 - 0xfe
    "11111111", -- 3672 - 0xe58  :  255 - 0xff -- plane 1
    "01111111", -- 3673 - 0xe59  :  127 - 0x7f
    "00011111", -- 3674 - 0xe5a  :   31 - 0x1f
    "00000111", -- 3675 - 0xe5b  :    7 - 0x7
    "00000011", -- 3676 - 0xe5c  :    3 - 0x3
    "00000011", -- 3677 - 0xe5d  :    3 - 0x3
    "00000001", -- 3678 - 0xe5e  :    1 - 0x1
    "10000001", -- 3679 - 0xe5f  :  129 - 0x81
    "01111111", -- 3680 - 0xe60  :  127 - 0x7f -- Background 0xe6
    "01111111", -- 3681 - 0xe61  :  127 - 0x7f
    "01111110", -- 3682 - 0xe62  :  126 - 0x7e
    "01111110", -- 3683 - 0xe63  :  126 - 0x7e
    "01111111", -- 3684 - 0xe64  :  127 - 0x7f
    "01111111", -- 3685 - 0xe65  :  127 - 0x7f
    "01111111", -- 3686 - 0xe66  :  127 - 0x7f
    "01111111", -- 3687 - 0xe67  :  127 - 0x7f
    "10000001", -- 3688 - 0xe68  :  129 - 0x81 -- plane 1
    "10000001", -- 3689 - 0xe69  :  129 - 0x81
    "10000001", -- 3690 - 0xe6a  :  129 - 0x81
    "10000001", -- 3691 - 0xe6b  :  129 - 0x81
    "10000001", -- 3692 - 0xe6c  :  129 - 0x81
    "10000001", -- 3693 - 0xe6d  :  129 - 0x81
    "10000001", -- 3694 - 0xe6e  :  129 - 0x81
    "10000001", -- 3695 - 0xe6f  :  129 - 0x81
    "01111110", -- 3696 - 0xe70  :  126 - 0x7e -- Background 0xe7
    "01111110", -- 3697 - 0xe71  :  126 - 0x7e
    "01111110", -- 3698 - 0xe72  :  126 - 0x7e
    "01111110", -- 3699 - 0xe73  :  126 - 0x7e
    "01111111", -- 3700 - 0xe74  :  127 - 0x7f
    "01111111", -- 3701 - 0xe75  :  127 - 0x7f
    "01111111", -- 3702 - 0xe76  :  127 - 0x7f
    "01111111", -- 3703 - 0xe77  :  127 - 0x7f
    "10000001", -- 3704 - 0xe78  :  129 - 0x81 -- plane 1
    "10000001", -- 3705 - 0xe79  :  129 - 0x81
    "10000001", -- 3706 - 0xe7a  :  129 - 0x81
    "10000001", -- 3707 - 0xe7b  :  129 - 0x81
    "10000001", -- 3708 - 0xe7c  :  129 - 0x81
    "10000001", -- 3709 - 0xe7d  :  129 - 0x81
    "10000001", -- 3710 - 0xe7e  :  129 - 0x81
    "10000001", -- 3711 - 0xe7f  :  129 - 0x81
    "10000001", -- 3712 - 0xe80  :  129 - 0x81 -- Background 0xe8
    "11000011", -- 3713 - 0xe81  :  195 - 0xc3
    "11000011", -- 3714 - 0xe82  :  195 - 0xc3
    "11100111", -- 3715 - 0xe83  :  231 - 0xe7
    "11100111", -- 3716 - 0xe84  :  231 - 0xe7
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "01111110", -- 3720 - 0xe88  :  126 - 0x7e -- plane 1
    "00111100", -- 3721 - 0xe89  :   60 - 0x3c
    "00111100", -- 3722 - 0xe8a  :   60 - 0x3c
    "00011000", -- 3723 - 0xe8b  :   24 - 0x18
    "00011000", -- 3724 - 0xe8c  :   24 - 0x18
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00001111", -- 3728 - 0xe90  :   15 - 0xf -- Background 0xe9
    "01000011", -- 3729 - 0xe91  :   67 - 0x43
    "01011011", -- 3730 - 0xe92  :   91 - 0x5b
    "01010011", -- 3731 - 0xe93  :   83 - 0x53
    "00110001", -- 3732 - 0xe94  :   49 - 0x31
    "00011001", -- 3733 - 0xe95  :   25 - 0x19
    "00001111", -- 3734 - 0xe96  :   15 - 0xf
    "00000111", -- 3735 - 0xe97  :    7 - 0x7
    "11110010", -- 3736 - 0xe98  :  242 - 0xf2 -- plane 1
    "11111110", -- 3737 - 0xe99  :  254 - 0xfe
    "11111110", -- 3738 - 0xe9a  :  254 - 0xfe
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111111", -- 3740 - 0xe9c  :  255 - 0xff
    "11101111", -- 3741 - 0xe9d  :  239 - 0xef
    "11110111", -- 3742 - 0xe9e  :  247 - 0xf7
    "11111000", -- 3743 - 0xe9f  :  248 - 0xf8
    "11000001", -- 3744 - 0xea0  :  193 - 0xc1 -- Background 0xea
    "11000011", -- 3745 - 0xea1  :  195 - 0xc3
    "11000110", -- 3746 - 0xea2  :  198 - 0xc6
    "10000100", -- 3747 - 0xea3  :  132 - 0x84
    "11111100", -- 3748 - 0xea4  :  252 - 0xfc
    "11111100", -- 3749 - 0xea5  :  252 - 0xfc
    "00001110", -- 3750 - 0xea6  :   14 - 0xe
    "00000010", -- 3751 - 0xea7  :    2 - 0x2
    "10111111", -- 3752 - 0xea8  :  191 - 0xbf -- plane 1
    "10111110", -- 3753 - 0xea9  :  190 - 0xbe
    "10111101", -- 3754 - 0xeaa  :  189 - 0xbd
    "01111011", -- 3755 - 0xeab  :  123 - 0x7b
    "01111011", -- 3756 - 0xeac  :  123 - 0x7b
    "00000111", -- 3757 - 0xead  :    7 - 0x7
    "11110011", -- 3758 - 0xeae  :  243 - 0xf3
    "11111101", -- 3759 - 0xeaf  :  253 - 0xfd
    "00010000", -- 3760 - 0xeb0  :   16 - 0x10 -- Background 0xeb
    "00100000", -- 3761 - 0xeb1  :   32 - 0x20
    "00100010", -- 3762 - 0xeb2  :   34 - 0x22
    "10111010", -- 3763 - 0xeb3  :  186 - 0xba
    "11100110", -- 3764 - 0xeb4  :  230 - 0xe6
    "11100001", -- 3765 - 0xeb5  :  225 - 0xe1
    "11000000", -- 3766 - 0xeb6  :  192 - 0xc0
    "11000000", -- 3767 - 0xeb7  :  192 - 0xc0
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff -- plane 1
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "01100111", -- 3771 - 0xebb  :  103 - 0x67
    "01011001", -- 3772 - 0xebc  :   89 - 0x59
    "10011110", -- 3773 - 0xebd  :  158 - 0x9e
    "10111111", -- 3774 - 0xebe  :  191 - 0xbf
    "10111111", -- 3775 - 0xebf  :  191 - 0xbf
    "00100000", -- 3776 - 0xec0  :   32 - 0x20 -- Background 0xec
    "10100110", -- 3777 - 0xec1  :  166 - 0xa6
    "01010100", -- 3778 - 0xec2  :   84 - 0x54
    "00100110", -- 3779 - 0xec3  :   38 - 0x26
    "00100000", -- 3780 - 0xec4  :   32 - 0x20
    "11000110", -- 3781 - 0xec5  :  198 - 0xc6
    "01010100", -- 3782 - 0xec6  :   84 - 0x54
    "00100110", -- 3783 - 0xec7  :   38 - 0x26
    "00100000", -- 3784 - 0xec8  :   32 - 0x20 -- plane 1
    "11100110", -- 3785 - 0xec9  :  230 - 0xe6
    "01010100", -- 3786 - 0xeca  :   84 - 0x54
    "00100110", -- 3787 - 0xecb  :   38 - 0x26
    "00100001", -- 3788 - 0xecc  :   33 - 0x21
    "00000110", -- 3789 - 0xecd  :    6 - 0x6
    "01010100", -- 3790 - 0xece  :   84 - 0x54
    "00100110", -- 3791 - 0xecf  :   38 - 0x26
    "00100000", -- 3792 - 0xed0  :   32 - 0x20 -- Background 0xed
    "10000101", -- 3793 - 0xed1  :  133 - 0x85
    "00000001", -- 3794 - 0xed2  :    1 - 0x1
    "01000100", -- 3795 - 0xed3  :   68 - 0x44
    "00100000", -- 3796 - 0xed4  :   32 - 0x20
    "10000110", -- 3797 - 0xed5  :  134 - 0x86
    "01010100", -- 3798 - 0xed6  :   84 - 0x54
    "01001000", -- 3799 - 0xed7  :   72 - 0x48
    "00100000", -- 3800 - 0xed8  :   32 - 0x20 -- plane 1
    "10011010", -- 3801 - 0xed9  :  154 - 0x9a
    "00000001", -- 3802 - 0xeda  :    1 - 0x1
    "01001001", -- 3803 - 0xedb  :   73 - 0x49
    "00100000", -- 3804 - 0xedc  :   32 - 0x20
    "10100101", -- 3805 - 0xedd  :  165 - 0xa5
    "11001001", -- 3806 - 0xede  :  201 - 0xc9
    "01000110", -- 3807 - 0xedf  :   70 - 0x46
    "00100000", -- 3808 - 0xee0  :   32 - 0x20 -- Background 0xee
    "10111010", -- 3809 - 0xee1  :  186 - 0xba
    "11001001", -- 3810 - 0xee2  :  201 - 0xc9
    "01001010", -- 3811 - 0xee3  :   74 - 0x4a
    "00100000", -- 3812 - 0xee4  :   32 - 0x20
    "10100110", -- 3813 - 0xee5  :  166 - 0xa6
    "00001010", -- 3814 - 0xee6  :   10 - 0xa
    "11010000", -- 3815 - 0xee7  :  208 - 0xd0
    "11010001", -- 3816 - 0xee8  :  209 - 0xd1 -- plane 1
    "11011000", -- 3817 - 0xee9  :  216 - 0xd8
    "11011000", -- 3818 - 0xeea  :  216 - 0xd8
    "11011110", -- 3819 - 0xeeb  :  222 - 0xde
    "11010001", -- 3820 - 0xeec  :  209 - 0xd1
    "11010000", -- 3821 - 0xeed  :  208 - 0xd0
    "11011010", -- 3822 - 0xeee  :  218 - 0xda
    "11011110", -- 3823 - 0xeef  :  222 - 0xde
    "11010001", -- 3824 - 0xef0  :  209 - 0xd1 -- Background 0xef
    "00100000", -- 3825 - 0xef1  :   32 - 0x20
    "11000110", -- 3826 - 0xef2  :  198 - 0xc6
    "00001010", -- 3827 - 0xef3  :   10 - 0xa
    "11010010", -- 3828 - 0xef4  :  210 - 0xd2
    "11010011", -- 3829 - 0xef5  :  211 - 0xd3
    "11011011", -- 3830 - 0xef6  :  219 - 0xdb
    "11011011", -- 3831 - 0xef7  :  219 - 0xdb
    "11011011", -- 3832 - 0xef8  :  219 - 0xdb -- plane 1
    "11011001", -- 3833 - 0xef9  :  217 - 0xd9
    "11011011", -- 3834 - 0xefa  :  219 - 0xdb
    "11011100", -- 3835 - 0xefb  :  220 - 0xdc
    "11011011", -- 3836 - 0xefc  :  219 - 0xdb
    "11011111", -- 3837 - 0xefd  :  223 - 0xdf
    "00100000", -- 3838 - 0xefe  :   32 - 0x20
    "11100110", -- 3839 - 0xeff  :  230 - 0xe6
    "00001010", -- 3840 - 0xf00  :   10 - 0xa -- Background 0xf0
    "11010100", -- 3841 - 0xf01  :  212 - 0xd4
    "11010101", -- 3842 - 0xf02  :  213 - 0xd5
    "11010100", -- 3843 - 0xf03  :  212 - 0xd4
    "11011001", -- 3844 - 0xf04  :  217 - 0xd9
    "11011011", -- 3845 - 0xf05  :  219 - 0xdb
    "11100010", -- 3846 - 0xf06  :  226 - 0xe2
    "11010100", -- 3847 - 0xf07  :  212 - 0xd4
    "11011010", -- 3848 - 0xf08  :  218 - 0xda -- plane 1
    "11011011", -- 3849 - 0xf09  :  219 - 0xdb
    "11100000", -- 3850 - 0xf0a  :  224 - 0xe0
    "00100001", -- 3851 - 0xf0b  :   33 - 0x21
    "00000110", -- 3852 - 0xf0c  :    6 - 0x6
    "00001010", -- 3853 - 0xf0d  :   10 - 0xa
    "11010110", -- 3854 - 0xf0e  :  214 - 0xd6
    "11010111", -- 3855 - 0xf0f  :  215 - 0xd7
    "11010110", -- 3856 - 0xf10  :  214 - 0xd6 -- Background 0xf1
    "11010111", -- 3857 - 0xf11  :  215 - 0xd7
    "11100001", -- 3858 - 0xf12  :  225 - 0xe1
    "00100110", -- 3859 - 0xf13  :   38 - 0x26
    "11010110", -- 3860 - 0xf14  :  214 - 0xd6
    "11011101", -- 3861 - 0xf15  :  221 - 0xdd
    "11100001", -- 3862 - 0xf16  :  225 - 0xe1
    "11100001", -- 3863 - 0xf17  :  225 - 0xe1
    "00100001", -- 3864 - 0xf18  :   33 - 0x21 -- plane 1
    "00100110", -- 3865 - 0xf19  :   38 - 0x26
    "00010100", -- 3866 - 0xf1a  :   20 - 0x14
    "11010000", -- 3867 - 0xf1b  :  208 - 0xd0
    "11101000", -- 3868 - 0xf1c  :  232 - 0xe8
    "11010001", -- 3869 - 0xf1d  :  209 - 0xd1
    "11010000", -- 3870 - 0xf1e  :  208 - 0xd0
    "11010001", -- 3871 - 0xf1f  :  209 - 0xd1
    "11011110", -- 3872 - 0xf20  :  222 - 0xde -- Background 0xf2
    "11010001", -- 3873 - 0xf21  :  209 - 0xd1
    "11011000", -- 3874 - 0xf22  :  216 - 0xd8
    "11010000", -- 3875 - 0xf23  :  208 - 0xd0
    "11010001", -- 3876 - 0xf24  :  209 - 0xd1
    "00100110", -- 3877 - 0xf25  :   38 - 0x26
    "11011110", -- 3878 - 0xf26  :  222 - 0xde
    "11010001", -- 3879 - 0xf27  :  209 - 0xd1
    "11011110", -- 3880 - 0xf28  :  222 - 0xde -- plane 1
    "11010001", -- 3881 - 0xf29  :  209 - 0xd1
    "11010000", -- 3882 - 0xf2a  :  208 - 0xd0
    "11010001", -- 3883 - 0xf2b  :  209 - 0xd1
    "11010000", -- 3884 - 0xf2c  :  208 - 0xd0
    "11010001", -- 3885 - 0xf2d  :  209 - 0xd1
    "00100110", -- 3886 - 0xf2e  :   38 - 0x26
    "00100001", -- 3887 - 0xf2f  :   33 - 0x21
    "01000110", -- 3888 - 0xf30  :   70 - 0x46 -- Background 0xf3
    "00010100", -- 3889 - 0xf31  :   20 - 0x14
    "11011011", -- 3890 - 0xf32  :  219 - 0xdb
    "01000010", -- 3891 - 0xf33  :   66 - 0x42
    "01000010", -- 3892 - 0xf34  :   66 - 0x42
    "11011011", -- 3893 - 0xf35  :  219 - 0xdb
    "01000010", -- 3894 - 0xf36  :   66 - 0x42
    "11011011", -- 3895 - 0xf37  :  219 - 0xdb
    "01000010", -- 3896 - 0xf38  :   66 - 0x42 -- plane 1
    "11011011", -- 3897 - 0xf39  :  219 - 0xdb
    "11011011", -- 3898 - 0xf3a  :  219 - 0xdb
    "01000010", -- 3899 - 0xf3b  :   66 - 0x42
    "00100110", -- 3900 - 0xf3c  :   38 - 0x26
    "11011011", -- 3901 - 0xf3d  :  219 - 0xdb
    "01000010", -- 3902 - 0xf3e  :   66 - 0x42
    "11011011", -- 3903 - 0xf3f  :  219 - 0xdb
    "01000010", -- 3904 - 0xf40  :   66 - 0x42 -- Background 0xf4
    "11011011", -- 3905 - 0xf41  :  219 - 0xdb
    "01000010", -- 3906 - 0xf42  :   66 - 0x42
    "11011011", -- 3907 - 0xf43  :  219 - 0xdb
    "01000010", -- 3908 - 0xf44  :   66 - 0x42
    "00100110", -- 3909 - 0xf45  :   38 - 0x26
    "00100001", -- 3910 - 0xf46  :   33 - 0x21
    "01100110", -- 3911 - 0xf47  :  102 - 0x66
    "01000110", -- 3912 - 0xf48  :   70 - 0x46 -- plane 1
    "11011011", -- 3913 - 0xf49  :  219 - 0xdb
    "00100001", -- 3914 - 0xf4a  :   33 - 0x21
    "01101100", -- 3915 - 0xf4b  :  108 - 0x6c
    "00001110", -- 3916 - 0xf4c  :   14 - 0xe
    "11011111", -- 3917 - 0xf4d  :  223 - 0xdf
    "11011011", -- 3918 - 0xf4e  :  219 - 0xdb
    "11011011", -- 3919 - 0xf4f  :  219 - 0xdb
    "11011011", -- 3920 - 0xf50  :  219 - 0xdb -- Background 0xf5
    "00100110", -- 3921 - 0xf51  :   38 - 0x26
    "11011011", -- 3922 - 0xf52  :  219 - 0xdb
    "11011111", -- 3923 - 0xf53  :  223 - 0xdf
    "11011011", -- 3924 - 0xf54  :  219 - 0xdb
    "11011111", -- 3925 - 0xf55  :  223 - 0xdf
    "11011011", -- 3926 - 0xf56  :  219 - 0xdb
    "11011011", -- 3927 - 0xf57  :  219 - 0xdb
    "11100100", -- 3928 - 0xf58  :  228 - 0xe4 -- plane 1
    "11100101", -- 3929 - 0xf59  :  229 - 0xe5
    "00100110", -- 3930 - 0xf5a  :   38 - 0x26
    "00100001", -- 3931 - 0xf5b  :   33 - 0x21
    "10000110", -- 3932 - 0xf5c  :  134 - 0x86
    "00010100", -- 3933 - 0xf5d  :   20 - 0x14
    "11011011", -- 3934 - 0xf5e  :  219 - 0xdb
    "11011011", -- 3935 - 0xf5f  :  219 - 0xdb
    "11011011", -- 3936 - 0xf60  :  219 - 0xdb -- Background 0xf6
    "11011110", -- 3937 - 0xf61  :  222 - 0xde
    "01000011", -- 3938 - 0xf62  :   67 - 0x43
    "11011011", -- 3939 - 0xf63  :  219 - 0xdb
    "11100000", -- 3940 - 0xf64  :  224 - 0xe0
    "11011011", -- 3941 - 0xf65  :  219 - 0xdb
    "11011011", -- 3942 - 0xf66  :  219 - 0xdb
    "11011011", -- 3943 - 0xf67  :  219 - 0xdb
    "00100110", -- 3944 - 0xf68  :   38 - 0x26 -- plane 1
    "11011011", -- 3945 - 0xf69  :  219 - 0xdb
    "11100011", -- 3946 - 0xf6a  :  227 - 0xe3
    "11011011", -- 3947 - 0xf6b  :  219 - 0xdb
    "11100000", -- 3948 - 0xf6c  :  224 - 0xe0
    "11011011", -- 3949 - 0xf6d  :  219 - 0xdb
    "11011011", -- 3950 - 0xf6e  :  219 - 0xdb
    "11100110", -- 3951 - 0xf6f  :  230 - 0xe6
    "11100011", -- 3952 - 0xf70  :  227 - 0xe3 -- Background 0xf7
    "00100110", -- 3953 - 0xf71  :   38 - 0x26
    "00100001", -- 3954 - 0xf72  :   33 - 0x21
    "10100110", -- 3955 - 0xf73  :  166 - 0xa6
    "00010100", -- 3956 - 0xf74  :   20 - 0x14
    "11011011", -- 3957 - 0xf75  :  219 - 0xdb
    "11011011", -- 3958 - 0xf76  :  219 - 0xdb
    "11011011", -- 3959 - 0xf77  :  219 - 0xdb
    "11011011", -- 3960 - 0xf78  :  219 - 0xdb -- plane 1
    "01000010", -- 3961 - 0xf79  :   66 - 0x42
    "11011011", -- 3962 - 0xf7a  :  219 - 0xdb
    "11011011", -- 3963 - 0xf7b  :  219 - 0xdb
    "11011011", -- 3964 - 0xf7c  :  219 - 0xdb
    "11010100", -- 3965 - 0xf7d  :  212 - 0xd4
    "11011001", -- 3966 - 0xf7e  :  217 - 0xd9
    "00100110", -- 3967 - 0xf7f  :   38 - 0x26
    "11011011", -- 3968 - 0xf80  :  219 - 0xdb -- Background 0xf8
    "11011001", -- 3969 - 0xf81  :  217 - 0xd9
    "11011011", -- 3970 - 0xf82  :  219 - 0xdb
    "11011011", -- 3971 - 0xf83  :  219 - 0xdb
    "11010100", -- 3972 - 0xf84  :  212 - 0xd4
    "11011001", -- 3973 - 0xf85  :  217 - 0xd9
    "11010100", -- 3974 - 0xf86  :  212 - 0xd4
    "11011001", -- 3975 - 0xf87  :  217 - 0xd9
    "11100111", -- 3976 - 0xf88  :  231 - 0xe7 -- plane 1
    "00100001", -- 3977 - 0xf89  :   33 - 0x21
    "11000101", -- 3978 - 0xf8a  :  197 - 0xc5
    "00010110", -- 3979 - 0xf8b  :   22 - 0x16
    "01011111", -- 3980 - 0xf8c  :   95 - 0x5f
    "10010101", -- 3981 - 0xf8d  :  149 - 0x95
    "10010101", -- 3982 - 0xf8e  :  149 - 0x95
    "10010101", -- 3983 - 0xf8f  :  149 - 0x95
    "10010101", -- 3984 - 0xf90  :  149 - 0x95 -- Background 0xf9
    "10010101", -- 3985 - 0xf91  :  149 - 0x95
    "10010101", -- 3986 - 0xf92  :  149 - 0x95
    "10010101", -- 3987 - 0xf93  :  149 - 0x95
    "10010101", -- 3988 - 0xf94  :  149 - 0x95
    "10010111", -- 3989 - 0xf95  :  151 - 0x97
    "10011000", -- 3990 - 0xf96  :  152 - 0x98
    "01111000", -- 3991 - 0xf97  :  120 - 0x78
    "10010101", -- 3992 - 0xf98  :  149 - 0x95 -- plane 1
    "10010110", -- 3993 - 0xf99  :  150 - 0x96
    "10010101", -- 3994 - 0xf9a  :  149 - 0x95
    "10010101", -- 3995 - 0xf9b  :  149 - 0x95
    "10010111", -- 3996 - 0xf9c  :  151 - 0x97
    "10011000", -- 3997 - 0xf9d  :  152 - 0x98
    "10010111", -- 3998 - 0xf9e  :  151 - 0x97
    "10011000", -- 3999 - 0xf9f  :  152 - 0x98
    "10010101", -- 4000 - 0xfa0  :  149 - 0x95 -- Background 0xfa
    "01111010", -- 4001 - 0xfa1  :  122 - 0x7a
    "00100001", -- 4002 - 0xfa2  :   33 - 0x21
    "11101101", -- 4003 - 0xfa3  :  237 - 0xed
    "00001110", -- 4004 - 0xfa4  :   14 - 0xe
    "11001111", -- 4005 - 0xfa5  :  207 - 0xcf
    "00000001", -- 4006 - 0xfa6  :    1 - 0x1
    "00001001", -- 4007 - 0xfa7  :    9 - 0x9
    "00001000", -- 4008 - 0xfa8  :    8 - 0x8 -- plane 1
    "00000101", -- 4009 - 0xfa9  :    5 - 0x5
    "00100100", -- 4010 - 0xfaa  :   36 - 0x24
    "00010111", -- 4011 - 0xfab  :   23 - 0x17
    "00010010", -- 4012 - 0xfac  :   18 - 0x12
    "00010111", -- 4013 - 0xfad  :   23 - 0x17
    "00011101", -- 4014 - 0xfae  :   29 - 0x1d
    "00001110", -- 4015 - 0xfaf  :   14 - 0xe
    "00010111", -- 4016 - 0xfb0  :   23 - 0x17 -- Background 0xfb
    "00001101", -- 4017 - 0xfb1  :   13 - 0xd
    "00011000", -- 4018 - 0xfb2  :   24 - 0x18
    "00100010", -- 4019 - 0xfb3  :   34 - 0x22
    "01001011", -- 4020 - 0xfb4  :   75 - 0x4b
    "00001101", -- 4021 - 0xfb5  :   13 - 0xd
    "00000001", -- 4022 - 0xfb6  :    1 - 0x1
    "00100100", -- 4023 - 0xfb7  :   36 - 0x24
    "00011001", -- 4024 - 0xfb8  :   25 - 0x19 -- plane 1
    "00010101", -- 4025 - 0xfb9  :   21 - 0x15
    "00001010", -- 4026 - 0xfba  :   10 - 0xa
    "00100010", -- 4027 - 0xfbb  :   34 - 0x22
    "00001110", -- 4028 - 0xfbc  :   14 - 0xe
    "00011011", -- 4029 - 0xfbd  :   27 - 0x1b
    "00100100", -- 4030 - 0xfbe  :   36 - 0x24
    "00010000", -- 4031 - 0xfbf  :   16 - 0x10
    "00001010", -- 4032 - 0xfc0  :   10 - 0xa -- Background 0xfc
    "00010110", -- 4033 - 0xfc1  :   22 - 0x16
    "00001110", -- 4034 - 0xfc2  :   14 - 0xe
    "00100010", -- 4035 - 0xfc3  :   34 - 0x22
    "10001011", -- 4036 - 0xfc4  :  139 - 0x8b
    "00001101", -- 4037 - 0xfc5  :   13 - 0xd
    "00000010", -- 4038 - 0xfc6  :    2 - 0x2
    "00100100", -- 4039 - 0xfc7  :   36 - 0x24
    "00011001", -- 4040 - 0xfc8  :   25 - 0x19 -- plane 1
    "00010101", -- 4041 - 0xfc9  :   21 - 0x15
    "00001010", -- 4042 - 0xfca  :   10 - 0xa
    "00100010", -- 4043 - 0xfcb  :   34 - 0x22
    "00001110", -- 4044 - 0xfcc  :   14 - 0xe
    "00011011", -- 4045 - 0xfcd  :   27 - 0x1b
    "00100100", -- 4046 - 0xfce  :   36 - 0x24
    "00010000", -- 4047 - 0xfcf  :   16 - 0x10
    "00001010", -- 4048 - 0xfd0  :   10 - 0xa -- Background 0xfd
    "00010110", -- 4049 - 0xfd1  :   22 - 0x16
    "00001110", -- 4050 - 0xfd2  :   14 - 0xe
    "00100010", -- 4051 - 0xfd3  :   34 - 0x22
    "11101100", -- 4052 - 0xfd4  :  236 - 0xec
    "00000100", -- 4053 - 0xfd5  :    4 - 0x4
    "00011101", -- 4054 - 0xfd6  :   29 - 0x1d
    "00011000", -- 4055 - 0xfd7  :   24 - 0x18
    "00011001", -- 4056 - 0xfd8  :   25 - 0x19 -- plane 1
    "00101000", -- 4057 - 0xfd9  :   40 - 0x28
    "00100010", -- 4058 - 0xfda  :   34 - 0x22
    "11110110", -- 4059 - 0xfdb  :  246 - 0xf6
    "00000001", -- 4060 - 0xfdc  :    1 - 0x1
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00100011", -- 4062 - 0xfde  :   35 - 0x23
    "11001001", -- 4063 - 0xfdf  :  201 - 0xc9
    "01010110", -- 4064 - 0xfe0  :   86 - 0x56 -- Background 0xfe
    "01010101", -- 4065 - 0xfe1  :   85 - 0x55
    "00100011", -- 4066 - 0xfe2  :   35 - 0x23
    "11100010", -- 4067 - 0xfe3  :  226 - 0xe2
    "00000100", -- 4068 - 0xfe4  :    4 - 0x4
    "10011001", -- 4069 - 0xfe5  :  153 - 0x99
    "10101010", -- 4070 - 0xfe6  :  170 - 0xaa
    "10101010", -- 4071 - 0xfe7  :  170 - 0xaa
    "10101010", -- 4072 - 0xfe8  :  170 - 0xaa -- plane 1
    "00100011", -- 4073 - 0xfe9  :   35 - 0x23
    "11101010", -- 4074 - 0xfea  :  234 - 0xea
    "00000100", -- 4075 - 0xfeb  :    4 - 0x4
    "10011001", -- 4076 - 0xfec  :  153 - 0x99
    "10101010", -- 4077 - 0xfed  :  170 - 0xaa
    "10101010", -- 4078 - 0xfee  :  170 - 0xaa
    "10101010", -- 4079 - 0xfef  :  170 - 0xaa
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff -- plane 1
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
