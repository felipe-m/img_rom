--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Pattern Table 0---------
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000011", --    1 -  0x1  :    3 - 0x3
    "00001111", --    2 -  0x2  :   15 - 0xf
    "00011111", --    3 -  0x3  :   31 - 0x1f
    "00111111", --    4 -  0x4  :   63 - 0x3f
    "00111111", --    5 -  0x5  :   63 - 0x3f
    "01111111", --    6 -  0x6  :  127 - 0x7f
    "01111111", --    7 -  0x7  :  127 - 0x7f
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x1
    "11000000", --   17 - 0x11  :  192 - 0xc0
    "11110000", --   18 - 0x12  :  240 - 0xf0
    "11111000", --   19 - 0x13  :  248 - 0xf8
    "11111000", --   20 - 0x14  :  248 - 0xf8
    "11111100", --   21 - 0x15  :  252 - 0xfc
    "11111100", --   22 - 0x16  :  252 - 0xfc
    "11111100", --   23 - 0x17  :  252 - 0xfc
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "00000111", --   33 - 0x21  :    7 - 0x7
    "00011111", --   34 - 0x22  :   31 - 0x1f
    "00111111", --   35 - 0x23  :   63 - 0x3f
    "00111111", --   36 - 0x24  :   63 - 0x3f
    "00001111", --   37 - 0x25  :   15 - 0xf
    "00000011", --   38 - 0x26  :    3 - 0x3
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000111", --   50 - 0x32  :    7 - 0x7
    "00011111", --   51 - 0x33  :   31 - 0x1f
    "00111111", --   52 - 0x34  :   63 - 0x3f
    "00111111", --   53 - 0x35  :   63 - 0x3f
    "01111111", --   54 - 0x36  :  127 - 0x7f
    "01111111", --   55 - 0x37  :  127 - 0x7f
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "01111110", --   64 - 0x40  :  126 - 0x7e -- Sprite 0x4
    "01111110", --   65 - 0x41  :  126 - 0x7e
    "01111100", --   66 - 0x42  :  124 - 0x7c
    "00111100", --   67 - 0x43  :   60 - 0x3c
    "00111000", --   68 - 0x44  :   56 - 0x38
    "00011000", --   69 - 0x45  :   24 - 0x18
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0x5
    "11000000", --   81 - 0x51  :  192 - 0xc0
    "11110000", --   82 - 0x52  :  240 - 0xf0
    "11111000", --   83 - 0x53  :  248 - 0xf8
    "11111000", --   84 - 0x54  :  248 - 0xf8
    "11111100", --   85 - 0x55  :  252 - 0xfc
    "01111100", --   86 - 0x56  :  124 - 0x7c
    "00111100", --   87 - 0x57  :   60 - 0x3c
    "00000000", --   88 - 0x58  :    0 - 0x0
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0x6
    "00000111", --   97 - 0x61  :    7 - 0x7
    "00000111", --   98 - 0x62  :    7 - 0x7
    "00000011", --   99 - 0x63  :    3 - 0x3
    "00000001", --  100 - 0x64  :    1 - 0x1
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0x7
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000111", --  114 - 0x72  :    7 - 0x7
    "00011111", --  115 - 0x73  :   31 - 0x1f
    "00111111", --  116 - 0x74  :   63 - 0x3f
    "00111111", --  117 - 0x75  :   63 - 0x3f
    "01111110", --  118 - 0x76  :  126 - 0x7e
    "01111100", --  119 - 0x77  :  124 - 0x7c
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "01111000", --  128 - 0x80  :  120 - 0x78 -- Sprite 0x8
    "01110000", --  129 - 0x81  :  112 - 0x70
    "01100000", --  130 - 0x82  :   96 - 0x60
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x9
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "01000000", --  149 - 0x95  :   64 - 0x40
    "11110000", --  150 - 0x96  :  240 - 0xf0
    "11111000", --  151 - 0x97  :  248 - 0xf8
    "00000000", --  152 - 0x98  :    0 - 0x0
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "11111110", --  160 - 0xa0  :  254 - 0xfe -- Sprite 0xa
    "01111111", --  161 - 0xa1  :  127 - 0x7f
    "01111111", --  162 - 0xa2  :  127 - 0x7f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00001110", --  164 - 0xa4  :   14 - 0xe
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0xb
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "11100000", --  183 - 0xb7  :  224 - 0xe0
    "00000000", --  184 - 0xb8  :    0 - 0x0
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "11111100", --  192 - 0xc0  :  252 - 0xfc -- Sprite 0xc
    "11111111", --  193 - 0xc1  :  255 - 0xff
    "01111111", --  194 - 0xc2  :  127 - 0x7f
    "00111111", --  195 - 0xc3  :   63 - 0x3f
    "00001110", --  196 - 0xc4  :   14 - 0xe
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "11110000", --  208 - 0xd0  :  240 - 0xf0 -- Sprite 0xd
    "11111111", --  209 - 0xd1  :  255 - 0xff
    "11111111", --  210 - 0xd2  :  255 - 0xff
    "01111111", --  211 - 0xd3  :  127 - 0x7f
    "00011110", --  212 - 0xd4  :   30 - 0x1e
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00001111", --  225 - 0xe1  :   15 - 0xf
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111111", --  227 - 0xe3  :  255 - 0xff
    "01111111", --  228 - 0xe4  :  127 - 0x7f
    "00011110", --  229 - 0xe5  :   30 - 0x1e
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0xf
    "00000011", --  241 - 0xf1  :    3 - 0x3
    "00001111", --  242 - 0xf2  :   15 - 0xf
    "01111111", --  243 - 0xf3  :  127 - 0x7f
    "11111111", --  244 - 0xf4  :  255 - 0xff
    "01111110", --  245 - 0xf5  :  126 - 0x7e
    "00011100", --  246 - 0xf6  :   28 - 0x1c
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000001", --  257 - 0x101  :    1 - 0x1
    "00000011", --  258 - 0x102  :    3 - 0x3
    "00001111", --  259 - 0x103  :   15 - 0xf
    "00011111", --  260 - 0x104  :   31 - 0x1f
    "01111111", --  261 - 0x105  :  127 - 0x7f
    "01111110", --  262 - 0x106  :  126 - 0x7e
    "00111100", --  263 - 0x107  :   60 - 0x3c
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x11
    "00000001", --  273 - 0x111  :    1 - 0x1
    "00000011", --  274 - 0x112  :    3 - 0x3
    "00000111", --  275 - 0x113  :    7 - 0x7
    "00000111", --  276 - 0x114  :    7 - 0x7
    "00001111", --  277 - 0x115  :   15 - 0xf
    "00011111", --  278 - 0x116  :   31 - 0x1f
    "00001110", --  279 - 0x117  :   14 - 0xe
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x12
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000001", --  290 - 0x122  :    1 - 0x1
    "00000011", --  291 - 0x123  :    3 - 0x3
    "00000011", --  292 - 0x124  :    3 - 0x3
    "00000011", --  293 - 0x125  :    3 - 0x3
    "00000111", --  294 - 0x126  :    7 - 0x7
    "00000010", --  295 - 0x127  :    2 - 0x2
    "00000000", --  296 - 0x128  :    0 - 0x0
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000001", --  306 - 0x132  :    1 - 0x1
    "00000001", --  307 - 0x133  :    1 - 0x1
    "00000001", --  308 - 0x134  :    1 - 0x1
    "00000001", --  309 - 0x135  :    1 - 0x1
    "00000001", --  310 - 0x136  :    1 - 0x1
    "00000001", --  311 - 0x137  :    1 - 0x1
    "00000000", --  312 - 0x138  :    0 - 0x0
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x14
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000100", --  326 - 0x146  :    4 - 0x4
    "00000010", --  327 - 0x147  :    2 - 0x2
    "00000000", --  328 - 0x148  :    0 - 0x0
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Sprite 0x15
    "00000000", --  337 - 0x151  :    0 - 0x0
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00100000", --  342 - 0x156  :   32 - 0x20
    "01001000", --  343 - 0x157  :   72 - 0x48
    "00000000", --  344 - 0x158  :    0 - 0x0
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00010000", --  352 - 0x160  :   16 - 0x10 -- Sprite 0x16
    "00001000", --  353 - 0x161  :    8 - 0x8
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00110000", --  355 - 0x163  :   48 - 0x30
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00001000", --  357 - 0x165  :    8 - 0x8
    "00010010", --  358 - 0x166  :   18 - 0x12
    "00000100", --  359 - 0x167  :    4 - 0x4
    "00000000", --  360 - 0x168  :    0 - 0x0
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00010000", --  368 - 0x170  :   16 - 0x10 -- Sprite 0x17
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00001100", --  370 - 0x172  :   12 - 0xc
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00010000", --  372 - 0x174  :   16 - 0x10
    "00001000", --  373 - 0x175  :    8 - 0x8
    "01000000", --  374 - 0x176  :   64 - 0x40
    "00100000", --  375 - 0x177  :   32 - 0x20
    "00000000", --  376 - 0x178  :    0 - 0x0
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000011", --  386 - 0x182  :    3 - 0x3
    "00000011", --  387 - 0x183  :    3 - 0x3
    "00000001", --  388 - 0x184  :    1 - 0x1
    "00100001", --  389 - 0x185  :   33 - 0x21
    "00100001", --  390 - 0x186  :   33 - 0x21
    "01110011", --  391 - 0x187  :  115 - 0x73
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000011", --  394 - 0x18a  :    3 - 0x3
    "00000011", --  395 - 0x18b  :    3 - 0x3
    "00010011", --  396 - 0x18c  :   19 - 0x13
    "00111111", --  397 - 0x18d  :   63 - 0x3f
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "01111111", --  399 - 0x18f  :  127 - 0x7f
    "01111111", --  400 - 0x190  :  127 - 0x7f -- Sprite 0x19
    "01111111", --  401 - 0x191  :  127 - 0x7f
    "01111111", --  402 - 0x192  :  127 - 0x7f
    "01111111", --  403 - 0x193  :  127 - 0x7f
    "01101110", --  404 - 0x194  :  110 - 0x6e
    "01000110", --  405 - 0x195  :   70 - 0x46
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "01111111", --  408 - 0x198  :  127 - 0x7f
    "01111111", --  409 - 0x199  :  127 - 0x7f
    "01111111", --  410 - 0x19a  :  127 - 0x7f
    "01111111", --  411 - 0x19b  :  127 - 0x7f
    "01101110", --  412 - 0x19c  :  110 - 0x6e
    "01000110", --  413 - 0x19d  :   70 - 0x46
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "01111111", --  416 - 0x1a0  :  127 - 0x7f -- Sprite 0x1a
    "01111111", --  417 - 0x1a1  :  127 - 0x7f
    "01111111", --  418 - 0x1a2  :  127 - 0x7f
    "01111111", --  419 - 0x1a3  :  127 - 0x7f
    "01111011", --  420 - 0x1a4  :  123 - 0x7b
    "00110001", --  421 - 0x1a5  :   49 - 0x31
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "01111111", --  424 - 0x1a8  :  127 - 0x7f
    "01111111", --  425 - 0x1a9  :  127 - 0x7f
    "01111111", --  426 - 0x1aa  :  127 - 0x7f
    "01111111", --  427 - 0x1ab  :  127 - 0x7f
    "01111011", --  428 - 0x1ac  :  123 - 0x7b
    "00110001", --  429 - 0x1ad  :   49 - 0x31
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "00000011", --  433 - 0x1b1  :    3 - 0x3
    "00001111", --  434 - 0x1b2  :   15 - 0xf
    "00011111", --  435 - 0x1b3  :   31 - 0x1f
    "00100111", --  436 - 0x1b4  :   39 - 0x27
    "00000011", --  437 - 0x1b5  :    3 - 0x3
    "00000011", --  438 - 0x1b6  :    3 - 0x3
    "01000011", --  439 - 0x1b7  :   67 - 0x43
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "00000011", --  441 - 0x1b9  :    3 - 0x3
    "00001111", --  442 - 0x1ba  :   15 - 0xf
    "00011111", --  443 - 0x1bb  :   31 - 0x1f
    "00111111", --  444 - 0x1bc  :   63 - 0x3f
    "00111111", --  445 - 0x1bd  :   63 - 0x3f
    "00001111", --  446 - 0x1be  :   15 - 0xf
    "01001111", --  447 - 0x1bf  :   79 - 0x4f
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x1c
    "11000000", --  449 - 0x1c1  :  192 - 0xc0
    "11110000", --  450 - 0x1c2  :  240 - 0xf0
    "11111000", --  451 - 0x1c3  :  248 - 0xf8
    "10011100", --  452 - 0x1c4  :  156 - 0x9c
    "00001100", --  453 - 0x1c5  :   12 - 0xc
    "00001100", --  454 - 0x1c6  :   12 - 0xc
    "00001110", --  455 - 0x1c7  :   14 - 0xe
    "00000000", --  456 - 0x1c8  :    0 - 0x0
    "11000000", --  457 - 0x1c9  :  192 - 0xc0
    "11110000", --  458 - 0x1ca  :  240 - 0xf0
    "11111000", --  459 - 0x1cb  :  248 - 0xf8
    "11111100", --  460 - 0x1cc  :  252 - 0xfc
    "11111100", --  461 - 0x1cd  :  252 - 0xfc
    "00111100", --  462 - 0x1ce  :   60 - 0x3c
    "00111110", --  463 - 0x1cf  :   62 - 0x3e
    "01100111", --  464 - 0x1d0  :  103 - 0x67 -- Sprite 0x1d
    "01111111", --  465 - 0x1d1  :  127 - 0x7f
    "01111111", --  466 - 0x1d2  :  127 - 0x7f
    "01111111", --  467 - 0x1d3  :  127 - 0x7f
    "01101110", --  468 - 0x1d4  :  110 - 0x6e
    "01000110", --  469 - 0x1d5  :   70 - 0x46
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "01111111", --  472 - 0x1d8  :  127 - 0x7f
    "01111111", --  473 - 0x1d9  :  127 - 0x7f
    "01111111", --  474 - 0x1da  :  127 - 0x7f
    "01111111", --  475 - 0x1db  :  127 - 0x7f
    "01101110", --  476 - 0x1dc  :  110 - 0x6e
    "01000110", --  477 - 0x1dd  :   70 - 0x46
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "01100111", --  480 - 0x1e0  :  103 - 0x67 -- Sprite 0x1e
    "01111111", --  481 - 0x1e1  :  127 - 0x7f
    "01111111", --  482 - 0x1e2  :  127 - 0x7f
    "01111111", --  483 - 0x1e3  :  127 - 0x7f
    "01111011", --  484 - 0x1e4  :  123 - 0x7b
    "00110001", --  485 - 0x1e5  :   49 - 0x31
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "01111111", --  488 - 0x1e8  :  127 - 0x7f
    "01111111", --  489 - 0x1e9  :  127 - 0x7f
    "01111111", --  490 - 0x1ea  :  127 - 0x7f
    "01111111", --  491 - 0x1eb  :  127 - 0x7f
    "01111011", --  492 - 0x1ec  :  123 - 0x7b
    "00110001", --  493 - 0x1ed  :   49 - 0x31
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "10011110", --  496 - 0x1f0  :  158 - 0x9e -- Sprite 0x1f
    "11111110", --  497 - 0x1f1  :  254 - 0xfe
    "11111110", --  498 - 0x1f2  :  254 - 0xfe
    "11111110", --  499 - 0x1f3  :  254 - 0xfe
    "01110110", --  500 - 0x1f4  :  118 - 0x76
    "01100010", --  501 - 0x1f5  :   98 - 0x62
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11111110", --  504 - 0x1f8  :  254 - 0xfe
    "11111110", --  505 - 0x1f9  :  254 - 0xfe
    "11111110", --  506 - 0x1fa  :  254 - 0xfe
    "11111110", --  507 - 0x1fb  :  254 - 0xfe
    "01110110", --  508 - 0x1fc  :  118 - 0x76
    "01100010", --  509 - 0x1fd  :   98 - 0x62
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "10011110", --  512 - 0x200  :  158 - 0x9e -- Sprite 0x20
    "11111110", --  513 - 0x201  :  254 - 0xfe
    "11111110", --  514 - 0x202  :  254 - 0xfe
    "11111110", --  515 - 0x203  :  254 - 0xfe
    "11011110", --  516 - 0x204  :  222 - 0xde
    "10001100", --  517 - 0x205  :  140 - 0x8c
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "11111110", --  520 - 0x208  :  254 - 0xfe
    "11111110", --  521 - 0x209  :  254 - 0xfe
    "11111110", --  522 - 0x20a  :  254 - 0xfe
    "11111110", --  523 - 0x20b  :  254 - 0xfe
    "11011110", --  524 - 0x20c  :  222 - 0xde
    "10001100", --  525 - 0x20d  :  140 - 0x8c
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x21
    "00000011", --  529 - 0x211  :    3 - 0x3
    "00001111", --  530 - 0x212  :   15 - 0xf
    "00011111", --  531 - 0x213  :   31 - 0x1f
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "00110011", --  533 - 0x215  :   51 - 0x33
    "00100001", --  534 - 0x216  :   33 - 0x21
    "01100001", --  535 - 0x217  :   97 - 0x61
    "00000000", --  536 - 0x218  :    0 - 0x0
    "00000011", --  537 - 0x219  :    3 - 0x3
    "00001111", --  538 - 0x21a  :   15 - 0xf
    "00011111", --  539 - 0x21b  :   31 - 0x1f
    "00111111", --  540 - 0x21c  :   63 - 0x3f
    "00111111", --  541 - 0x21d  :   63 - 0x3f
    "00111111", --  542 - 0x21e  :   63 - 0x3f
    "01111111", --  543 - 0x21f  :  127 - 0x7f
    "01100001", --  544 - 0x220  :   97 - 0x61 -- Sprite 0x22
    "01110011", --  545 - 0x221  :  115 - 0x73
    "01111111", --  546 - 0x222  :  127 - 0x7f
    "01111111", --  547 - 0x223  :  127 - 0x7f
    "01101110", --  548 - 0x224  :  110 - 0x6e
    "01000110", --  549 - 0x225  :   70 - 0x46
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "01110011", --  552 - 0x228  :  115 - 0x73
    "01110011", --  553 - 0x229  :  115 - 0x73
    "01111111", --  554 - 0x22a  :  127 - 0x7f
    "01111111", --  555 - 0x22b  :  127 - 0x7f
    "01101110", --  556 - 0x22c  :  110 - 0x6e
    "01000110", --  557 - 0x22d  :   70 - 0x46
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "01100001", --  560 - 0x230  :   97 - 0x61 -- Sprite 0x23
    "01110011", --  561 - 0x231  :  115 - 0x73
    "01111111", --  562 - 0x232  :  127 - 0x7f
    "01111111", --  563 - 0x233  :  127 - 0x7f
    "01110111", --  564 - 0x234  :  119 - 0x77
    "00100011", --  565 - 0x235  :   35 - 0x23
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "01110011", --  568 - 0x238  :  115 - 0x73
    "01110011", --  569 - 0x239  :  115 - 0x73
    "01111111", --  570 - 0x23a  :  127 - 0x7f
    "01111111", --  571 - 0x23b  :  127 - 0x7f
    "01110111", --  572 - 0x23c  :  119 - 0x77
    "00100011", --  573 - 0x23d  :   35 - 0x23
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x24
    "00000011", --  577 - 0x241  :    3 - 0x3
    "00001111", --  578 - 0x242  :   15 - 0xf
    "00011111", --  579 - 0x243  :   31 - 0x1f
    "00111111", --  580 - 0x244  :   63 - 0x3f
    "00111111", --  581 - 0x245  :   63 - 0x3f
    "00111111", --  582 - 0x246  :   63 - 0x3f
    "01111111", --  583 - 0x247  :  127 - 0x7f
    "00000000", --  584 - 0x248  :    0 - 0x0
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000110", --  589 - 0x24d  :    6 - 0x6
    "00000110", --  590 - 0x24e  :    6 - 0x6
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "01111111", --  592 - 0x250  :  127 - 0x7f -- Sprite 0x25
    "01111111", --  593 - 0x251  :  127 - 0x7f
    "01111111", --  594 - 0x252  :  127 - 0x7f
    "01111111", --  595 - 0x253  :  127 - 0x7f
    "01101110", --  596 - 0x254  :  110 - 0x6e
    "01000110", --  597 - 0x255  :   70 - 0x46
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00011001", --  601 - 0x259  :   25 - 0x19
    "00100110", --  602 - 0x25a  :   38 - 0x26
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "01111111", --  608 - 0x260  :  127 - 0x7f -- Sprite 0x26
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "01111111", --  610 - 0x262  :  127 - 0x7f
    "01111111", --  611 - 0x263  :  127 - 0x7f
    "01111011", --  612 - 0x264  :  123 - 0x7b
    "00110001", --  613 - 0x265  :   49 - 0x31
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0
    "00011001", --  617 - 0x269  :   25 - 0x19
    "00100110", --  618 - 0x26a  :   38 - 0x26
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x27
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0
    "00001100", --  633 - 0x279  :   12 - 0xc
    "00010010", --  634 - 0x27a  :   18 - 0x12
    "00010010", --  635 - 0x27b  :   18 - 0x12
    "00011110", --  636 - 0x27c  :   30 - 0x1e
    "00001100", --  637 - 0x27d  :   12 - 0xc
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00111000", --  653 - 0x28d  :   56 - 0x38
    "01001101", --  654 - 0x28e  :   77 - 0x4d
    "01001101", --  655 - 0x28f  :   77 - 0x4d
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x29
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "11100000", --  669 - 0x29d  :  224 - 0xe0
    "00110000", --  670 - 0x29e  :   48 - 0x30
    "00110000", --  671 - 0x29f  :   48 - 0x30
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x2a
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00111000", --  680 - 0x2a8  :   56 - 0x38
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Sprite 0x2b
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "11100000", --  696 - 0x2b8  :  224 - 0xe0
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00001100", --  718 - 0x2ce  :   12 - 0xc
    "00011110", --  719 - 0x2cf  :   30 - 0x1e
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00010010", --  728 - 0x2d8  :   18 - 0x12
    "00010010", --  729 - 0x2d9  :   18 - 0x12
    "00001100", --  730 - 0x2da  :   12 - 0xc
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00010001", --  747 - 0x2eb  :   17 - 0x11
    "00110010", --  748 - 0x2ec  :   50 - 0x32
    "00010010", --  749 - 0x2ed  :   18 - 0x12
    "00010010", --  750 - 0x2ee  :   18 - 0x12
    "00010010", --  751 - 0x2ef  :   18 - 0x12
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "10001100", --  763 - 0x2fb  :  140 - 0x8c
    "01010010", --  764 - 0x2fc  :   82 - 0x52
    "01010010", --  765 - 0x2fd  :   82 - 0x52
    "01010010", --  766 - 0x2fe  :   82 - 0x52
    "01010010", --  767 - 0x2ff  :   82 - 0x52
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00010010", --  776 - 0x308  :   18 - 0x12
    "00111001", --  777 - 0x309  :   57 - 0x39
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x31
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "01010010", --  792 - 0x318  :   82 - 0x52
    "10001100", --  793 - 0x319  :  140 - 0x8c
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "01110001", --  811 - 0x32b  :  113 - 0x71
    "10001010", --  812 - 0x32c  :  138 - 0x8a
    "00001010", --  813 - 0x32d  :   10 - 0xa
    "00010010", --  814 - 0x32e  :   18 - 0x12
    "00100010", --  815 - 0x32f  :   34 - 0x22
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x33
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "01000010", --  824 - 0x338  :   66 - 0x42
    "11111001", --  825 - 0x339  :  249 - 0xf9
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00110001", --  843 - 0x34b  :   49 - 0x31
    "01001010", --  844 - 0x34c  :   74 - 0x4a
    "00001010", --  845 - 0x34d  :   10 - 0xa
    "00110010", --  846 - 0x34e  :   50 - 0x32
    "00001010", --  847 - 0x34f  :   10 - 0xa
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x35
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "01001010", --  856 - 0x358  :   74 - 0x4a
    "00110001", --  857 - 0x359  :   49 - 0x31
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00010001", --  875 - 0x36b  :   17 - 0x11
    "00110010", --  876 - 0x36c  :   50 - 0x32
    "01010010", --  877 - 0x36d  :   82 - 0x52
    "10010010", --  878 - 0x36e  :  146 - 0x92
    "11111010", --  879 - 0x36f  :  250 - 0xfa
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x37
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00010010", --  888 - 0x378  :   18 - 0x12
    "00010001", --  889 - 0x379  :   17 - 0x11
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "01110001", --  907 - 0x38b  :  113 - 0x71
    "01000010", --  908 - 0x38c  :   66 - 0x42
    "01000010", --  909 - 0x38d  :   66 - 0x42
    "01110010", --  910 - 0x38e  :  114 - 0x72
    "00001010", --  911 - 0x38f  :   10 - 0xa
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00001010", --  920 - 0x398  :   10 - 0xa
    "01110001", --  921 - 0x399  :  113 - 0x71
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "01110001", --  939 - 0x3ab  :  113 - 0x71
    "00001010", --  940 - 0x3ac  :   10 - 0xa
    "00010010", --  941 - 0x3ad  :   18 - 0x12
    "00010010", --  942 - 0x3ae  :   18 - 0x12
    "00100010", --  943 - 0x3af  :   34 - 0x22
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00100010", --  952 - 0x3b8  :   34 - 0x22
    "00100001", --  953 - 0x3b9  :   33 - 0x21
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "01110001", --  971 - 0x3cb  :  113 - 0x71
    "10001010", --  972 - 0x3cc  :  138 - 0x8a
    "10001010", --  973 - 0x3cd  :  138 - 0x8a
    "01110010", --  974 - 0x3ce  :  114 - 0x72
    "10001010", --  975 - 0x3cf  :  138 - 0x8a
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "10001010", --  984 - 0x3d8  :  138 - 0x8a
    "01110001", --  985 - 0x3d9  :  113 - 0x71
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "10011000", -- 1003 - 0x3eb  :  152 - 0x98
    "10100101", -- 1004 - 0x3ec  :  165 - 0xa5
    "10100101", -- 1005 - 0x3ed  :  165 - 0xa5
    "10100101", -- 1006 - 0x3ee  :  165 - 0xa5
    "10100101", -- 1007 - 0x3ef  :  165 - 0xa5
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "11000110", -- 1019 - 0x3fb  :  198 - 0xc6
    "00101001", -- 1020 - 0x3fc  :   41 - 0x29
    "00101001", -- 1021 - 0x3fd  :   41 - 0x29
    "00101001", -- 1022 - 0x3fe  :   41 - 0x29
    "00101001", -- 1023 - 0x3ff  :   41 - 0x29
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x40
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "10100101", -- 1032 - 0x408  :  165 - 0xa5
    "10011000", -- 1033 - 0x409  :  152 - 0x98
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x41
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00101001", -- 1048 - 0x418  :   41 - 0x29
    "11000110", -- 1049 - 0x419  :  198 - 0xc6
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Sprite 0x42
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "10011100", -- 1067 - 0x42b  :  156 - 0x9c
    "10100001", -- 1068 - 0x42c  :  161 - 0xa1
    "10100001", -- 1069 - 0x42d  :  161 - 0xa1
    "10111101", -- 1070 - 0x42e  :  189 - 0xbd
    "10100101", -- 1071 - 0x42f  :  165 - 0xa5
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x43
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "10100101", -- 1080 - 0x438  :  165 - 0xa5
    "10011000", -- 1081 - 0x439  :  152 - 0x98
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x44
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "01100010", -- 1099 - 0x44b  :   98 - 0x62
    "10010101", -- 1100 - 0x44c  :  149 - 0x95
    "00010101", -- 1101 - 0x44d  :   21 - 0x15
    "00100101", -- 1102 - 0x44e  :   37 - 0x25
    "01000101", -- 1103 - 0x44f  :   69 - 0x45
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x45
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00100010", -- 1115 - 0x45b  :   34 - 0x22
    "01010101", -- 1116 - 0x45c  :   85 - 0x55
    "01010101", -- 1117 - 0x45d  :   85 - 0x55
    "01010101", -- 1118 - 0x45e  :   85 - 0x55
    "01010101", -- 1119 - 0x45f  :   85 - 0x55
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x46
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "10000101", -- 1128 - 0x468  :  133 - 0x85
    "11110010", -- 1129 - 0x469  :  242 - 0xf2
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Sprite 0x47
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "01010101", -- 1144 - 0x478  :   85 - 0x55
    "00100010", -- 1145 - 0x479  :   34 - 0x22
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x48
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "01100010", -- 1163 - 0x48b  :   98 - 0x62
    "10010101", -- 1164 - 0x48c  :  149 - 0x95
    "00010101", -- 1165 - 0x48d  :   21 - 0x15
    "01100101", -- 1166 - 0x48e  :  101 - 0x65
    "00010101", -- 1167 - 0x48f  :   21 - 0x15
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x49
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "10010101", -- 1176 - 0x498  :  149 - 0x95
    "01100010", -- 1177 - 0x499  :   98 - 0x62
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x4a
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "11100010", -- 1195 - 0x4ab  :  226 - 0xe2
    "10000101", -- 1196 - 0x4ac  :  133 - 0x85
    "10000101", -- 1197 - 0x4ad  :  133 - 0x85
    "11100101", -- 1198 - 0x4ae  :  229 - 0xe5
    "00010101", -- 1199 - 0x4af  :   21 - 0x15
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x4b
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00010101", -- 1208 - 0x4b8  :   21 - 0x15
    "11100010", -- 1209 - 0x4b9  :  226 - 0xe2
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x4c
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x4d
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000001", -- 1235 - 0x4d3  :    1 - 0x1
    "00000011", -- 1236 - 0x4d4  :    3 - 0x3
    "00000111", -- 1237 - 0x4d5  :    7 - 0x7
    "00001111", -- 1238 - 0x4d6  :   15 - 0xf
    "00011111", -- 1239 - 0x4d7  :   31 - 0x1f
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Sprite 0x4e
    "00001111", -- 1249 - 0x4e1  :   15 - 0xf
    "01111111", -- 1250 - 0x4e2  :  127 - 0x7f
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111111", -- 1254 - 0x4e6  :  255 - 0xff
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00011111", -- 1264 - 0x4f0  :   31 - 0x1f -- Sprite 0x4f
    "00111111", -- 1265 - 0x4f1  :   63 - 0x3f
    "00111111", -- 1266 - 0x4f2  :   63 - 0x3f
    "00111111", -- 1267 - 0x4f3  :   63 - 0x3f
    "01111111", -- 1268 - 0x4f4  :  127 - 0x7f
    "01111111", -- 1269 - 0x4f5  :  127 - 0x7f
    "01111111", -- 1270 - 0x4f6  :  127 - 0x7f
    "01111111", -- 1271 - 0x4f7  :  127 - 0x7f
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0x50
    "11111111", -- 1281 - 0x501  :  255 - 0xff
    "11111111", -- 1282 - 0x502  :  255 - 0xff
    "11111111", -- 1283 - 0x503  :  255 - 0xff
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Sprite 0x51
    "11111111", -- 1297 - 0x511  :  255 - 0xff
    "11111111", -- 1298 - 0x512  :  255 - 0xff
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "11111111", -- 1300 - 0x514  :  255 - 0xff
    "11111111", -- 1301 - 0x515  :  255 - 0xff
    "11111111", -- 1302 - 0x516  :  255 - 0xff
    "11111110", -- 1303 - 0x517  :  254 - 0xfe
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0x52
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "10000000", -- 1315 - 0x523  :  128 - 0x80
    "11000000", -- 1316 - 0x524  :  192 - 0xc0
    "11100000", -- 1317 - 0x525  :  224 - 0xe0
    "11110000", -- 1318 - 0x526  :  240 - 0xf0
    "11110000", -- 1319 - 0x527  :  240 - 0xf0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Sprite 0x53
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "11111110", -- 1330 - 0x532  :  254 - 0xfe
    "11111100", -- 1331 - 0x533  :  252 - 0xfc
    "11110000", -- 1332 - 0x534  :  240 - 0xf0
    "11100000", -- 1333 - 0x535  :  224 - 0xe0
    "10000000", -- 1334 - 0x536  :  128 - 0x80
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "11000000", -- 1344 - 0x540  :  192 - 0xc0 -- Sprite 0x54
    "10000000", -- 1345 - 0x541  :  128 - 0x80
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0x55
    "11110000", -- 1361 - 0x551  :  240 - 0xf0
    "11111110", -- 1362 - 0x552  :  254 - 0xfe
    "11111110", -- 1363 - 0x553  :  254 - 0xfe
    "11111110", -- 1364 - 0x554  :  254 - 0xfe
    "11111100", -- 1365 - 0x555  :  252 - 0xfc
    "11111000", -- 1366 - 0x556  :  248 - 0xf8
    "11111000", -- 1367 - 0x557  :  248 - 0xf8
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "11110000", -- 1376 - 0x560  :  240 - 0xf0 -- Sprite 0x56
    "11100000", -- 1377 - 0x561  :  224 - 0xe0
    "11100000", -- 1378 - 0x562  :  224 - 0xe0
    "11000000", -- 1379 - 0x563  :  192 - 0xc0
    "10000000", -- 1380 - 0x564  :  128 - 0x80
    "10000000", -- 1381 - 0x565  :  128 - 0x80
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0x57
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000100", -- 1399 - 0x577  :    4 - 0x4
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000100", -- 1407 - 0x57f  :    4 - 0x4
    "00000110", -- 1408 - 0x580  :    6 - 0x6 -- Sprite 0x58
    "00000110", -- 1409 - 0x581  :    6 - 0x6
    "00000111", -- 1410 - 0x582  :    7 - 0x7
    "00000111", -- 1411 - 0x583  :    7 - 0x7
    "00000111", -- 1412 - 0x584  :    7 - 0x7
    "00000111", -- 1413 - 0x585  :    7 - 0x7
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000110", -- 1416 - 0x588  :    6 - 0x6
    "00000110", -- 1417 - 0x589  :    6 - 0x6
    "00000111", -- 1418 - 0x58a  :    7 - 0x7
    "00000111", -- 1419 - 0x58b  :    7 - 0x7
    "00000111", -- 1420 - 0x58c  :    7 - 0x7
    "00000111", -- 1421 - 0x58d  :    7 - 0x7
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0x59
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00010000", -- 1431 - 0x597  :   16 - 0x10
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00010000", -- 1439 - 0x59f  :   16 - 0x10
    "00011100", -- 1440 - 0x5a0  :   28 - 0x1c -- Sprite 0x5a
    "00011110", -- 1441 - 0x5a1  :   30 - 0x1e
    "00011111", -- 1442 - 0x5a2  :   31 - 0x1f
    "00011111", -- 1443 - 0x5a3  :   31 - 0x1f
    "00011111", -- 1444 - 0x5a4  :   31 - 0x1f
    "00011111", -- 1445 - 0x5a5  :   31 - 0x1f
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00011100", -- 1448 - 0x5a8  :   28 - 0x1c
    "00011110", -- 1449 - 0x5a9  :   30 - 0x1e
    "00011111", -- 1450 - 0x5aa  :   31 - 0x1f
    "00011111", -- 1451 - 0x5ab  :   31 - 0x1f
    "00011111", -- 1452 - 0x5ac  :   31 - 0x1f
    "00011111", -- 1453 - 0x5ad  :   31 - 0x1f
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "11000000", -- 1463 - 0x5b7  :  192 - 0xc0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "11000000", -- 1471 - 0x5bf  :  192 - 0xc0
    "11110000", -- 1472 - 0x5c0  :  240 - 0xf0 -- Sprite 0x5c
    "11111100", -- 1473 - 0x5c1  :  252 - 0xfc
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "11110000", -- 1480 - 0x5c8  :  240 - 0xf0
    "11111100", -- 1481 - 0x5c9  :  252 - 0xfc
    "11111111", -- 1482 - 0x5ca  :  255 - 0xff
    "11111111", -- 1483 - 0x5cb  :  255 - 0xff
    "11111111", -- 1484 - 0x5cc  :  255 - 0xff
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0x5d
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000001", -- 1490 - 0x5d2  :    1 - 0x1
    "00000011", -- 1491 - 0x5d3  :    3 - 0x3
    "00001111", -- 1492 - 0x5d4  :   15 - 0xf
    "00001111", -- 1493 - 0x5d5  :   15 - 0xf
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000001", -- 1498 - 0x5da  :    1 - 0x1
    "00000011", -- 1499 - 0x5db  :    3 - 0x3
    "00001111", -- 1500 - 0x5dc  :   15 - 0xf
    "00001111", -- 1501 - 0x5dd  :   15 - 0xf
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "11111100", -- 1504 - 0x5e0  :  252 - 0xfc -- Sprite 0x5e
    "11111100", -- 1505 - 0x5e1  :  252 - 0xfc
    "11111100", -- 1506 - 0x5e2  :  252 - 0xfc
    "11111100", -- 1507 - 0x5e3  :  252 - 0xfc
    "11111000", -- 1508 - 0x5e4  :  248 - 0xf8
    "11111100", -- 1509 - 0x5e5  :  252 - 0xfc
    "00111100", -- 1510 - 0x5e6  :   60 - 0x3c
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "11111000", -- 1512 - 0x5e8  :  248 - 0xf8
    "11110000", -- 1513 - 0x5e9  :  240 - 0xf0
    "11100000", -- 1514 - 0x5ea  :  224 - 0xe0
    "11110000", -- 1515 - 0x5eb  :  240 - 0xf0
    "11100000", -- 1516 - 0x5ec  :  224 - 0xe0
    "11000000", -- 1517 - 0x5ed  :  192 - 0xc0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000100", -- 1520 - 0x5f0  :    4 - 0x4 -- Sprite 0x5f
    "00001100", -- 1521 - 0x5f1  :   12 - 0xc
    "00011100", -- 1522 - 0x5f2  :   28 - 0x1c
    "00001100", -- 1523 - 0x5f3  :   12 - 0xc
    "00011000", -- 1524 - 0x5f4  :   24 - 0x18
    "00111100", -- 1525 - 0x5f5  :   60 - 0x3c
    "00111100", -- 1526 - 0x5f6  :   60 - 0x3c
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000011", -- 1537 - 0x601  :    3 - 0x3
    "00001111", -- 1538 - 0x602  :   15 - 0xf
    "00010011", -- 1539 - 0x603  :   19 - 0x13
    "00100001", -- 1540 - 0x604  :   33 - 0x21
    "00100001", -- 1541 - 0x605  :   33 - 0x21
    "00100001", -- 1542 - 0x606  :   33 - 0x21
    "01110011", -- 1543 - 0x607  :  115 - 0x73
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000011", -- 1545 - 0x609  :    3 - 0x3
    "00001111", -- 1546 - 0x60a  :   15 - 0xf
    "00011111", -- 1547 - 0x60b  :   31 - 0x1f
    "00111111", -- 1548 - 0x60c  :   63 - 0x3f
    "00111111", -- 1549 - 0x60d  :   63 - 0x3f
    "00111001", -- 1550 - 0x60e  :   57 - 0x39
    "01111011", -- 1551 - 0x60f  :  123 - 0x7b
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0x61
    "11000000", -- 1553 - 0x611  :  192 - 0xc0
    "11110000", -- 1554 - 0x612  :  240 - 0xf0
    "11001000", -- 1555 - 0x613  :  200 - 0xc8
    "10000100", -- 1556 - 0x614  :  132 - 0x84
    "10000100", -- 1557 - 0x615  :  132 - 0x84
    "10000100", -- 1558 - 0x616  :  132 - 0x84
    "11001110", -- 1559 - 0x617  :  206 - 0xce
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "11000000", -- 1561 - 0x619  :  192 - 0xc0
    "11110000", -- 1562 - 0x61a  :  240 - 0xf0
    "11111000", -- 1563 - 0x61b  :  248 - 0xf8
    "11111100", -- 1564 - 0x61c  :  252 - 0xfc
    "11111100", -- 1565 - 0x61d  :  252 - 0xfc
    "11100100", -- 1566 - 0x61e  :  228 - 0xe4
    "11101110", -- 1567 - 0x61f  :  238 - 0xee
    "10010100", -- 1568 - 0x620  :  148 - 0x94 -- Sprite 0x62
    "11101010", -- 1569 - 0x621  :  234 - 0xea
    "11011110", -- 1570 - 0x622  :  222 - 0xde
    "11101110", -- 1571 - 0x623  :  238 - 0xee
    "11011110", -- 1572 - 0x624  :  222 - 0xde
    "01100110", -- 1573 - 0x625  :  102 - 0x66
    "01000010", -- 1574 - 0x626  :   66 - 0x42
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "11111110", -- 1576 - 0x628  :  254 - 0xfe
    "11111110", -- 1577 - 0x629  :  254 - 0xfe
    "11111110", -- 1578 - 0x62a  :  254 - 0xfe
    "11111110", -- 1579 - 0x62b  :  254 - 0xfe
    "11111110", -- 1580 - 0x62c  :  254 - 0xfe
    "01100110", -- 1581 - 0x62d  :  102 - 0x66
    "01000010", -- 1582 - 0x62e  :   66 - 0x42
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "10010100", -- 1584 - 0x630  :  148 - 0x94 -- Sprite 0x63
    "11101010", -- 1585 - 0x631  :  234 - 0xea
    "11011110", -- 1586 - 0x632  :  222 - 0xde
    "11101110", -- 1587 - 0x633  :  238 - 0xee
    "11011110", -- 1588 - 0x634  :  222 - 0xde
    "11001110", -- 1589 - 0x635  :  206 - 0xce
    "10001100", -- 1590 - 0x636  :  140 - 0x8c
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "11111110", -- 1592 - 0x638  :  254 - 0xfe
    "11111110", -- 1593 - 0x639  :  254 - 0xfe
    "11111110", -- 1594 - 0x63a  :  254 - 0xfe
    "11111110", -- 1595 - 0x63b  :  254 - 0xfe
    "11111110", -- 1596 - 0x63c  :  254 - 0xfe
    "11011110", -- 1597 - 0x63d  :  222 - 0xde
    "10001100", -- 1598 - 0x63e  :  140 - 0x8c
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000001", -- 1607 - 0x647  :    1 - 0x1
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00110110", -- 1621 - 0x655  :   54 - 0x36
    "00110110", -- 1622 - 0x656  :   54 - 0x36
    "10010000", -- 1623 - 0x657  :  144 - 0x90
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "01101100", -- 1628 - 0x65c  :  108 - 0x6c
    "11111110", -- 1629 - 0x65d  :  254 - 0xfe
    "11111110", -- 1630 - 0x65e  :  254 - 0xfe
    "11111100", -- 1631 - 0x65f  :  252 - 0xfc
    "00000001", -- 1632 - 0x660  :    1 - 0x1 -- Sprite 0x66
    "00000011", -- 1633 - 0x661  :    3 - 0x3
    "00000111", -- 1634 - 0x662  :    7 - 0x7
    "00000111", -- 1635 - 0x663  :    7 - 0x7
    "00011111", -- 1636 - 0x664  :   31 - 0x1f
    "00011111", -- 1637 - 0x665  :   31 - 0x1f
    "00011100", -- 1638 - 0x666  :   28 - 0x1c
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11111000", -- 1648 - 0x670  :  248 - 0xf8 -- Sprite 0x67
    "11111000", -- 1649 - 0x671  :  248 - 0xf8
    "11111000", -- 1650 - 0x672  :  248 - 0xf8
    "11111000", -- 1651 - 0x673  :  248 - 0xf8
    "11111110", -- 1652 - 0x674  :  254 - 0xfe
    "11111110", -- 1653 - 0x675  :  254 - 0xfe
    "00001110", -- 1654 - 0x676  :   14 - 0xe
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000111", -- 1664 - 0x680  :    7 - 0x7 -- Sprite 0x68
    "00001111", -- 1665 - 0x681  :   15 - 0xf
    "00011111", -- 1666 - 0x682  :   31 - 0x1f
    "00011111", -- 1667 - 0x683  :   31 - 0x1f
    "00111111", -- 1668 - 0x684  :   63 - 0x3f
    "00111111", -- 1669 - 0x685  :   63 - 0x3f
    "00111000", -- 1670 - 0x686  :   56 - 0x38
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "11111000", -- 1680 - 0x690  :  248 - 0xf8 -- Sprite 0x69
    "11110000", -- 1681 - 0x691  :  240 - 0xf0
    "11110000", -- 1682 - 0x692  :  240 - 0xf0
    "11100000", -- 1683 - 0x693  :  224 - 0xe0
    "11111000", -- 1684 - 0x694  :  248 - 0xf8
    "11111000", -- 1685 - 0x695  :  248 - 0xf8
    "00111000", -- 1686 - 0x696  :   56 - 0x38
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "00011111", -- 1697 - 0x6a1  :   31 - 0x1f
    "01111111", -- 1698 - 0x6a2  :  127 - 0x7f
    "00111111", -- 1699 - 0x6a3  :   63 - 0x3f
    "00001111", -- 1700 - 0x6a4  :   15 - 0xf
    "00000111", -- 1701 - 0x6a5  :    7 - 0x7
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00011111", -- 1705 - 0x6a9  :   31 - 0x1f
    "01111111", -- 1706 - 0x6aa  :  127 - 0x7f
    "00111111", -- 1707 - 0x6ab  :   63 - 0x3f
    "00001111", -- 1708 - 0x6ac  :   15 - 0xf
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0x6b
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "11000000", -- 1714 - 0x6b2  :  192 - 0xc0
    "11110000", -- 1715 - 0x6b3  :  240 - 0xf0
    "11111000", -- 1716 - 0x6b4  :  248 - 0xf8
    "11111000", -- 1717 - 0x6b5  :  248 - 0xf8
    "11100000", -- 1718 - 0x6b6  :  224 - 0xe0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "11000000", -- 1722 - 0x6ba  :  192 - 0xc0
    "11110000", -- 1723 - 0x6bb  :  240 - 0xf0
    "11111000", -- 1724 - 0x6bc  :  248 - 0xf8
    "11111000", -- 1725 - 0x6bd  :  248 - 0xf8
    "11100000", -- 1726 - 0x6be  :  224 - 0xe0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0x6c
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0x6d
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0x6f
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "11111111", -- 1792 - 0x700  :  255 - 0xff -- Sprite 0x70
    "11111111", -- 1793 - 0x701  :  255 - 0xff
    "11111111", -- 1794 - 0x702  :  255 - 0xff
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "11111111", -- 1796 - 0x704  :  255 - 0xff
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "11111111", -- 1802 - 0x70a  :  255 - 0xff
    "11111111", -- 1803 - 0x70b  :  255 - 0xff
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Sprite 0x71
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11111111", -- 1816 - 0x718  :  255 - 0xff
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "11111111", -- 1818 - 0x71a  :  255 - 0xff
    "11111111", -- 1819 - 0x71b  :  255 - 0xff
    "11111111", -- 1820 - 0x71c  :  255 - 0xff
    "11111111", -- 1821 - 0x71d  :  255 - 0xff
    "11111111", -- 1822 - 0x71e  :  255 - 0xff
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "11111111", -- 1824 - 0x720  :  255 - 0xff -- Sprite 0x72
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "11111111", -- 1826 - 0x722  :  255 - 0xff
    "11111111", -- 1827 - 0x723  :  255 - 0xff
    "11111111", -- 1828 - 0x724  :  255 - 0xff
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "11111111", -- 1834 - 0x72a  :  255 - 0xff
    "11111111", -- 1835 - 0x72b  :  255 - 0xff
    "11111111", -- 1836 - 0x72c  :  255 - 0xff
    "11111111", -- 1837 - 0x72d  :  255 - 0xff
    "11111111", -- 1838 - 0x72e  :  255 - 0xff
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Sprite 0x73
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11111111", -- 1843 - 0x733  :  255 - 0xff
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11111111", -- 1845 - 0x735  :  255 - 0xff
    "11111111", -- 1846 - 0x736  :  255 - 0xff
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "11111111", -- 1850 - 0x73a  :  255 - 0xff
    "11111111", -- 1851 - 0x73b  :  255 - 0xff
    "11111111", -- 1852 - 0x73c  :  255 - 0xff
    "11111111", -- 1853 - 0x73d  :  255 - 0xff
    "11111111", -- 1854 - 0x73e  :  255 - 0xff
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0x74
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11111111", -- 1864 - 0x748  :  255 - 0xff
    "11111111", -- 1865 - 0x749  :  255 - 0xff
    "11111111", -- 1866 - 0x74a  :  255 - 0xff
    "11111111", -- 1867 - 0x74b  :  255 - 0xff
    "11111111", -- 1868 - 0x74c  :  255 - 0xff
    "11111111", -- 1869 - 0x74d  :  255 - 0xff
    "11111111", -- 1870 - 0x74e  :  255 - 0xff
    "11111111", -- 1871 - 0x74f  :  255 - 0xff
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0x75
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "11111111", -- 1880 - 0x758  :  255 - 0xff
    "11111111", -- 1881 - 0x759  :  255 - 0xff
    "11111111", -- 1882 - 0x75a  :  255 - 0xff
    "11111111", -- 1883 - 0x75b  :  255 - 0xff
    "11111111", -- 1884 - 0x75c  :  255 - 0xff
    "11111111", -- 1885 - 0x75d  :  255 - 0xff
    "11111111", -- 1886 - 0x75e  :  255 - 0xff
    "11111111", -- 1887 - 0x75f  :  255 - 0xff
    "11111111", -- 1888 - 0x760  :  255 - 0xff -- Sprite 0x76
    "11111111", -- 1889 - 0x761  :  255 - 0xff
    "11111111", -- 1890 - 0x762  :  255 - 0xff
    "11111111", -- 1891 - 0x763  :  255 - 0xff
    "11111111", -- 1892 - 0x764  :  255 - 0xff
    "11111111", -- 1893 - 0x765  :  255 - 0xff
    "11111111", -- 1894 - 0x766  :  255 - 0xff
    "11111111", -- 1895 - 0x767  :  255 - 0xff
    "11111111", -- 1896 - 0x768  :  255 - 0xff
    "11111111", -- 1897 - 0x769  :  255 - 0xff
    "11111111", -- 1898 - 0x76a  :  255 - 0xff
    "11111111", -- 1899 - 0x76b  :  255 - 0xff
    "11111111", -- 1900 - 0x76c  :  255 - 0xff
    "11111111", -- 1901 - 0x76d  :  255 - 0xff
    "11111111", -- 1902 - 0x76e  :  255 - 0xff
    "11111111", -- 1903 - 0x76f  :  255 - 0xff
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Sprite 0x77
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "11111111", -- 1906 - 0x772  :  255 - 0xff
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111111", -- 1909 - 0x775  :  255 - 0xff
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "11111111", -- 1912 - 0x778  :  255 - 0xff
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111111", -- 1914 - 0x77a  :  255 - 0xff
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111111", -- 1916 - 0x77c  :  255 - 0xff
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11111111", -- 1919 - 0x77f  :  255 - 0xff
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0x78
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0x79
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "11111111", -- 1944 - 0x798  :  255 - 0xff
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Sprite 0x7a
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Sprite 0x7b
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0x7c
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0x7d
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Sprite 0x7e
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff
    "11111111", -- 2025 - 0x7e9  :  255 - 0xff
    "11111111", -- 2026 - 0x7ea  :  255 - 0xff
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111111", -- 2028 - 0x7ec  :  255 - 0xff
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Sprite 0x7f
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111", -- 2047 - 0x7ff  :  255 - 0xff
    "11111111", -- 2048 - 0x800  :  255 - 0xff -- Sprite 0x80
    "11111111", -- 2049 - 0x801  :  255 - 0xff
    "11111111", -- 2050 - 0x802  :  255 - 0xff
    "11111111", -- 2051 - 0x803  :  255 - 0xff
    "11111111", -- 2052 - 0x804  :  255 - 0xff
    "11111111", -- 2053 - 0x805  :  255 - 0xff
    "11111111", -- 2054 - 0x806  :  255 - 0xff
    "11111111", -- 2055 - 0x807  :  255 - 0xff
    "11111111", -- 2056 - 0x808  :  255 - 0xff
    "11111111", -- 2057 - 0x809  :  255 - 0xff
    "11111111", -- 2058 - 0x80a  :  255 - 0xff
    "11111111", -- 2059 - 0x80b  :  255 - 0xff
    "11111111", -- 2060 - 0x80c  :  255 - 0xff
    "11111111", -- 2061 - 0x80d  :  255 - 0xff
    "11111111", -- 2062 - 0x80e  :  255 - 0xff
    "11111111", -- 2063 - 0x80f  :  255 - 0xff
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Sprite 0x81
    "11111111", -- 2065 - 0x811  :  255 - 0xff
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "11111111", -- 2067 - 0x813  :  255 - 0xff
    "11111111", -- 2068 - 0x814  :  255 - 0xff
    "11111111", -- 2069 - 0x815  :  255 - 0xff
    "11111111", -- 2070 - 0x816  :  255 - 0xff
    "11111111", -- 2071 - 0x817  :  255 - 0xff
    "11111111", -- 2072 - 0x818  :  255 - 0xff
    "11111111", -- 2073 - 0x819  :  255 - 0xff
    "11111111", -- 2074 - 0x81a  :  255 - 0xff
    "11111111", -- 2075 - 0x81b  :  255 - 0xff
    "11111111", -- 2076 - 0x81c  :  255 - 0xff
    "11111111", -- 2077 - 0x81d  :  255 - 0xff
    "11111111", -- 2078 - 0x81e  :  255 - 0xff
    "11111111", -- 2079 - 0x81f  :  255 - 0xff
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Sprite 0x82
    "11111111", -- 2081 - 0x821  :  255 - 0xff
    "11111111", -- 2082 - 0x822  :  255 - 0xff
    "11111111", -- 2083 - 0x823  :  255 - 0xff
    "11111111", -- 2084 - 0x824  :  255 - 0xff
    "11111111", -- 2085 - 0x825  :  255 - 0xff
    "11111111", -- 2086 - 0x826  :  255 - 0xff
    "11111111", -- 2087 - 0x827  :  255 - 0xff
    "11111111", -- 2088 - 0x828  :  255 - 0xff
    "11111111", -- 2089 - 0x829  :  255 - 0xff
    "11111111", -- 2090 - 0x82a  :  255 - 0xff
    "11111111", -- 2091 - 0x82b  :  255 - 0xff
    "11111111", -- 2092 - 0x82c  :  255 - 0xff
    "11111111", -- 2093 - 0x82d  :  255 - 0xff
    "11111111", -- 2094 - 0x82e  :  255 - 0xff
    "11111111", -- 2095 - 0x82f  :  255 - 0xff
    "11111111", -- 2096 - 0x830  :  255 - 0xff -- Sprite 0x83
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "11111111", -- 2098 - 0x832  :  255 - 0xff
    "11111111", -- 2099 - 0x833  :  255 - 0xff
    "11111111", -- 2100 - 0x834  :  255 - 0xff
    "11111111", -- 2101 - 0x835  :  255 - 0xff
    "11111111", -- 2102 - 0x836  :  255 - 0xff
    "11111111", -- 2103 - 0x837  :  255 - 0xff
    "11111111", -- 2104 - 0x838  :  255 - 0xff
    "11111111", -- 2105 - 0x839  :  255 - 0xff
    "11111111", -- 2106 - 0x83a  :  255 - 0xff
    "11111111", -- 2107 - 0x83b  :  255 - 0xff
    "11111111", -- 2108 - 0x83c  :  255 - 0xff
    "11111111", -- 2109 - 0x83d  :  255 - 0xff
    "11111111", -- 2110 - 0x83e  :  255 - 0xff
    "11111111", -- 2111 - 0x83f  :  255 - 0xff
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Sprite 0x84
    "11111111", -- 2113 - 0x841  :  255 - 0xff
    "11111111", -- 2114 - 0x842  :  255 - 0xff
    "11111111", -- 2115 - 0x843  :  255 - 0xff
    "11111111", -- 2116 - 0x844  :  255 - 0xff
    "11111111", -- 2117 - 0x845  :  255 - 0xff
    "11111111", -- 2118 - 0x846  :  255 - 0xff
    "11111111", -- 2119 - 0x847  :  255 - 0xff
    "11111111", -- 2120 - 0x848  :  255 - 0xff
    "11111111", -- 2121 - 0x849  :  255 - 0xff
    "11111111", -- 2122 - 0x84a  :  255 - 0xff
    "11111111", -- 2123 - 0x84b  :  255 - 0xff
    "11111111", -- 2124 - 0x84c  :  255 - 0xff
    "11111111", -- 2125 - 0x84d  :  255 - 0xff
    "11111111", -- 2126 - 0x84e  :  255 - 0xff
    "11111111", -- 2127 - 0x84f  :  255 - 0xff
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Sprite 0x85
    "11111111", -- 2129 - 0x851  :  255 - 0xff
    "11111111", -- 2130 - 0x852  :  255 - 0xff
    "11111111", -- 2131 - 0x853  :  255 - 0xff
    "11111111", -- 2132 - 0x854  :  255 - 0xff
    "11111111", -- 2133 - 0x855  :  255 - 0xff
    "11111111", -- 2134 - 0x856  :  255 - 0xff
    "11111111", -- 2135 - 0x857  :  255 - 0xff
    "11111111", -- 2136 - 0x858  :  255 - 0xff
    "11111111", -- 2137 - 0x859  :  255 - 0xff
    "11111111", -- 2138 - 0x85a  :  255 - 0xff
    "11111111", -- 2139 - 0x85b  :  255 - 0xff
    "11111111", -- 2140 - 0x85c  :  255 - 0xff
    "11111111", -- 2141 - 0x85d  :  255 - 0xff
    "11111111", -- 2142 - 0x85e  :  255 - 0xff
    "11111111", -- 2143 - 0x85f  :  255 - 0xff
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11111111", -- 2147 - 0x863  :  255 - 0xff
    "11111111", -- 2148 - 0x864  :  255 - 0xff
    "11111111", -- 2149 - 0x865  :  255 - 0xff
    "11111111", -- 2150 - 0x866  :  255 - 0xff
    "11111111", -- 2151 - 0x867  :  255 - 0xff
    "11111111", -- 2152 - 0x868  :  255 - 0xff
    "11111111", -- 2153 - 0x869  :  255 - 0xff
    "11111111", -- 2154 - 0x86a  :  255 - 0xff
    "11111111", -- 2155 - 0x86b  :  255 - 0xff
    "11111111", -- 2156 - 0x86c  :  255 - 0xff
    "11111111", -- 2157 - 0x86d  :  255 - 0xff
    "11111111", -- 2158 - 0x86e  :  255 - 0xff
    "11111111", -- 2159 - 0x86f  :  255 - 0xff
    "11111111", -- 2160 - 0x870  :  255 - 0xff -- Sprite 0x87
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "11111111", -- 2165 - 0x875  :  255 - 0xff
    "11111111", -- 2166 - 0x876  :  255 - 0xff
    "11111111", -- 2167 - 0x877  :  255 - 0xff
    "11111111", -- 2168 - 0x878  :  255 - 0xff
    "11111111", -- 2169 - 0x879  :  255 - 0xff
    "11111111", -- 2170 - 0x87a  :  255 - 0xff
    "11111111", -- 2171 - 0x87b  :  255 - 0xff
    "11111111", -- 2172 - 0x87c  :  255 - 0xff
    "11111111", -- 2173 - 0x87d  :  255 - 0xff
    "11111111", -- 2174 - 0x87e  :  255 - 0xff
    "11111111", -- 2175 - 0x87f  :  255 - 0xff
    "11111111", -- 2176 - 0x880  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "11111111", -- 2178 - 0x882  :  255 - 0xff
    "11111111", -- 2179 - 0x883  :  255 - 0xff
    "11111111", -- 2180 - 0x884  :  255 - 0xff
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "11111111", -- 2182 - 0x886  :  255 - 0xff
    "11111111", -- 2183 - 0x887  :  255 - 0xff
    "11111111", -- 2184 - 0x888  :  255 - 0xff
    "11111111", -- 2185 - 0x889  :  255 - 0xff
    "11111111", -- 2186 - 0x88a  :  255 - 0xff
    "11111111", -- 2187 - 0x88b  :  255 - 0xff
    "11111111", -- 2188 - 0x88c  :  255 - 0xff
    "11111111", -- 2189 - 0x88d  :  255 - 0xff
    "11111111", -- 2190 - 0x88e  :  255 - 0xff
    "11111111", -- 2191 - 0x88f  :  255 - 0xff
    "11111111", -- 2192 - 0x890  :  255 - 0xff -- Sprite 0x89
    "11111111", -- 2193 - 0x891  :  255 - 0xff
    "11111111", -- 2194 - 0x892  :  255 - 0xff
    "11111111", -- 2195 - 0x893  :  255 - 0xff
    "11111111", -- 2196 - 0x894  :  255 - 0xff
    "11111111", -- 2197 - 0x895  :  255 - 0xff
    "11111111", -- 2198 - 0x896  :  255 - 0xff
    "11111111", -- 2199 - 0x897  :  255 - 0xff
    "11111111", -- 2200 - 0x898  :  255 - 0xff
    "11111111", -- 2201 - 0x899  :  255 - 0xff
    "11111111", -- 2202 - 0x89a  :  255 - 0xff
    "11111111", -- 2203 - 0x89b  :  255 - 0xff
    "11111111", -- 2204 - 0x89c  :  255 - 0xff
    "11111111", -- 2205 - 0x89d  :  255 - 0xff
    "11111111", -- 2206 - 0x89e  :  255 - 0xff
    "11111111", -- 2207 - 0x89f  :  255 - 0xff
    "11111111", -- 2208 - 0x8a0  :  255 - 0xff -- Sprite 0x8a
    "11111111", -- 2209 - 0x8a1  :  255 - 0xff
    "11111111", -- 2210 - 0x8a2  :  255 - 0xff
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "11111111", -- 2212 - 0x8a4  :  255 - 0xff
    "11111111", -- 2213 - 0x8a5  :  255 - 0xff
    "11111111", -- 2214 - 0x8a6  :  255 - 0xff
    "11111111", -- 2215 - 0x8a7  :  255 - 0xff
    "11111111", -- 2216 - 0x8a8  :  255 - 0xff
    "11111111", -- 2217 - 0x8a9  :  255 - 0xff
    "11111111", -- 2218 - 0x8aa  :  255 - 0xff
    "11111111", -- 2219 - 0x8ab  :  255 - 0xff
    "11111111", -- 2220 - 0x8ac  :  255 - 0xff
    "11111111", -- 2221 - 0x8ad  :  255 - 0xff
    "11111111", -- 2222 - 0x8ae  :  255 - 0xff
    "11111111", -- 2223 - 0x8af  :  255 - 0xff
    "11111111", -- 2224 - 0x8b0  :  255 - 0xff -- Sprite 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11111111", -- 2226 - 0x8b2  :  255 - 0xff
    "11111111", -- 2227 - 0x8b3  :  255 - 0xff
    "11111111", -- 2228 - 0x8b4  :  255 - 0xff
    "11111111", -- 2229 - 0x8b5  :  255 - 0xff
    "11111111", -- 2230 - 0x8b6  :  255 - 0xff
    "11111111", -- 2231 - 0x8b7  :  255 - 0xff
    "11111111", -- 2232 - 0x8b8  :  255 - 0xff
    "11111111", -- 2233 - 0x8b9  :  255 - 0xff
    "11111111", -- 2234 - 0x8ba  :  255 - 0xff
    "11111111", -- 2235 - 0x8bb  :  255 - 0xff
    "11111111", -- 2236 - 0x8bc  :  255 - 0xff
    "11111111", -- 2237 - 0x8bd  :  255 - 0xff
    "11111111", -- 2238 - 0x8be  :  255 - 0xff
    "11111111", -- 2239 - 0x8bf  :  255 - 0xff
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Sprite 0x8c
    "11111111", -- 2241 - 0x8c1  :  255 - 0xff
    "11111111", -- 2242 - 0x8c2  :  255 - 0xff
    "11111111", -- 2243 - 0x8c3  :  255 - 0xff
    "11111111", -- 2244 - 0x8c4  :  255 - 0xff
    "11111111", -- 2245 - 0x8c5  :  255 - 0xff
    "11111111", -- 2246 - 0x8c6  :  255 - 0xff
    "11111111", -- 2247 - 0x8c7  :  255 - 0xff
    "11111111", -- 2248 - 0x8c8  :  255 - 0xff
    "11111111", -- 2249 - 0x8c9  :  255 - 0xff
    "11111111", -- 2250 - 0x8ca  :  255 - 0xff
    "11111111", -- 2251 - 0x8cb  :  255 - 0xff
    "11111111", -- 2252 - 0x8cc  :  255 - 0xff
    "11111111", -- 2253 - 0x8cd  :  255 - 0xff
    "11111111", -- 2254 - 0x8ce  :  255 - 0xff
    "11111111", -- 2255 - 0x8cf  :  255 - 0xff
    "11111111", -- 2256 - 0x8d0  :  255 - 0xff -- Sprite 0x8d
    "11111111", -- 2257 - 0x8d1  :  255 - 0xff
    "11111111", -- 2258 - 0x8d2  :  255 - 0xff
    "11111111", -- 2259 - 0x8d3  :  255 - 0xff
    "11111111", -- 2260 - 0x8d4  :  255 - 0xff
    "11111111", -- 2261 - 0x8d5  :  255 - 0xff
    "11111111", -- 2262 - 0x8d6  :  255 - 0xff
    "11111111", -- 2263 - 0x8d7  :  255 - 0xff
    "11111111", -- 2264 - 0x8d8  :  255 - 0xff
    "11111111", -- 2265 - 0x8d9  :  255 - 0xff
    "11111111", -- 2266 - 0x8da  :  255 - 0xff
    "11111111", -- 2267 - 0x8db  :  255 - 0xff
    "11111111", -- 2268 - 0x8dc  :  255 - 0xff
    "11111111", -- 2269 - 0x8dd  :  255 - 0xff
    "11111111", -- 2270 - 0x8de  :  255 - 0xff
    "11111111", -- 2271 - 0x8df  :  255 - 0xff
    "11111111", -- 2272 - 0x8e0  :  255 - 0xff -- Sprite 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11111111", -- 2274 - 0x8e2  :  255 - 0xff
    "11111111", -- 2275 - 0x8e3  :  255 - 0xff
    "11111111", -- 2276 - 0x8e4  :  255 - 0xff
    "11111111", -- 2277 - 0x8e5  :  255 - 0xff
    "11111111", -- 2278 - 0x8e6  :  255 - 0xff
    "11111111", -- 2279 - 0x8e7  :  255 - 0xff
    "11111111", -- 2280 - 0x8e8  :  255 - 0xff
    "11111111", -- 2281 - 0x8e9  :  255 - 0xff
    "11111111", -- 2282 - 0x8ea  :  255 - 0xff
    "11111111", -- 2283 - 0x8eb  :  255 - 0xff
    "11111111", -- 2284 - 0x8ec  :  255 - 0xff
    "11111111", -- 2285 - 0x8ed  :  255 - 0xff
    "11111111", -- 2286 - 0x8ee  :  255 - 0xff
    "11111111", -- 2287 - 0x8ef  :  255 - 0xff
    "11111111", -- 2288 - 0x8f0  :  255 - 0xff -- Sprite 0x8f
    "11111111", -- 2289 - 0x8f1  :  255 - 0xff
    "11111111", -- 2290 - 0x8f2  :  255 - 0xff
    "11111111", -- 2291 - 0x8f3  :  255 - 0xff
    "11111111", -- 2292 - 0x8f4  :  255 - 0xff
    "11111111", -- 2293 - 0x8f5  :  255 - 0xff
    "11111111", -- 2294 - 0x8f6  :  255 - 0xff
    "11111111", -- 2295 - 0x8f7  :  255 - 0xff
    "11111111", -- 2296 - 0x8f8  :  255 - 0xff
    "11111111", -- 2297 - 0x8f9  :  255 - 0xff
    "11111111", -- 2298 - 0x8fa  :  255 - 0xff
    "11111111", -- 2299 - 0x8fb  :  255 - 0xff
    "11111111", -- 2300 - 0x8fc  :  255 - 0xff
    "11111111", -- 2301 - 0x8fd  :  255 - 0xff
    "11111111", -- 2302 - 0x8fe  :  255 - 0xff
    "11111111", -- 2303 - 0x8ff  :  255 - 0xff
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000000", -- 2308 - 0x904  :    0 - 0x0
    "00000001", -- 2309 - 0x905  :    1 - 0x1
    "00011110", -- 2310 - 0x906  :   30 - 0x1e
    "00111011", -- 2311 - 0x907  :   59 - 0x3b
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00000000", -- 2316 - 0x90c  :    0 - 0x0
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "00000000", -- 2318 - 0x90e  :    0 - 0x0
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "00000000", -- 2320 - 0x910  :    0 - 0x0 -- Sprite 0x91
    "00000000", -- 2321 - 0x911  :    0 - 0x0
    "00001100", -- 2322 - 0x912  :   12 - 0xc
    "00111100", -- 2323 - 0x913  :   60 - 0x3c
    "11010000", -- 2324 - 0x914  :  208 - 0xd0
    "00010000", -- 2325 - 0x915  :   16 - 0x10
    "00100000", -- 2326 - 0x916  :   32 - 0x20
    "01000000", -- 2327 - 0x917  :   64 - 0x40
    "00000000", -- 2328 - 0x918  :    0 - 0x0
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00000000", -- 2331 - 0x91b  :    0 - 0x0
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00111110", -- 2336 - 0x920  :   62 - 0x3e -- Sprite 0x92
    "00101101", -- 2337 - 0x921  :   45 - 0x2d
    "00110101", -- 2338 - 0x922  :   53 - 0x35
    "00011101", -- 2339 - 0x923  :   29 - 0x1d
    "00000001", -- 2340 - 0x924  :    1 - 0x1
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00000000", -- 2344 - 0x928  :    0 - 0x0
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "00000000", -- 2349 - 0x92d  :    0 - 0x0
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "10110000", -- 2352 - 0x930  :  176 - 0xb0 -- Sprite 0x93
    "10111000", -- 2353 - 0x931  :  184 - 0xb8
    "11111000", -- 2354 - 0x932  :  248 - 0xf8
    "01111000", -- 2355 - 0x933  :  120 - 0x78
    "10011000", -- 2356 - 0x934  :  152 - 0x98
    "11110000", -- 2357 - 0x935  :  240 - 0xf0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "00000000", -- 2362 - 0x93a  :    0 - 0x0
    "00000000", -- 2363 - 0x93b  :    0 - 0x0
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000111", -- 2370 - 0x942  :    7 - 0x7
    "00000011", -- 2371 - 0x943  :    3 - 0x3
    "00001101", -- 2372 - 0x944  :   13 - 0xd
    "00011110", -- 2373 - 0x945  :   30 - 0x1e
    "00010111", -- 2374 - 0x946  :   23 - 0x17
    "00011101", -- 2375 - 0x947  :   29 - 0x1d
    "00000000", -- 2376 - 0x948  :    0 - 0x0
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00000000", -- 2380 - 0x94c  :    0 - 0x0
    "00000000", -- 2381 - 0x94d  :    0 - 0x0
    "00000000", -- 2382 - 0x94e  :    0 - 0x0
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00000000", -- 2384 - 0x950  :    0 - 0x0 -- Sprite 0x95
    "10000000", -- 2385 - 0x951  :  128 - 0x80
    "01110000", -- 2386 - 0x952  :  112 - 0x70
    "11100000", -- 2387 - 0x953  :  224 - 0xe0
    "11011000", -- 2388 - 0x954  :  216 - 0xd8
    "10111100", -- 2389 - 0x955  :  188 - 0xbc
    "01110100", -- 2390 - 0x956  :  116 - 0x74
    "11011100", -- 2391 - 0x957  :  220 - 0xdc
    "00000000", -- 2392 - 0x958  :    0 - 0x0
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00011111", -- 2400 - 0x960  :   31 - 0x1f -- Sprite 0x96
    "00001011", -- 2401 - 0x961  :   11 - 0xb
    "00001111", -- 2402 - 0x962  :   15 - 0xf
    "00000101", -- 2403 - 0x963  :    5 - 0x5
    "00000011", -- 2404 - 0x964  :    3 - 0x3
    "00000001", -- 2405 - 0x965  :    1 - 0x1
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "00000000", -- 2410 - 0x96a  :    0 - 0x0
    "00000000", -- 2411 - 0x96b  :    0 - 0x0
    "00000000", -- 2412 - 0x96c  :    0 - 0x0
    "00000000", -- 2413 - 0x96d  :    0 - 0x0
    "00000000", -- 2414 - 0x96e  :    0 - 0x0
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "11111100", -- 2416 - 0x970  :  252 - 0xfc -- Sprite 0x97
    "01101000", -- 2417 - 0x971  :  104 - 0x68
    "11111000", -- 2418 - 0x972  :  248 - 0xf8
    "10110000", -- 2419 - 0x973  :  176 - 0xb0
    "11100000", -- 2420 - 0x974  :  224 - 0xe0
    "10000000", -- 2421 - 0x975  :  128 - 0x80
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000000", -- 2424 - 0x978  :    0 - 0x0
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "00000000", -- 2426 - 0x97a  :    0 - 0x0
    "00000000", -- 2427 - 0x97b  :    0 - 0x0
    "00000000", -- 2428 - 0x97c  :    0 - 0x0
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Sprite 0x98
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000001", -- 2435 - 0x983  :    1 - 0x1
    "00000001", -- 2436 - 0x984  :    1 - 0x1
    "00001011", -- 2437 - 0x985  :   11 - 0xb
    "00011100", -- 2438 - 0x986  :   28 - 0x1c
    "00111111", -- 2439 - 0x987  :   63 - 0x3f
    "00000000", -- 2440 - 0x988  :    0 - 0x0
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Sprite 0x99
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00110000", -- 2450 - 0x992  :   48 - 0x30
    "01111000", -- 2451 - 0x993  :  120 - 0x78
    "10000000", -- 2452 - 0x994  :  128 - 0x80
    "11110000", -- 2453 - 0x995  :  240 - 0xf0
    "11111000", -- 2454 - 0x996  :  248 - 0xf8
    "11111100", -- 2455 - 0x997  :  252 - 0xfc
    "00000000", -- 2456 - 0x998  :    0 - 0x0
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00111111", -- 2464 - 0x9a0  :   63 - 0x3f -- Sprite 0x9a
    "00111111", -- 2465 - 0x9a1  :   63 - 0x3f
    "00111111", -- 2466 - 0x9a2  :   63 - 0x3f
    "00011111", -- 2467 - 0x9a3  :   31 - 0x1f
    "00011111", -- 2468 - 0x9a4  :   31 - 0x1f
    "00000111", -- 2469 - 0x9a5  :    7 - 0x7
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "11111100", -- 2480 - 0x9b0  :  252 - 0xfc -- Sprite 0x9b
    "11101100", -- 2481 - 0x9b1  :  236 - 0xec
    "11101100", -- 2482 - 0x9b2  :  236 - 0xec
    "11011000", -- 2483 - 0x9b3  :  216 - 0xd8
    "11111000", -- 2484 - 0x9b4  :  248 - 0xf8
    "11100000", -- 2485 - 0x9b5  :  224 - 0xe0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Sprite 0x9c
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000001", -- 2498 - 0x9c2  :    1 - 0x1
    "00011101", -- 2499 - 0x9c3  :   29 - 0x1d
    "00111110", -- 2500 - 0x9c4  :   62 - 0x3e
    "00111111", -- 2501 - 0x9c5  :   63 - 0x3f
    "00111111", -- 2502 - 0x9c6  :   63 - 0x3f
    "00111111", -- 2503 - 0x9c7  :   63 - 0x3f
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Sprite 0x9d
    "10000000", -- 2513 - 0x9d1  :  128 - 0x80
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "01110000", -- 2515 - 0x9d3  :  112 - 0x70
    "11111000", -- 2516 - 0x9d4  :  248 - 0xf8
    "11111100", -- 2517 - 0x9d5  :  252 - 0xfc
    "11111100", -- 2518 - 0x9d6  :  252 - 0xfc
    "11111100", -- 2519 - 0x9d7  :  252 - 0xfc
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00111111", -- 2528 - 0x9e0  :   63 - 0x3f -- Sprite 0x9e
    "00111111", -- 2529 - 0x9e1  :   63 - 0x3f
    "00011111", -- 2530 - 0x9e2  :   31 - 0x1f
    "00011111", -- 2531 - 0x9e3  :   31 - 0x1f
    "00001111", -- 2532 - 0x9e4  :   15 - 0xf
    "00000110", -- 2533 - 0x9e5  :    6 - 0x6
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "11101100", -- 2544 - 0x9f0  :  236 - 0xec -- Sprite 0x9f
    "11101100", -- 2545 - 0x9f1  :  236 - 0xec
    "11011000", -- 2546 - 0x9f2  :  216 - 0xd8
    "11111000", -- 2547 - 0x9f3  :  248 - 0xf8
    "11110000", -- 2548 - 0x9f4  :  240 - 0xf0
    "11100000", -- 2549 - 0x9f5  :  224 - 0xe0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Sprite 0xa0
    "00000100", -- 2561 - 0xa01  :    4 - 0x4
    "00000011", -- 2562 - 0xa02  :    3 - 0x3
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000001", -- 2564 - 0xa04  :    1 - 0x1
    "00000111", -- 2565 - 0xa05  :    7 - 0x7
    "00001111", -- 2566 - 0xa06  :   15 - 0xf
    "00001100", -- 2567 - 0xa07  :   12 - 0xc
    "00000000", -- 2568 - 0xa08  :    0 - 0x0
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Sprite 0xa1
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "11100000", -- 2578 - 0xa12  :  224 - 0xe0
    "10000000", -- 2579 - 0xa13  :  128 - 0x80
    "01000000", -- 2580 - 0xa14  :   64 - 0x40
    "11110000", -- 2581 - 0xa15  :  240 - 0xf0
    "10011000", -- 2582 - 0xa16  :  152 - 0x98
    "11111000", -- 2583 - 0xa17  :  248 - 0xf8
    "00000000", -- 2584 - 0xa18  :    0 - 0x0
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00011111", -- 2592 - 0xa20  :   31 - 0x1f -- Sprite 0xa2
    "00010011", -- 2593 - 0xa21  :   19 - 0x13
    "00011111", -- 2594 - 0xa22  :   31 - 0x1f
    "00001111", -- 2595 - 0xa23  :   15 - 0xf
    "00001001", -- 2596 - 0xa24  :    9 - 0x9
    "00000111", -- 2597 - 0xa25  :    7 - 0x7
    "00000001", -- 2598 - 0xa26  :    1 - 0x1
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "11100100", -- 2608 - 0xa30  :  228 - 0xe4 -- Sprite 0xa3
    "00111100", -- 2609 - 0xa31  :   60 - 0x3c
    "11100100", -- 2610 - 0xa32  :  228 - 0xe4
    "00111000", -- 2611 - 0xa33  :   56 - 0x38
    "11111000", -- 2612 - 0xa34  :  248 - 0xf8
    "11110000", -- 2613 - 0xa35  :  240 - 0xf0
    "11000000", -- 2614 - 0xa36  :  192 - 0xc0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Sprite 0xa4
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00010001", -- 2628 - 0xa44  :   17 - 0x11
    "00010011", -- 2629 - 0xa45  :   19 - 0x13
    "00011111", -- 2630 - 0xa46  :   31 - 0x1f
    "00011111", -- 2631 - 0xa47  :   31 - 0x1f
    "00000000", -- 2632 - 0xa48  :    0 - 0x0
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "10000000", -- 2643 - 0xa53  :  128 - 0x80
    "11000100", -- 2644 - 0xa54  :  196 - 0xc4
    "11100100", -- 2645 - 0xa55  :  228 - 0xe4
    "11111100", -- 2646 - 0xa56  :  252 - 0xfc
    "11111100", -- 2647 - 0xa57  :  252 - 0xfc
    "00000000", -- 2648 - 0xa58  :    0 - 0x0
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00011111", -- 2656 - 0xa60  :   31 - 0x1f -- Sprite 0xa6
    "00001110", -- 2657 - 0xa61  :   14 - 0xe
    "00000110", -- 2658 - 0xa62  :    6 - 0x6
    "00000010", -- 2659 - 0xa63  :    2 - 0x2
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "11111100", -- 2672 - 0xa70  :  252 - 0xfc -- Sprite 0xa7
    "10111000", -- 2673 - 0xa71  :  184 - 0xb8
    "10110000", -- 2674 - 0xa72  :  176 - 0xb0
    "10100000", -- 2675 - 0xa73  :  160 - 0xa0
    "10000000", -- 2676 - 0xa74  :  128 - 0x80
    "00000000", -- 2677 - 0xa75  :    0 - 0x0
    "00000000", -- 2678 - 0xa76  :    0 - 0x0
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00000000", -- 2680 - 0xa78  :    0 - 0x0
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000000", -- 2685 - 0xa7d  :    0 - 0x0
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000001", -- 2691 - 0xa83  :    1 - 0x1
    "00000011", -- 2692 - 0xa84  :    3 - 0x3
    "00000110", -- 2693 - 0xa85  :    6 - 0x6
    "00000110", -- 2694 - 0xa86  :    6 - 0x6
    "00001111", -- 2695 - 0xa87  :   15 - 0xf
    "00000000", -- 2696 - 0xa88  :    0 - 0x0
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000000", -- 2703 - 0xa8f  :    0 - 0x0
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Sprite 0xa9
    "00011000", -- 2705 - 0xa91  :   24 - 0x18
    "11110100", -- 2706 - 0xa92  :  244 - 0xf4
    "11111000", -- 2707 - 0xa93  :  248 - 0xf8
    "00111000", -- 2708 - 0xa94  :   56 - 0x38
    "01111100", -- 2709 - 0xa95  :  124 - 0x7c
    "11111100", -- 2710 - 0xa96  :  252 - 0xfc
    "11111100", -- 2711 - 0xa97  :  252 - 0xfc
    "00000000", -- 2712 - 0xa98  :    0 - 0x0
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00001111", -- 2720 - 0xaa0  :   15 - 0xf -- Sprite 0xaa
    "00011111", -- 2721 - 0xaa1  :   31 - 0x1f
    "00110000", -- 2722 - 0xaa2  :   48 - 0x30
    "00111000", -- 2723 - 0xaa3  :   56 - 0x38
    "00011101", -- 2724 - 0xaa4  :   29 - 0x1d
    "00000011", -- 2725 - 0xaa5  :    3 - 0x3
    "00000011", -- 2726 - 0xaa6  :    3 - 0x3
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "00000000", -- 2733 - 0xaad  :    0 - 0x0
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "11111100", -- 2736 - 0xab0  :  252 - 0xfc -- Sprite 0xab
    "11111100", -- 2737 - 0xab1  :  252 - 0xfc
    "01111100", -- 2738 - 0xab2  :  124 - 0x7c
    "10001110", -- 2739 - 0xab3  :  142 - 0x8e
    "10000110", -- 2740 - 0xab4  :  134 - 0x86
    "10011100", -- 2741 - 0xab5  :  156 - 0x9c
    "01111000", -- 2742 - 0xab6  :  120 - 0x78
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000001", -- 2753 - 0xac1  :    1 - 0x1
    "00000110", -- 2754 - 0xac2  :    6 - 0x6
    "00000111", -- 2755 - 0xac3  :    7 - 0x7
    "00000111", -- 2756 - 0xac4  :    7 - 0x7
    "00000111", -- 2757 - 0xac5  :    7 - 0x7
    "00000001", -- 2758 - 0xac6  :    1 - 0x1
    "00000011", -- 2759 - 0xac7  :    3 - 0x3
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Sprite 0xad
    "11000000", -- 2769 - 0xad1  :  192 - 0xc0
    "00110000", -- 2770 - 0xad2  :   48 - 0x30
    "11110000", -- 2771 - 0xad3  :  240 - 0xf0
    "11110000", -- 2772 - 0xad4  :  240 - 0xf0
    "11110000", -- 2773 - 0xad5  :  240 - 0xf0
    "01000000", -- 2774 - 0xad6  :   64 - 0x40
    "01000000", -- 2775 - 0xad7  :   64 - 0x40
    "00000000", -- 2776 - 0xad8  :    0 - 0x0
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000001", -- 2784 - 0xae0  :    1 - 0x1 -- Sprite 0xae
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000001", -- 2786 - 0xae2  :    1 - 0x1
    "00000011", -- 2787 - 0xae3  :    3 - 0x3
    "00000001", -- 2788 - 0xae4  :    1 - 0x1
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "01000000", -- 2800 - 0xaf0  :   64 - 0x40 -- Sprite 0xaf
    "01000000", -- 2801 - 0xaf1  :   64 - 0x40
    "01000000", -- 2802 - 0xaf2  :   64 - 0x40
    "01000000", -- 2803 - 0xaf3  :   64 - 0x40
    "01000000", -- 2804 - 0xaf4  :   64 - 0x40
    "10000000", -- 2805 - 0xaf5  :  128 - 0x80
    "00000000", -- 2806 - 0xaf6  :    0 - 0x0
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "01111110", -- 2816 - 0xb00  :  126 - 0x7e -- Sprite 0xb0
    "01100011", -- 2817 - 0xb01  :   99 - 0x63
    "01100011", -- 2818 - 0xb02  :   99 - 0x63
    "01100011", -- 2819 - 0xb03  :   99 - 0x63
    "01111110", -- 2820 - 0xb04  :  126 - 0x7e
    "01100000", -- 2821 - 0xb05  :   96 - 0x60
    "01100000", -- 2822 - 0xb06  :   96 - 0x60
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "01111110", -- 2824 - 0xb08  :  126 - 0x7e
    "01100011", -- 2825 - 0xb09  :   99 - 0x63
    "01100011", -- 2826 - 0xb0a  :   99 - 0x63
    "01100011", -- 2827 - 0xb0b  :   99 - 0x63
    "01111110", -- 2828 - 0xb0c  :  126 - 0x7e
    "01100000", -- 2829 - 0xb0d  :   96 - 0x60
    "01100000", -- 2830 - 0xb0e  :   96 - 0x60
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "01100000", -- 2832 - 0xb10  :   96 - 0x60 -- Sprite 0xb1
    "01100000", -- 2833 - 0xb11  :   96 - 0x60
    "01100000", -- 2834 - 0xb12  :   96 - 0x60
    "01100000", -- 2835 - 0xb13  :   96 - 0x60
    "01100000", -- 2836 - 0xb14  :   96 - 0x60
    "01100000", -- 2837 - 0xb15  :   96 - 0x60
    "01111111", -- 2838 - 0xb16  :  127 - 0x7f
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "01100000", -- 2840 - 0xb18  :   96 - 0x60
    "01100000", -- 2841 - 0xb19  :   96 - 0x60
    "01100000", -- 2842 - 0xb1a  :   96 - 0x60
    "01100000", -- 2843 - 0xb1b  :   96 - 0x60
    "01100000", -- 2844 - 0xb1c  :   96 - 0x60
    "01100000", -- 2845 - 0xb1d  :   96 - 0x60
    "01111111", -- 2846 - 0xb1e  :  127 - 0x7f
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00011100", -- 2848 - 0xb20  :   28 - 0x1c -- Sprite 0xb2
    "00110110", -- 2849 - 0xb21  :   54 - 0x36
    "01100011", -- 2850 - 0xb22  :   99 - 0x63
    "01100011", -- 2851 - 0xb23  :   99 - 0x63
    "01111111", -- 2852 - 0xb24  :  127 - 0x7f
    "01100011", -- 2853 - 0xb25  :   99 - 0x63
    "01100011", -- 2854 - 0xb26  :   99 - 0x63
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00011100", -- 2856 - 0xb28  :   28 - 0x1c
    "00110110", -- 2857 - 0xb29  :   54 - 0x36
    "01100011", -- 2858 - 0xb2a  :   99 - 0x63
    "01100011", -- 2859 - 0xb2b  :   99 - 0x63
    "01111111", -- 2860 - 0xb2c  :  127 - 0x7f
    "01100011", -- 2861 - 0xb2d  :   99 - 0x63
    "01100011", -- 2862 - 0xb2e  :   99 - 0x63
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00110011", -- 2864 - 0xb30  :   51 - 0x33 -- Sprite 0xb3
    "00110011", -- 2865 - 0xb31  :   51 - 0x33
    "00110011", -- 2866 - 0xb32  :   51 - 0x33
    "00011110", -- 2867 - 0xb33  :   30 - 0x1e
    "00001100", -- 2868 - 0xb34  :   12 - 0xc
    "00001100", -- 2869 - 0xb35  :   12 - 0xc
    "00001100", -- 2870 - 0xb36  :   12 - 0xc
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "00110011", -- 2872 - 0xb38  :   51 - 0x33
    "00110011", -- 2873 - 0xb39  :   51 - 0x33
    "00110011", -- 2874 - 0xb3a  :   51 - 0x33
    "00011110", -- 2875 - 0xb3b  :   30 - 0x1e
    "00001100", -- 2876 - 0xb3c  :   12 - 0xc
    "00001100", -- 2877 - 0xb3d  :   12 - 0xc
    "00001100", -- 2878 - 0xb3e  :   12 - 0xc
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "01111111", -- 2880 - 0xb40  :  127 - 0x7f -- Sprite 0xb4
    "01100000", -- 2881 - 0xb41  :   96 - 0x60
    "01100000", -- 2882 - 0xb42  :   96 - 0x60
    "01111110", -- 2883 - 0xb43  :  126 - 0x7e
    "01100000", -- 2884 - 0xb44  :   96 - 0x60
    "01100000", -- 2885 - 0xb45  :   96 - 0x60
    "01111111", -- 2886 - 0xb46  :  127 - 0x7f
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "01111111", -- 2888 - 0xb48  :  127 - 0x7f
    "01100000", -- 2889 - 0xb49  :   96 - 0x60
    "01100000", -- 2890 - 0xb4a  :   96 - 0x60
    "01111110", -- 2891 - 0xb4b  :  126 - 0x7e
    "01100000", -- 2892 - 0xb4c  :   96 - 0x60
    "01100000", -- 2893 - 0xb4d  :   96 - 0x60
    "01111111", -- 2894 - 0xb4e  :  127 - 0x7f
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "01111110", -- 2896 - 0xb50  :  126 - 0x7e -- Sprite 0xb5
    "01100011", -- 2897 - 0xb51  :   99 - 0x63
    "01100011", -- 2898 - 0xb52  :   99 - 0x63
    "01100111", -- 2899 - 0xb53  :  103 - 0x67
    "01111100", -- 2900 - 0xb54  :  124 - 0x7c
    "01101110", -- 2901 - 0xb55  :  110 - 0x6e
    "01100111", -- 2902 - 0xb56  :  103 - 0x67
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "01111110", -- 2904 - 0xb58  :  126 - 0x7e
    "01100011", -- 2905 - 0xb59  :   99 - 0x63
    "01100011", -- 2906 - 0xb5a  :   99 - 0x63
    "01100111", -- 2907 - 0xb5b  :  103 - 0x67
    "01111100", -- 2908 - 0xb5c  :  124 - 0x7c
    "01101110", -- 2909 - 0xb5d  :  110 - 0x6e
    "01100111", -- 2910 - 0xb5e  :  103 - 0x67
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00111110", -- 2912 - 0xb60  :   62 - 0x3e -- Sprite 0xb6
    "01100011", -- 2913 - 0xb61  :   99 - 0x63
    "01100011", -- 2914 - 0xb62  :   99 - 0x63
    "01100011", -- 2915 - 0xb63  :   99 - 0x63
    "01100011", -- 2916 - 0xb64  :   99 - 0x63
    "01100011", -- 2917 - 0xb65  :   99 - 0x63
    "00111110", -- 2918 - 0xb66  :   62 - 0x3e
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00111110", -- 2920 - 0xb68  :   62 - 0x3e
    "01100011", -- 2921 - 0xb69  :   99 - 0x63
    "01100011", -- 2922 - 0xb6a  :   99 - 0x63
    "01100011", -- 2923 - 0xb6b  :   99 - 0x63
    "01100011", -- 2924 - 0xb6c  :   99 - 0x63
    "01100011", -- 2925 - 0xb6d  :   99 - 0x63
    "00111110", -- 2926 - 0xb6e  :   62 - 0x3e
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "01100011", -- 2928 - 0xb70  :   99 - 0x63 -- Sprite 0xb7
    "01110011", -- 2929 - 0xb71  :  115 - 0x73
    "01111011", -- 2930 - 0xb72  :  123 - 0x7b
    "01111111", -- 2931 - 0xb73  :  127 - 0x7f
    "01101111", -- 2932 - 0xb74  :  111 - 0x6f
    "01100111", -- 2933 - 0xb75  :  103 - 0x67
    "01100011", -- 2934 - 0xb76  :   99 - 0x63
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "01100011", -- 2936 - 0xb78  :   99 - 0x63
    "01110011", -- 2937 - 0xb79  :  115 - 0x73
    "01111011", -- 2938 - 0xb7a  :  123 - 0x7b
    "01111111", -- 2939 - 0xb7b  :  127 - 0x7f
    "01101111", -- 2940 - 0xb7c  :  111 - 0x6f
    "01100111", -- 2941 - 0xb7d  :  103 - 0x67
    "01100011", -- 2942 - 0xb7e  :   99 - 0x63
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00111111", -- 2944 - 0xb80  :   63 - 0x3f -- Sprite 0xb8
    "00001100", -- 2945 - 0xb81  :   12 - 0xc
    "00001100", -- 2946 - 0xb82  :   12 - 0xc
    "00001100", -- 2947 - 0xb83  :   12 - 0xc
    "00001100", -- 2948 - 0xb84  :   12 - 0xc
    "00001100", -- 2949 - 0xb85  :   12 - 0xc
    "00001100", -- 2950 - 0xb86  :   12 - 0xc
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00111111", -- 2952 - 0xb88  :   63 - 0x3f
    "00001100", -- 2953 - 0xb89  :   12 - 0xc
    "00001100", -- 2954 - 0xb8a  :   12 - 0xc
    "00001100", -- 2955 - 0xb8b  :   12 - 0xc
    "00001100", -- 2956 - 0xb8c  :   12 - 0xc
    "00001100", -- 2957 - 0xb8d  :   12 - 0xc
    "00001100", -- 2958 - 0xb8e  :   12 - 0xc
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "01100011", -- 2960 - 0xb90  :   99 - 0x63 -- Sprite 0xb9
    "01100011", -- 2961 - 0xb91  :   99 - 0x63
    "01101011", -- 2962 - 0xb92  :  107 - 0x6b
    "01111111", -- 2963 - 0xb93  :  127 - 0x7f
    "01111111", -- 2964 - 0xb94  :  127 - 0x7f
    "01110111", -- 2965 - 0xb95  :  119 - 0x77
    "01100011", -- 2966 - 0xb96  :   99 - 0x63
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "01100011", -- 2968 - 0xb98  :   99 - 0x63
    "01100011", -- 2969 - 0xb99  :   99 - 0x63
    "01101011", -- 2970 - 0xb9a  :  107 - 0x6b
    "01111111", -- 2971 - 0xb9b  :  127 - 0x7f
    "01111111", -- 2972 - 0xb9c  :  127 - 0x7f
    "01110111", -- 2973 - 0xb9d  :  119 - 0x77
    "01100011", -- 2974 - 0xb9e  :   99 - 0x63
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "01111100", -- 2976 - 0xba0  :  124 - 0x7c -- Sprite 0xba
    "01100110", -- 2977 - 0xba1  :  102 - 0x66
    "01100011", -- 2978 - 0xba2  :   99 - 0x63
    "01100011", -- 2979 - 0xba3  :   99 - 0x63
    "01100011", -- 2980 - 0xba4  :   99 - 0x63
    "01100110", -- 2981 - 0xba5  :  102 - 0x66
    "01111100", -- 2982 - 0xba6  :  124 - 0x7c
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "00000000", -- 2984 - 0xba8  :    0 - 0x0
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00011100", -- 2992 - 0xbb0  :   28 - 0x1c -- Sprite 0xbb
    "00011100", -- 2993 - 0xbb1  :   28 - 0x1c
    "00011100", -- 2994 - 0xbb2  :   28 - 0x1c
    "00011000", -- 2995 - 0xbb3  :   24 - 0x18
    "00011000", -- 2996 - 0xbb4  :   24 - 0x18
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00011000", -- 2998 - 0xbb6  :   24 - 0x18
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00011111", -- 3008 - 0xbc0  :   31 - 0x1f -- Sprite 0xbc
    "00110000", -- 3009 - 0xbc1  :   48 - 0x30
    "01100000", -- 3010 - 0xbc2  :   96 - 0x60
    "01100111", -- 3011 - 0xbc3  :  103 - 0x67
    "01100011", -- 3012 - 0xbc4  :   99 - 0x63
    "00110011", -- 3013 - 0xbc5  :   51 - 0x33
    "00011111", -- 3014 - 0xbc6  :   31 - 0x1f
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00011111", -- 3016 - 0xbc8  :   31 - 0x1f
    "00110000", -- 3017 - 0xbc9  :   48 - 0x30
    "01100000", -- 3018 - 0xbca  :   96 - 0x60
    "01100111", -- 3019 - 0xbcb  :  103 - 0x67
    "01100011", -- 3020 - 0xbcc  :   99 - 0x63
    "00110011", -- 3021 - 0xbcd  :   51 - 0x33
    "00011111", -- 3022 - 0xbce  :   31 - 0x1f
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "01100011", -- 3024 - 0xbd0  :   99 - 0x63 -- Sprite 0xbd
    "01110111", -- 3025 - 0xbd1  :  119 - 0x77
    "01111111", -- 3026 - 0xbd2  :  127 - 0x7f
    "01111111", -- 3027 - 0xbd3  :  127 - 0x7f
    "01101011", -- 3028 - 0xbd4  :  107 - 0x6b
    "01100011", -- 3029 - 0xbd5  :   99 - 0x63
    "01100011", -- 3030 - 0xbd6  :   99 - 0x63
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "01100011", -- 3032 - 0xbd8  :   99 - 0x63
    "01110111", -- 3033 - 0xbd9  :  119 - 0x77
    "01111111", -- 3034 - 0xbda  :  127 - 0x7f
    "01111111", -- 3035 - 0xbdb  :  127 - 0x7f
    "01101011", -- 3036 - 0xbdc  :  107 - 0x6b
    "01100011", -- 3037 - 0xbdd  :   99 - 0x63
    "01100011", -- 3038 - 0xbde  :   99 - 0x63
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "01100011", -- 3040 - 0xbe0  :   99 - 0x63 -- Sprite 0xbe
    "01100011", -- 3041 - 0xbe1  :   99 - 0x63
    "01100011", -- 3042 - 0xbe2  :   99 - 0x63
    "01110111", -- 3043 - 0xbe3  :  119 - 0x77
    "00111110", -- 3044 - 0xbe4  :   62 - 0x3e
    "00011100", -- 3045 - 0xbe5  :   28 - 0x1c
    "00001000", -- 3046 - 0xbe6  :    8 - 0x8
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "01100011", -- 3048 - 0xbe8  :   99 - 0x63
    "01100011", -- 3049 - 0xbe9  :   99 - 0x63
    "01100011", -- 3050 - 0xbea  :   99 - 0x63
    "01110111", -- 3051 - 0xbeb  :  119 - 0x77
    "00111110", -- 3052 - 0xbec  :   62 - 0x3e
    "00011100", -- 3053 - 0xbed  :   28 - 0x1c
    "00001000", -- 3054 - 0xbee  :    8 - 0x8
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00011111", -- 3072 - 0xc00  :   31 - 0x1f -- Sprite 0xc0
    "00110000", -- 3073 - 0xc01  :   48 - 0x30
    "01100000", -- 3074 - 0xc02  :   96 - 0x60
    "01100111", -- 3075 - 0xc03  :  103 - 0x67
    "01100011", -- 3076 - 0xc04  :   99 - 0x63
    "00110011", -- 3077 - 0xc05  :   51 - 0x33
    "00011111", -- 3078 - 0xc06  :   31 - 0x1f
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00011100", -- 3088 - 0xc10  :   28 - 0x1c -- Sprite 0xc1
    "00110110", -- 3089 - 0xc11  :   54 - 0x36
    "01100011", -- 3090 - 0xc12  :   99 - 0x63
    "01100011", -- 3091 - 0xc13  :   99 - 0x63
    "01111111", -- 3092 - 0xc14  :  127 - 0x7f
    "01100011", -- 3093 - 0xc15  :   99 - 0x63
    "01100011", -- 3094 - 0xc16  :   99 - 0x63
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "01100011", -- 3104 - 0xc20  :   99 - 0x63 -- Sprite 0xc2
    "01110111", -- 3105 - 0xc21  :  119 - 0x77
    "01111111", -- 3106 - 0xc22  :  127 - 0x7f
    "01111111", -- 3107 - 0xc23  :  127 - 0x7f
    "01101011", -- 3108 - 0xc24  :  107 - 0x6b
    "01100011", -- 3109 - 0xc25  :   99 - 0x63
    "01100011", -- 3110 - 0xc26  :   99 - 0x63
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "01111111", -- 3120 - 0xc30  :  127 - 0x7f -- Sprite 0xc3
    "01100000", -- 3121 - 0xc31  :   96 - 0x60
    "01100000", -- 3122 - 0xc32  :   96 - 0x60
    "01111110", -- 3123 - 0xc33  :  126 - 0x7e
    "01100000", -- 3124 - 0xc34  :   96 - 0x60
    "01100000", -- 3125 - 0xc35  :   96 - 0x60
    "01111111", -- 3126 - 0xc36  :  127 - 0x7f
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00111110", -- 3136 - 0xc40  :   62 - 0x3e -- Sprite 0xc4
    "01100011", -- 3137 - 0xc41  :   99 - 0x63
    "01100011", -- 3138 - 0xc42  :   99 - 0x63
    "01100011", -- 3139 - 0xc43  :   99 - 0x63
    "01100011", -- 3140 - 0xc44  :   99 - 0x63
    "01100011", -- 3141 - 0xc45  :   99 - 0x63
    "00111110", -- 3142 - 0xc46  :   62 - 0x3e
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "01100011", -- 3152 - 0xc50  :   99 - 0x63 -- Sprite 0xc5
    "01100011", -- 3153 - 0xc51  :   99 - 0x63
    "01100011", -- 3154 - 0xc52  :   99 - 0x63
    "01110111", -- 3155 - 0xc53  :  119 - 0x77
    "00111110", -- 3156 - 0xc54  :   62 - 0x3e
    "00011100", -- 3157 - 0xc55  :   28 - 0x1c
    "00001000", -- 3158 - 0xc56  :    8 - 0x8
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "00000000", -- 3160 - 0xc58  :    0 - 0x0
    "00000000", -- 3161 - 0xc59  :    0 - 0x0
    "00000000", -- 3162 - 0xc5a  :    0 - 0x0
    "00000000", -- 3163 - 0xc5b  :    0 - 0x0
    "00000000", -- 3164 - 0xc5c  :    0 - 0x0
    "00000000", -- 3165 - 0xc5d  :    0 - 0x0
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "01111110", -- 3168 - 0xc60  :  126 - 0x7e -- Sprite 0xc6
    "01100011", -- 3169 - 0xc61  :   99 - 0x63
    "01100011", -- 3170 - 0xc62  :   99 - 0x63
    "01100111", -- 3171 - 0xc63  :  103 - 0x67
    "01111100", -- 3172 - 0xc64  :  124 - 0x7c
    "01101110", -- 3173 - 0xc65  :  110 - 0x6e
    "01100111", -- 3174 - 0xc66  :  103 - 0x67
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "00000000", -- 3181 - 0xc6d  :    0 - 0x0
    "00000000", -- 3182 - 0xc6e  :    0 - 0x0
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00110011", -- 3184 - 0xc70  :   51 - 0x33 -- Sprite 0xc7
    "00110011", -- 3185 - 0xc71  :   51 - 0x33
    "00110011", -- 3186 - 0xc72  :   51 - 0x33
    "00011110", -- 3187 - 0xc73  :   30 - 0x1e
    "00001100", -- 3188 - 0xc74  :   12 - 0xc
    "00001100", -- 3189 - 0xc75  :   12 - 0xc
    "00001100", -- 3190 - 0xc76  :   12 - 0xc
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "00000000", -- 3192 - 0xc78  :    0 - 0x0
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000000", -- 3196 - 0xc7c  :    0 - 0x0
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00000000", -- 3208 - 0xc88  :    0 - 0x0
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0 -- Sprite 0xc9
    "00000000", -- 3217 - 0xc91  :    0 - 0x0
    "00000000", -- 3218 - 0xc92  :    0 - 0x0
    "00000000", -- 3219 - 0xc93  :    0 - 0x0
    "00000000", -- 3220 - 0xc94  :    0 - 0x0
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00000000", -- 3224 - 0xc98  :    0 - 0x0
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00000000", -- 3226 - 0xc9a  :    0 - 0x0
    "00000000", -- 3227 - 0xc9b  :    0 - 0x0
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00000000", -- 3235 - 0xca3  :    0 - 0x0
    "00000000", -- 3236 - 0xca4  :    0 - 0x0
    "00000000", -- 3237 - 0xca5  :    0 - 0x0
    "00000000", -- 3238 - 0xca6  :    0 - 0x0
    "00000000", -- 3239 - 0xca7  :    0 - 0x0
    "00000000", -- 3240 - 0xca8  :    0 - 0x0
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00000000", -- 3243 - 0xcab  :    0 - 0x0
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00000000", -- 3250 - 0xcb2  :    0 - 0x0
    "00000000", -- 3251 - 0xcb3  :    0 - 0x0
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0
    "00000000", -- 3257 - 0xcb9  :    0 - 0x0
    "00000000", -- 3258 - 0xcba  :    0 - 0x0
    "00000000", -- 3259 - 0xcbb  :    0 - 0x0
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00000000", -- 3261 - 0xcbd  :    0 - 0x0
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000000", -- 3302 - 0xce6  :    0 - 0x0
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000000", -- 3309 - 0xced  :    0 - 0x0
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "11111111", -- 3328 - 0xd00  :  255 - 0xff -- Sprite 0xd0
    "11111111", -- 3329 - 0xd01  :  255 - 0xff
    "11111111", -- 3330 - 0xd02  :  255 - 0xff
    "11111111", -- 3331 - 0xd03  :  255 - 0xff
    "11111111", -- 3332 - 0xd04  :  255 - 0xff
    "11111111", -- 3333 - 0xd05  :  255 - 0xff
    "11111111", -- 3334 - 0xd06  :  255 - 0xff
    "11111111", -- 3335 - 0xd07  :  255 - 0xff
    "11111111", -- 3336 - 0xd08  :  255 - 0xff
    "11111111", -- 3337 - 0xd09  :  255 - 0xff
    "11111111", -- 3338 - 0xd0a  :  255 - 0xff
    "11111111", -- 3339 - 0xd0b  :  255 - 0xff
    "11111111", -- 3340 - 0xd0c  :  255 - 0xff
    "11111111", -- 3341 - 0xd0d  :  255 - 0xff
    "11111111", -- 3342 - 0xd0e  :  255 - 0xff
    "11111111", -- 3343 - 0xd0f  :  255 - 0xff
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Sprite 0xd1
    "11111111", -- 3345 - 0xd11  :  255 - 0xff
    "11111111", -- 3346 - 0xd12  :  255 - 0xff
    "11111111", -- 3347 - 0xd13  :  255 - 0xff
    "11111111", -- 3348 - 0xd14  :  255 - 0xff
    "11111111", -- 3349 - 0xd15  :  255 - 0xff
    "11111111", -- 3350 - 0xd16  :  255 - 0xff
    "11111111", -- 3351 - 0xd17  :  255 - 0xff
    "11111111", -- 3352 - 0xd18  :  255 - 0xff
    "11111111", -- 3353 - 0xd19  :  255 - 0xff
    "11111111", -- 3354 - 0xd1a  :  255 - 0xff
    "11111111", -- 3355 - 0xd1b  :  255 - 0xff
    "11111111", -- 3356 - 0xd1c  :  255 - 0xff
    "11111111", -- 3357 - 0xd1d  :  255 - 0xff
    "11111111", -- 3358 - 0xd1e  :  255 - 0xff
    "11111111", -- 3359 - 0xd1f  :  255 - 0xff
    "11111111", -- 3360 - 0xd20  :  255 - 0xff -- Sprite 0xd2
    "11111111", -- 3361 - 0xd21  :  255 - 0xff
    "11111111", -- 3362 - 0xd22  :  255 - 0xff
    "11111111", -- 3363 - 0xd23  :  255 - 0xff
    "11111111", -- 3364 - 0xd24  :  255 - 0xff
    "11111111", -- 3365 - 0xd25  :  255 - 0xff
    "11111111", -- 3366 - 0xd26  :  255 - 0xff
    "11111111", -- 3367 - 0xd27  :  255 - 0xff
    "11111111", -- 3368 - 0xd28  :  255 - 0xff
    "11111111", -- 3369 - 0xd29  :  255 - 0xff
    "11111111", -- 3370 - 0xd2a  :  255 - 0xff
    "11111111", -- 3371 - 0xd2b  :  255 - 0xff
    "11111111", -- 3372 - 0xd2c  :  255 - 0xff
    "11111111", -- 3373 - 0xd2d  :  255 - 0xff
    "11111111", -- 3374 - 0xd2e  :  255 - 0xff
    "11111111", -- 3375 - 0xd2f  :  255 - 0xff
    "11111111", -- 3376 - 0xd30  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11111111", -- 3380 - 0xd34  :  255 - 0xff
    "11111111", -- 3381 - 0xd35  :  255 - 0xff
    "11111111", -- 3382 - 0xd36  :  255 - 0xff
    "11111111", -- 3383 - 0xd37  :  255 - 0xff
    "11111111", -- 3384 - 0xd38  :  255 - 0xff
    "11111111", -- 3385 - 0xd39  :  255 - 0xff
    "11111111", -- 3386 - 0xd3a  :  255 - 0xff
    "11111111", -- 3387 - 0xd3b  :  255 - 0xff
    "11111111", -- 3388 - 0xd3c  :  255 - 0xff
    "11111111", -- 3389 - 0xd3d  :  255 - 0xff
    "11111111", -- 3390 - 0xd3e  :  255 - 0xff
    "11111111", -- 3391 - 0xd3f  :  255 - 0xff
    "11111111", -- 3392 - 0xd40  :  255 - 0xff -- Sprite 0xd4
    "11111111", -- 3393 - 0xd41  :  255 - 0xff
    "11111111", -- 3394 - 0xd42  :  255 - 0xff
    "11111111", -- 3395 - 0xd43  :  255 - 0xff
    "11111111", -- 3396 - 0xd44  :  255 - 0xff
    "11111111", -- 3397 - 0xd45  :  255 - 0xff
    "11111111", -- 3398 - 0xd46  :  255 - 0xff
    "11111111", -- 3399 - 0xd47  :  255 - 0xff
    "11111111", -- 3400 - 0xd48  :  255 - 0xff
    "11111111", -- 3401 - 0xd49  :  255 - 0xff
    "11111111", -- 3402 - 0xd4a  :  255 - 0xff
    "11111111", -- 3403 - 0xd4b  :  255 - 0xff
    "11111111", -- 3404 - 0xd4c  :  255 - 0xff
    "11111111", -- 3405 - 0xd4d  :  255 - 0xff
    "11111111", -- 3406 - 0xd4e  :  255 - 0xff
    "11111111", -- 3407 - 0xd4f  :  255 - 0xff
    "11111111", -- 3408 - 0xd50  :  255 - 0xff -- Sprite 0xd5
    "11111111", -- 3409 - 0xd51  :  255 - 0xff
    "11111111", -- 3410 - 0xd52  :  255 - 0xff
    "11111111", -- 3411 - 0xd53  :  255 - 0xff
    "11111111", -- 3412 - 0xd54  :  255 - 0xff
    "11111111", -- 3413 - 0xd55  :  255 - 0xff
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "11111111", -- 3416 - 0xd58  :  255 - 0xff
    "11111111", -- 3417 - 0xd59  :  255 - 0xff
    "11111111", -- 3418 - 0xd5a  :  255 - 0xff
    "11111111", -- 3419 - 0xd5b  :  255 - 0xff
    "11111111", -- 3420 - 0xd5c  :  255 - 0xff
    "11111111", -- 3421 - 0xd5d  :  255 - 0xff
    "11111111", -- 3422 - 0xd5e  :  255 - 0xff
    "11111111", -- 3423 - 0xd5f  :  255 - 0xff
    "11111111", -- 3424 - 0xd60  :  255 - 0xff -- Sprite 0xd6
    "11111111", -- 3425 - 0xd61  :  255 - 0xff
    "11111111", -- 3426 - 0xd62  :  255 - 0xff
    "11111111", -- 3427 - 0xd63  :  255 - 0xff
    "11111111", -- 3428 - 0xd64  :  255 - 0xff
    "11111111", -- 3429 - 0xd65  :  255 - 0xff
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "11111111", -- 3432 - 0xd68  :  255 - 0xff
    "11111111", -- 3433 - 0xd69  :  255 - 0xff
    "11111111", -- 3434 - 0xd6a  :  255 - 0xff
    "11111111", -- 3435 - 0xd6b  :  255 - 0xff
    "11111111", -- 3436 - 0xd6c  :  255 - 0xff
    "11111111", -- 3437 - 0xd6d  :  255 - 0xff
    "11111111", -- 3438 - 0xd6e  :  255 - 0xff
    "11111111", -- 3439 - 0xd6f  :  255 - 0xff
    "11111111", -- 3440 - 0xd70  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "11111111", -- 3442 - 0xd72  :  255 - 0xff
    "11111111", -- 3443 - 0xd73  :  255 - 0xff
    "11111111", -- 3444 - 0xd74  :  255 - 0xff
    "11111111", -- 3445 - 0xd75  :  255 - 0xff
    "11111111", -- 3446 - 0xd76  :  255 - 0xff
    "11111111", -- 3447 - 0xd77  :  255 - 0xff
    "11111111", -- 3448 - 0xd78  :  255 - 0xff
    "11111111", -- 3449 - 0xd79  :  255 - 0xff
    "11111111", -- 3450 - 0xd7a  :  255 - 0xff
    "11111111", -- 3451 - 0xd7b  :  255 - 0xff
    "11111111", -- 3452 - 0xd7c  :  255 - 0xff
    "11111111", -- 3453 - 0xd7d  :  255 - 0xff
    "11111111", -- 3454 - 0xd7e  :  255 - 0xff
    "11111111", -- 3455 - 0xd7f  :  255 - 0xff
    "11111111", -- 3456 - 0xd80  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 3457 - 0xd81  :  255 - 0xff
    "11111111", -- 3458 - 0xd82  :  255 - 0xff
    "11111111", -- 3459 - 0xd83  :  255 - 0xff
    "11111111", -- 3460 - 0xd84  :  255 - 0xff
    "11111111", -- 3461 - 0xd85  :  255 - 0xff
    "11111111", -- 3462 - 0xd86  :  255 - 0xff
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11111111", -- 3464 - 0xd88  :  255 - 0xff
    "11111111", -- 3465 - 0xd89  :  255 - 0xff
    "11111111", -- 3466 - 0xd8a  :  255 - 0xff
    "11111111", -- 3467 - 0xd8b  :  255 - 0xff
    "11111111", -- 3468 - 0xd8c  :  255 - 0xff
    "11111111", -- 3469 - 0xd8d  :  255 - 0xff
    "11111111", -- 3470 - 0xd8e  :  255 - 0xff
    "11111111", -- 3471 - 0xd8f  :  255 - 0xff
    "11111111", -- 3472 - 0xd90  :  255 - 0xff -- Sprite 0xd9
    "11111111", -- 3473 - 0xd91  :  255 - 0xff
    "11111111", -- 3474 - 0xd92  :  255 - 0xff
    "11111111", -- 3475 - 0xd93  :  255 - 0xff
    "11111111", -- 3476 - 0xd94  :  255 - 0xff
    "11111111", -- 3477 - 0xd95  :  255 - 0xff
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111111", -- 3479 - 0xd97  :  255 - 0xff
    "11111111", -- 3480 - 0xd98  :  255 - 0xff
    "11111111", -- 3481 - 0xd99  :  255 - 0xff
    "11111111", -- 3482 - 0xd9a  :  255 - 0xff
    "11111111", -- 3483 - 0xd9b  :  255 - 0xff
    "11111111", -- 3484 - 0xd9c  :  255 - 0xff
    "11111111", -- 3485 - 0xd9d  :  255 - 0xff
    "11111111", -- 3486 - 0xd9e  :  255 - 0xff
    "11111111", -- 3487 - 0xd9f  :  255 - 0xff
    "11111111", -- 3488 - 0xda0  :  255 - 0xff -- Sprite 0xda
    "11111111", -- 3489 - 0xda1  :  255 - 0xff
    "11111111", -- 3490 - 0xda2  :  255 - 0xff
    "11111111", -- 3491 - 0xda3  :  255 - 0xff
    "11111111", -- 3492 - 0xda4  :  255 - 0xff
    "11111111", -- 3493 - 0xda5  :  255 - 0xff
    "11111111", -- 3494 - 0xda6  :  255 - 0xff
    "11111111", -- 3495 - 0xda7  :  255 - 0xff
    "11111111", -- 3496 - 0xda8  :  255 - 0xff
    "11111111", -- 3497 - 0xda9  :  255 - 0xff
    "11111111", -- 3498 - 0xdaa  :  255 - 0xff
    "11111111", -- 3499 - 0xdab  :  255 - 0xff
    "11111111", -- 3500 - 0xdac  :  255 - 0xff
    "11111111", -- 3501 - 0xdad  :  255 - 0xff
    "11111111", -- 3502 - 0xdae  :  255 - 0xff
    "11111111", -- 3503 - 0xdaf  :  255 - 0xff
    "11111111", -- 3504 - 0xdb0  :  255 - 0xff -- Sprite 0xdb
    "11111111", -- 3505 - 0xdb1  :  255 - 0xff
    "11111111", -- 3506 - 0xdb2  :  255 - 0xff
    "11111111", -- 3507 - 0xdb3  :  255 - 0xff
    "11111111", -- 3508 - 0xdb4  :  255 - 0xff
    "11111111", -- 3509 - 0xdb5  :  255 - 0xff
    "11111111", -- 3510 - 0xdb6  :  255 - 0xff
    "11111111", -- 3511 - 0xdb7  :  255 - 0xff
    "11111111", -- 3512 - 0xdb8  :  255 - 0xff
    "11111111", -- 3513 - 0xdb9  :  255 - 0xff
    "11111111", -- 3514 - 0xdba  :  255 - 0xff
    "11111111", -- 3515 - 0xdbb  :  255 - 0xff
    "11111111", -- 3516 - 0xdbc  :  255 - 0xff
    "11111111", -- 3517 - 0xdbd  :  255 - 0xff
    "11111111", -- 3518 - 0xdbe  :  255 - 0xff
    "11111111", -- 3519 - 0xdbf  :  255 - 0xff
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Sprite 0xdc
    "11111111", -- 3521 - 0xdc1  :  255 - 0xff
    "11111111", -- 3522 - 0xdc2  :  255 - 0xff
    "11111111", -- 3523 - 0xdc3  :  255 - 0xff
    "11111111", -- 3524 - 0xdc4  :  255 - 0xff
    "11111111", -- 3525 - 0xdc5  :  255 - 0xff
    "11111111", -- 3526 - 0xdc6  :  255 - 0xff
    "11111111", -- 3527 - 0xdc7  :  255 - 0xff
    "11111111", -- 3528 - 0xdc8  :  255 - 0xff
    "11111111", -- 3529 - 0xdc9  :  255 - 0xff
    "11111111", -- 3530 - 0xdca  :  255 - 0xff
    "11111111", -- 3531 - 0xdcb  :  255 - 0xff
    "11111111", -- 3532 - 0xdcc  :  255 - 0xff
    "11111111", -- 3533 - 0xdcd  :  255 - 0xff
    "11111111", -- 3534 - 0xdce  :  255 - 0xff
    "11111111", -- 3535 - 0xdcf  :  255 - 0xff
    "11111111", -- 3536 - 0xdd0  :  255 - 0xff -- Sprite 0xdd
    "11111111", -- 3537 - 0xdd1  :  255 - 0xff
    "11111111", -- 3538 - 0xdd2  :  255 - 0xff
    "11111111", -- 3539 - 0xdd3  :  255 - 0xff
    "11111111", -- 3540 - 0xdd4  :  255 - 0xff
    "11111111", -- 3541 - 0xdd5  :  255 - 0xff
    "11111111", -- 3542 - 0xdd6  :  255 - 0xff
    "11111111", -- 3543 - 0xdd7  :  255 - 0xff
    "11111111", -- 3544 - 0xdd8  :  255 - 0xff
    "11111111", -- 3545 - 0xdd9  :  255 - 0xff
    "11111111", -- 3546 - 0xdda  :  255 - 0xff
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "11111111", -- 3548 - 0xddc  :  255 - 0xff
    "11111111", -- 3549 - 0xddd  :  255 - 0xff
    "11111111", -- 3550 - 0xdde  :  255 - 0xff
    "11111111", -- 3551 - 0xddf  :  255 - 0xff
    "11111111", -- 3552 - 0xde0  :  255 - 0xff -- Sprite 0xde
    "11111111", -- 3553 - 0xde1  :  255 - 0xff
    "11111111", -- 3554 - 0xde2  :  255 - 0xff
    "11111111", -- 3555 - 0xde3  :  255 - 0xff
    "11111111", -- 3556 - 0xde4  :  255 - 0xff
    "11111111", -- 3557 - 0xde5  :  255 - 0xff
    "11111111", -- 3558 - 0xde6  :  255 - 0xff
    "11111111", -- 3559 - 0xde7  :  255 - 0xff
    "11111111", -- 3560 - 0xde8  :  255 - 0xff
    "11111111", -- 3561 - 0xde9  :  255 - 0xff
    "11111111", -- 3562 - 0xdea  :  255 - 0xff
    "11111111", -- 3563 - 0xdeb  :  255 - 0xff
    "11111111", -- 3564 - 0xdec  :  255 - 0xff
    "11111111", -- 3565 - 0xded  :  255 - 0xff
    "11111111", -- 3566 - 0xdee  :  255 - 0xff
    "11111111", -- 3567 - 0xdef  :  255 - 0xff
    "11111111", -- 3568 - 0xdf0  :  255 - 0xff -- Sprite 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "11111111", -- 3570 - 0xdf2  :  255 - 0xff
    "11111111", -- 3571 - 0xdf3  :  255 - 0xff
    "11111111", -- 3572 - 0xdf4  :  255 - 0xff
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111111", -- 3575 - 0xdf7  :  255 - 0xff
    "11111111", -- 3576 - 0xdf8  :  255 - 0xff
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11111111", -- 3580 - 0xdfc  :  255 - 0xff
    "11111111", -- 3581 - 0xdfd  :  255 - 0xff
    "11111111", -- 3582 - 0xdfe  :  255 - 0xff
    "11111111", -- 3583 - 0xdff  :  255 - 0xff
    "11111111", -- 3584 - 0xe00  :  255 - 0xff -- Sprite 0xe0
    "11111111", -- 3585 - 0xe01  :  255 - 0xff
    "11111111", -- 3586 - 0xe02  :  255 - 0xff
    "11111111", -- 3587 - 0xe03  :  255 - 0xff
    "11111111", -- 3588 - 0xe04  :  255 - 0xff
    "11111111", -- 3589 - 0xe05  :  255 - 0xff
    "11111111", -- 3590 - 0xe06  :  255 - 0xff
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "11111111", -- 3592 - 0xe08  :  255 - 0xff
    "11111111", -- 3593 - 0xe09  :  255 - 0xff
    "11111111", -- 3594 - 0xe0a  :  255 - 0xff
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "11111111", -- 3596 - 0xe0c  :  255 - 0xff
    "11111111", -- 3597 - 0xe0d  :  255 - 0xff
    "11111111", -- 3598 - 0xe0e  :  255 - 0xff
    "11111111", -- 3599 - 0xe0f  :  255 - 0xff
    "11111111", -- 3600 - 0xe10  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "11111111", -- 3602 - 0xe12  :  255 - 0xff
    "11111111", -- 3603 - 0xe13  :  255 - 0xff
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111111", -- 3605 - 0xe15  :  255 - 0xff
    "11111111", -- 3606 - 0xe16  :  255 - 0xff
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "11111111", -- 3608 - 0xe18  :  255 - 0xff
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "11111111", -- 3610 - 0xe1a  :  255 - 0xff
    "11111111", -- 3611 - 0xe1b  :  255 - 0xff
    "11111111", -- 3612 - 0xe1c  :  255 - 0xff
    "11111111", -- 3613 - 0xe1d  :  255 - 0xff
    "11111111", -- 3614 - 0xe1e  :  255 - 0xff
    "11111111", -- 3615 - 0xe1f  :  255 - 0xff
    "11111111", -- 3616 - 0xe20  :  255 - 0xff -- Sprite 0xe2
    "11111111", -- 3617 - 0xe21  :  255 - 0xff
    "11111111", -- 3618 - 0xe22  :  255 - 0xff
    "11111111", -- 3619 - 0xe23  :  255 - 0xff
    "11111111", -- 3620 - 0xe24  :  255 - 0xff
    "11111111", -- 3621 - 0xe25  :  255 - 0xff
    "11111111", -- 3622 - 0xe26  :  255 - 0xff
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111111", -- 3624 - 0xe28  :  255 - 0xff
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "11111111", -- 3631 - 0xe2f  :  255 - 0xff
    "11111111", -- 3632 - 0xe30  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 3633 - 0xe31  :  255 - 0xff
    "11111111", -- 3634 - 0xe32  :  255 - 0xff
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "11111111", -- 3636 - 0xe34  :  255 - 0xff
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "11111111", -- 3640 - 0xe38  :  255 - 0xff
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "11111111", -- 3642 - 0xe3a  :  255 - 0xff
    "11111111", -- 3643 - 0xe3b  :  255 - 0xff
    "11111111", -- 3644 - 0xe3c  :  255 - 0xff
    "11111111", -- 3645 - 0xe3d  :  255 - 0xff
    "11111111", -- 3646 - 0xe3e  :  255 - 0xff
    "11111111", -- 3647 - 0xe3f  :  255 - 0xff
    "11111111", -- 3648 - 0xe40  :  255 - 0xff -- Sprite 0xe4
    "11111111", -- 3649 - 0xe41  :  255 - 0xff
    "11111111", -- 3650 - 0xe42  :  255 - 0xff
    "11111111", -- 3651 - 0xe43  :  255 - 0xff
    "11111111", -- 3652 - 0xe44  :  255 - 0xff
    "11111111", -- 3653 - 0xe45  :  255 - 0xff
    "11111111", -- 3654 - 0xe46  :  255 - 0xff
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11111111", -- 3656 - 0xe48  :  255 - 0xff
    "11111111", -- 3657 - 0xe49  :  255 - 0xff
    "11111111", -- 3658 - 0xe4a  :  255 - 0xff
    "11111111", -- 3659 - 0xe4b  :  255 - 0xff
    "11111111", -- 3660 - 0xe4c  :  255 - 0xff
    "11111111", -- 3661 - 0xe4d  :  255 - 0xff
    "11111111", -- 3662 - 0xe4e  :  255 - 0xff
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "11111111", -- 3664 - 0xe50  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 3665 - 0xe51  :  255 - 0xff
    "11111111", -- 3666 - 0xe52  :  255 - 0xff
    "11111111", -- 3667 - 0xe53  :  255 - 0xff
    "11111111", -- 3668 - 0xe54  :  255 - 0xff
    "11111111", -- 3669 - 0xe55  :  255 - 0xff
    "11111111", -- 3670 - 0xe56  :  255 - 0xff
    "11111111", -- 3671 - 0xe57  :  255 - 0xff
    "11111111", -- 3672 - 0xe58  :  255 - 0xff
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "11111111", -- 3674 - 0xe5a  :  255 - 0xff
    "11111111", -- 3675 - 0xe5b  :  255 - 0xff
    "11111111", -- 3676 - 0xe5c  :  255 - 0xff
    "11111111", -- 3677 - 0xe5d  :  255 - 0xff
    "11111111", -- 3678 - 0xe5e  :  255 - 0xff
    "11111111", -- 3679 - 0xe5f  :  255 - 0xff
    "11111111", -- 3680 - 0xe60  :  255 - 0xff -- Sprite 0xe6
    "11111111", -- 3681 - 0xe61  :  255 - 0xff
    "11111111", -- 3682 - 0xe62  :  255 - 0xff
    "11111111", -- 3683 - 0xe63  :  255 - 0xff
    "11111111", -- 3684 - 0xe64  :  255 - 0xff
    "11111111", -- 3685 - 0xe65  :  255 - 0xff
    "11111111", -- 3686 - 0xe66  :  255 - 0xff
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "11111111", -- 3688 - 0xe68  :  255 - 0xff
    "11111111", -- 3689 - 0xe69  :  255 - 0xff
    "11111111", -- 3690 - 0xe6a  :  255 - 0xff
    "11111111", -- 3691 - 0xe6b  :  255 - 0xff
    "11111111", -- 3692 - 0xe6c  :  255 - 0xff
    "11111111", -- 3693 - 0xe6d  :  255 - 0xff
    "11111111", -- 3694 - 0xe6e  :  255 - 0xff
    "11111111", -- 3695 - 0xe6f  :  255 - 0xff
    "11111111", -- 3696 - 0xe70  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 3697 - 0xe71  :  255 - 0xff
    "11111111", -- 3698 - 0xe72  :  255 - 0xff
    "11111111", -- 3699 - 0xe73  :  255 - 0xff
    "11111111", -- 3700 - 0xe74  :  255 - 0xff
    "11111111", -- 3701 - 0xe75  :  255 - 0xff
    "11111111", -- 3702 - 0xe76  :  255 - 0xff
    "11111111", -- 3703 - 0xe77  :  255 - 0xff
    "11111111", -- 3704 - 0xe78  :  255 - 0xff
    "11111111", -- 3705 - 0xe79  :  255 - 0xff
    "11111111", -- 3706 - 0xe7a  :  255 - 0xff
    "11111111", -- 3707 - 0xe7b  :  255 - 0xff
    "11111111", -- 3708 - 0xe7c  :  255 - 0xff
    "11111111", -- 3709 - 0xe7d  :  255 - 0xff
    "11111111", -- 3710 - 0xe7e  :  255 - 0xff
    "11111111", -- 3711 - 0xe7f  :  255 - 0xff
    "11111111", -- 3712 - 0xe80  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "11111111", -- 3715 - 0xe83  :  255 - 0xff
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11111111", -- 3720 - 0xe88  :  255 - 0xff
    "11111111", -- 3721 - 0xe89  :  255 - 0xff
    "11111111", -- 3722 - 0xe8a  :  255 - 0xff
    "11111111", -- 3723 - 0xe8b  :  255 - 0xff
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11111111", -- 3728 - 0xe90  :  255 - 0xff -- Sprite 0xe9
    "11111111", -- 3729 - 0xe91  :  255 - 0xff
    "11111111", -- 3730 - 0xe92  :  255 - 0xff
    "11111111", -- 3731 - 0xe93  :  255 - 0xff
    "11111111", -- 3732 - 0xe94  :  255 - 0xff
    "11111111", -- 3733 - 0xe95  :  255 - 0xff
    "11111111", -- 3734 - 0xe96  :  255 - 0xff
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111111", -- 3736 - 0xe98  :  255 - 0xff
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111111", -- 3740 - 0xe9c  :  255 - 0xff
    "11111111", -- 3741 - 0xe9d  :  255 - 0xff
    "11111111", -- 3742 - 0xe9e  :  255 - 0xff
    "11111111", -- 3743 - 0xe9f  :  255 - 0xff
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "11111111", -- 3748 - 0xea4  :  255 - 0xff
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "11111111", -- 3751 - 0xea7  :  255 - 0xff
    "11111111", -- 3752 - 0xea8  :  255 - 0xff
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "11111111", -- 3760 - 0xeb0  :  255 - 0xff -- Sprite 0xeb
    "11111111", -- 3761 - 0xeb1  :  255 - 0xff
    "11111111", -- 3762 - 0xeb2  :  255 - 0xff
    "11111111", -- 3763 - 0xeb3  :  255 - 0xff
    "11111111", -- 3764 - 0xeb4  :  255 - 0xff
    "11111111", -- 3765 - 0xeb5  :  255 - 0xff
    "11111111", -- 3766 - 0xeb6  :  255 - 0xff
    "11111111", -- 3767 - 0xeb7  :  255 - 0xff
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "11111111", -- 3772 - 0xebc  :  255 - 0xff
    "11111111", -- 3773 - 0xebd  :  255 - 0xff
    "11111111", -- 3774 - 0xebe  :  255 - 0xff
    "11111111", -- 3775 - 0xebf  :  255 - 0xff
    "11111111", -- 3776 - 0xec0  :  255 - 0xff -- Sprite 0xec
    "11111111", -- 3777 - 0xec1  :  255 - 0xff
    "11111111", -- 3778 - 0xec2  :  255 - 0xff
    "11111111", -- 3779 - 0xec3  :  255 - 0xff
    "11111111", -- 3780 - 0xec4  :  255 - 0xff
    "11111111", -- 3781 - 0xec5  :  255 - 0xff
    "11111111", -- 3782 - 0xec6  :  255 - 0xff
    "11111111", -- 3783 - 0xec7  :  255 - 0xff
    "11111111", -- 3784 - 0xec8  :  255 - 0xff
    "11111111", -- 3785 - 0xec9  :  255 - 0xff
    "11111111", -- 3786 - 0xeca  :  255 - 0xff
    "11111111", -- 3787 - 0xecb  :  255 - 0xff
    "11111111", -- 3788 - 0xecc  :  255 - 0xff
    "11111111", -- 3789 - 0xecd  :  255 - 0xff
    "11111111", -- 3790 - 0xece  :  255 - 0xff
    "11111111", -- 3791 - 0xecf  :  255 - 0xff
    "11111111", -- 3792 - 0xed0  :  255 - 0xff -- Sprite 0xed
    "11111111", -- 3793 - 0xed1  :  255 - 0xff
    "11111111", -- 3794 - 0xed2  :  255 - 0xff
    "11111111", -- 3795 - 0xed3  :  255 - 0xff
    "11111111", -- 3796 - 0xed4  :  255 - 0xff
    "11111111", -- 3797 - 0xed5  :  255 - 0xff
    "11111111", -- 3798 - 0xed6  :  255 - 0xff
    "11111111", -- 3799 - 0xed7  :  255 - 0xff
    "11111111", -- 3800 - 0xed8  :  255 - 0xff
    "11111111", -- 3801 - 0xed9  :  255 - 0xff
    "11111111", -- 3802 - 0xeda  :  255 - 0xff
    "11111111", -- 3803 - 0xedb  :  255 - 0xff
    "11111111", -- 3804 - 0xedc  :  255 - 0xff
    "11111111", -- 3805 - 0xedd  :  255 - 0xff
    "11111111", -- 3806 - 0xede  :  255 - 0xff
    "11111111", -- 3807 - 0xedf  :  255 - 0xff
    "11111111", -- 3808 - 0xee0  :  255 - 0xff -- Sprite 0xee
    "11111111", -- 3809 - 0xee1  :  255 - 0xff
    "11111111", -- 3810 - 0xee2  :  255 - 0xff
    "11111111", -- 3811 - 0xee3  :  255 - 0xff
    "11111111", -- 3812 - 0xee4  :  255 - 0xff
    "11111111", -- 3813 - 0xee5  :  255 - 0xff
    "11111111", -- 3814 - 0xee6  :  255 - 0xff
    "11111111", -- 3815 - 0xee7  :  255 - 0xff
    "11111111", -- 3816 - 0xee8  :  255 - 0xff
    "11111111", -- 3817 - 0xee9  :  255 - 0xff
    "11111111", -- 3818 - 0xeea  :  255 - 0xff
    "11111111", -- 3819 - 0xeeb  :  255 - 0xff
    "11111111", -- 3820 - 0xeec  :  255 - 0xff
    "11111111", -- 3821 - 0xeed  :  255 - 0xff
    "11111111", -- 3822 - 0xeee  :  255 - 0xff
    "11111111", -- 3823 - 0xeef  :  255 - 0xff
    "11111111", -- 3824 - 0xef0  :  255 - 0xff -- Sprite 0xef
    "11111111", -- 3825 - 0xef1  :  255 - 0xff
    "11111111", -- 3826 - 0xef2  :  255 - 0xff
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11111111", -- 3828 - 0xef4  :  255 - 0xff
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11111111", -- 3830 - 0xef6  :  255 - 0xff
    "11111111", -- 3831 - 0xef7  :  255 - 0xff
    "11111111", -- 3832 - 0xef8  :  255 - 0xff
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "11111111", -- 3834 - 0xefa  :  255 - 0xff
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111111", -- 3836 - 0xefc  :  255 - 0xff
    "11111111", -- 3837 - 0xefd  :  255 - 0xff
    "11111111", -- 3838 - 0xefe  :  255 - 0xff
    "11111111", -- 3839 - 0xeff  :  255 - 0xff
    "11111111", -- 3840 - 0xf00  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 3841 - 0xf01  :  255 - 0xff
    "11111111", -- 3842 - 0xf02  :  255 - 0xff
    "11111111", -- 3843 - 0xf03  :  255 - 0xff
    "11111111", -- 3844 - 0xf04  :  255 - 0xff
    "11111111", -- 3845 - 0xf05  :  255 - 0xff
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11111111", -- 3848 - 0xf08  :  255 - 0xff
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "11111111", -- 3850 - 0xf0a  :  255 - 0xff
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "11111111", -- 3860 - 0xf14  :  255 - 0xff
    "11111111", -- 3861 - 0xf15  :  255 - 0xff
    "11111111", -- 3862 - 0xf16  :  255 - 0xff
    "11111111", -- 3863 - 0xf17  :  255 - 0xff
    "11111111", -- 3864 - 0xf18  :  255 - 0xff
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11111111", -- 3867 - 0xf1b  :  255 - 0xff
    "11111111", -- 3868 - 0xf1c  :  255 - 0xff
    "11111111", -- 3869 - 0xf1d  :  255 - 0xff
    "11111111", -- 3870 - 0xf1e  :  255 - 0xff
    "11111111", -- 3871 - 0xf1f  :  255 - 0xff
    "11111111", -- 3872 - 0xf20  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 3873 - 0xf21  :  255 - 0xff
    "11111111", -- 3874 - 0xf22  :  255 - 0xff
    "11111111", -- 3875 - 0xf23  :  255 - 0xff
    "11111111", -- 3876 - 0xf24  :  255 - 0xff
    "11111111", -- 3877 - 0xf25  :  255 - 0xff
    "11111111", -- 3878 - 0xf26  :  255 - 0xff
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11111111", -- 3883 - 0xf2b  :  255 - 0xff
    "11111111", -- 3884 - 0xf2c  :  255 - 0xff
    "11111111", -- 3885 - 0xf2d  :  255 - 0xff
    "11111111", -- 3886 - 0xf2e  :  255 - 0xff
    "11111111", -- 3887 - 0xf2f  :  255 - 0xff
    "11111111", -- 3888 - 0xf30  :  255 - 0xff -- Sprite 0xf3
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "11111111", -- 3891 - 0xf33  :  255 - 0xff
    "11111111", -- 3892 - 0xf34  :  255 - 0xff
    "11111111", -- 3893 - 0xf35  :  255 - 0xff
    "11111111", -- 3894 - 0xf36  :  255 - 0xff
    "11111111", -- 3895 - 0xf37  :  255 - 0xff
    "11111111", -- 3896 - 0xf38  :  255 - 0xff
    "11111111", -- 3897 - 0xf39  :  255 - 0xff
    "11111111", -- 3898 - 0xf3a  :  255 - 0xff
    "11111111", -- 3899 - 0xf3b  :  255 - 0xff
    "11111111", -- 3900 - 0xf3c  :  255 - 0xff
    "11111111", -- 3901 - 0xf3d  :  255 - 0xff
    "11111111", -- 3902 - 0xf3e  :  255 - 0xff
    "11111111", -- 3903 - 0xf3f  :  255 - 0xff
    "11111111", -- 3904 - 0xf40  :  255 - 0xff -- Sprite 0xf4
    "11111111", -- 3905 - 0xf41  :  255 - 0xff
    "11111111", -- 3906 - 0xf42  :  255 - 0xff
    "11111111", -- 3907 - 0xf43  :  255 - 0xff
    "11111111", -- 3908 - 0xf44  :  255 - 0xff
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "11111111", -- 3912 - 0xf48  :  255 - 0xff
    "11111111", -- 3913 - 0xf49  :  255 - 0xff
    "11111111", -- 3914 - 0xf4a  :  255 - 0xff
    "11111111", -- 3915 - 0xf4b  :  255 - 0xff
    "11111111", -- 3916 - 0xf4c  :  255 - 0xff
    "11111111", -- 3917 - 0xf4d  :  255 - 0xff
    "11111111", -- 3918 - 0xf4e  :  255 - 0xff
    "11111111", -- 3919 - 0xf4f  :  255 - 0xff
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Sprite 0xf5
    "11111111", -- 3921 - 0xf51  :  255 - 0xff
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "11111111", -- 3923 - 0xf53  :  255 - 0xff
    "11111111", -- 3924 - 0xf54  :  255 - 0xff
    "11111111", -- 3925 - 0xf55  :  255 - 0xff
    "11111111", -- 3926 - 0xf56  :  255 - 0xff
    "11111111", -- 3927 - 0xf57  :  255 - 0xff
    "11111111", -- 3928 - 0xf58  :  255 - 0xff
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "11111111", -- 3931 - 0xf5b  :  255 - 0xff
    "11111111", -- 3932 - 0xf5c  :  255 - 0xff
    "11111111", -- 3933 - 0xf5d  :  255 - 0xff
    "11111111", -- 3934 - 0xf5e  :  255 - 0xff
    "11111111", -- 3935 - 0xf5f  :  255 - 0xff
    "11111111", -- 3936 - 0xf60  :  255 - 0xff -- Sprite 0xf6
    "11111111", -- 3937 - 0xf61  :  255 - 0xff
    "11111111", -- 3938 - 0xf62  :  255 - 0xff
    "11111111", -- 3939 - 0xf63  :  255 - 0xff
    "11111111", -- 3940 - 0xf64  :  255 - 0xff
    "11111111", -- 3941 - 0xf65  :  255 - 0xff
    "11111111", -- 3942 - 0xf66  :  255 - 0xff
    "11111111", -- 3943 - 0xf67  :  255 - 0xff
    "11111111", -- 3944 - 0xf68  :  255 - 0xff
    "11111111", -- 3945 - 0xf69  :  255 - 0xff
    "11111111", -- 3946 - 0xf6a  :  255 - 0xff
    "11111111", -- 3947 - 0xf6b  :  255 - 0xff
    "11111111", -- 3948 - 0xf6c  :  255 - 0xff
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "11111111", -- 3952 - 0xf70  :  255 - 0xff -- Sprite 0xf7
    "11111111", -- 3953 - 0xf71  :  255 - 0xff
    "11111111", -- 3954 - 0xf72  :  255 - 0xff
    "11111111", -- 3955 - 0xf73  :  255 - 0xff
    "11111111", -- 3956 - 0xf74  :  255 - 0xff
    "11111111", -- 3957 - 0xf75  :  255 - 0xff
    "11111111", -- 3958 - 0xf76  :  255 - 0xff
    "11111111", -- 3959 - 0xf77  :  255 - 0xff
    "11111111", -- 3960 - 0xf78  :  255 - 0xff
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "11111111", -- 3968 - 0xf80  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "11111111", -- 3970 - 0xf82  :  255 - 0xff
    "11111111", -- 3971 - 0xf83  :  255 - 0xff
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "11111111", -- 3974 - 0xf86  :  255 - 0xff
    "11111111", -- 3975 - 0xf87  :  255 - 0xff
    "11111111", -- 3976 - 0xf88  :  255 - 0xff
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111111", -- 3982 - 0xf8e  :  255 - 0xff
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "11111111", -- 3992 - 0xf98  :  255 - 0xff
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111111", -- 3999 - 0xf9f  :  255 - 0xff
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "11111111", -- 4007 - 0xfa7  :  255 - 0xff
    "11111111", -- 4008 - 0xfa8  :  255 - 0xff
    "11111111", -- 4009 - 0xfa9  :  255 - 0xff
    "11111111", -- 4010 - 0xfaa  :  255 - 0xff
    "11111111", -- 4011 - 0xfab  :  255 - 0xff
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "11111111", -- 4015 - 0xfaf  :  255 - 0xff
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "11111111", -- 4024 - 0xfb8  :  255 - 0xff
    "11111111", -- 4025 - 0xfb9  :  255 - 0xff
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "11111111", -- 4031 - 0xfbf  :  255 - 0xff
    "11111111", -- 4032 - 0xfc0  :  255 - 0xff -- Sprite 0xfc
    "11111111", -- 4033 - 0xfc1  :  255 - 0xff
    "11111111", -- 4034 - 0xfc2  :  255 - 0xff
    "11111111", -- 4035 - 0xfc3  :  255 - 0xff
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "11111111", -- 4040 - 0xfc8  :  255 - 0xff
    "11111111", -- 4041 - 0xfc9  :  255 - 0xff
    "11111111", -- 4042 - 0xfca  :  255 - 0xff
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "11111111", -- 4048 - 0xfd0  :  255 - 0xff -- Sprite 0xfd
    "11111111", -- 4049 - 0xfd1  :  255 - 0xff
    "11111111", -- 4050 - 0xfd2  :  255 - 0xff
    "11111111", -- 4051 - 0xfd3  :  255 - 0xff
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "11111111", -- 4064 - 0xfe0  :  255 - 0xff -- Sprite 0xfe
    "11111111", -- 4065 - 0xfe1  :  255 - 0xff
    "11111111", -- 4066 - 0xfe2  :  255 - 0xff
    "11111111", -- 4067 - 0xfe3  :  255 - 0xff
    "11111111", -- 4068 - 0xfe4  :  255 - 0xff
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11111111", -- 4075 - 0xfeb  :  255 - 0xff
    "11111111", -- 4076 - 0xfec  :  255 - 0xff
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111", -- 4095 - 0xfff  :  255 - 0xff
          -- Pattern Table 1---------
    "00000000", -- 4096 - 0x1000  :    0 - 0x0 -- Background 0x0
    "00000000", -- 4097 - 0x1001  :    0 - 0x0
    "00000000", -- 4098 - 0x1002  :    0 - 0x0
    "00000000", -- 4099 - 0x1003  :    0 - 0x0
    "00000000", -- 4100 - 0x1004  :    0 - 0x0
    "00000000", -- 4101 - 0x1005  :    0 - 0x0
    "00000000", -- 4102 - 0x1006  :    0 - 0x0
    "00000000", -- 4103 - 0x1007  :    0 - 0x0
    "00000000", -- 4104 - 0x1008  :    0 - 0x0
    "00000000", -- 4105 - 0x1009  :    0 - 0x0
    "00000000", -- 4106 - 0x100a  :    0 - 0x0
    "00000000", -- 4107 - 0x100b  :    0 - 0x0
    "00000000", -- 4108 - 0x100c  :    0 - 0x0
    "00000000", -- 4109 - 0x100d  :    0 - 0x0
    "00000000", -- 4110 - 0x100e  :    0 - 0x0
    "00000000", -- 4111 - 0x100f  :    0 - 0x0
    "00000000", -- 4112 - 0x1010  :    0 - 0x0 -- Background 0x1
    "00111000", -- 4113 - 0x1011  :   56 - 0x38
    "01111100", -- 4114 - 0x1012  :  124 - 0x7c
    "11111110", -- 4115 - 0x1013  :  254 - 0xfe
    "11111110", -- 4116 - 0x1014  :  254 - 0xfe
    "11111110", -- 4117 - 0x1015  :  254 - 0xfe
    "01111100", -- 4118 - 0x1016  :  124 - 0x7c
    "00111000", -- 4119 - 0x1017  :   56 - 0x38
    "00000000", -- 4120 - 0x1018  :    0 - 0x0
    "00111000", -- 4121 - 0x1019  :   56 - 0x38
    "01111100", -- 4122 - 0x101a  :  124 - 0x7c
    "11111110", -- 4123 - 0x101b  :  254 - 0xfe
    "11111110", -- 4124 - 0x101c  :  254 - 0xfe
    "11111110", -- 4125 - 0x101d  :  254 - 0xfe
    "01111100", -- 4126 - 0x101e  :  124 - 0x7c
    "00111000", -- 4127 - 0x101f  :   56 - 0x38
    "00000000", -- 4128 - 0x1020  :    0 - 0x0 -- Background 0x2
    "00000000", -- 4129 - 0x1021  :    0 - 0x0
    "00000000", -- 4130 - 0x1022  :    0 - 0x0
    "00000000", -- 4131 - 0x1023  :    0 - 0x0
    "00000000", -- 4132 - 0x1024  :    0 - 0x0
    "00000000", -- 4133 - 0x1025  :    0 - 0x0
    "00000000", -- 4134 - 0x1026  :    0 - 0x0
    "00000000", -- 4135 - 0x1027  :    0 - 0x0
    "00000000", -- 4136 - 0x1028  :    0 - 0x0
    "00000000", -- 4137 - 0x1029  :    0 - 0x0
    "00000000", -- 4138 - 0x102a  :    0 - 0x0
    "00000000", -- 4139 - 0x102b  :    0 - 0x0
    "00000000", -- 4140 - 0x102c  :    0 - 0x0
    "00000000", -- 4141 - 0x102d  :    0 - 0x0
    "00000000", -- 4142 - 0x102e  :    0 - 0x0
    "00000000", -- 4143 - 0x102f  :    0 - 0x0
    "00000000", -- 4144 - 0x1030  :    0 - 0x0 -- Background 0x3
    "00000000", -- 4145 - 0x1031  :    0 - 0x0
    "00000000", -- 4146 - 0x1032  :    0 - 0x0
    "00011000", -- 4147 - 0x1033  :   24 - 0x18
    "00011000", -- 4148 - 0x1034  :   24 - 0x18
    "00000000", -- 4149 - 0x1035  :    0 - 0x0
    "00000000", -- 4150 - 0x1036  :    0 - 0x0
    "00000000", -- 4151 - 0x1037  :    0 - 0x0
    "00000000", -- 4152 - 0x1038  :    0 - 0x0
    "00000000", -- 4153 - 0x1039  :    0 - 0x0
    "00000000", -- 4154 - 0x103a  :    0 - 0x0
    "00011000", -- 4155 - 0x103b  :   24 - 0x18
    "00011000", -- 4156 - 0x103c  :   24 - 0x18
    "00000000", -- 4157 - 0x103d  :    0 - 0x0
    "00000000", -- 4158 - 0x103e  :    0 - 0x0
    "00000000", -- 4159 - 0x103f  :    0 - 0x0
    "00000000", -- 4160 - 0x1040  :    0 - 0x0 -- Background 0x4
    "00000000", -- 4161 - 0x1041  :    0 - 0x0
    "00000000", -- 4162 - 0x1042  :    0 - 0x0
    "00000000", -- 4163 - 0x1043  :    0 - 0x0
    "00000000", -- 4164 - 0x1044  :    0 - 0x0
    "00000000", -- 4165 - 0x1045  :    0 - 0x0
    "00000000", -- 4166 - 0x1046  :    0 - 0x0
    "00000000", -- 4167 - 0x1047  :    0 - 0x0
    "11111111", -- 4168 - 0x1048  :  255 - 0xff
    "11111111", -- 4169 - 0x1049  :  255 - 0xff
    "11111111", -- 4170 - 0x104a  :  255 - 0xff
    "11111111", -- 4171 - 0x104b  :  255 - 0xff
    "11111111", -- 4172 - 0x104c  :  255 - 0xff
    "11111111", -- 4173 - 0x104d  :  255 - 0xff
    "11111111", -- 4174 - 0x104e  :  255 - 0xff
    "11111111", -- 4175 - 0x104f  :  255 - 0xff
    "00000000", -- 4176 - 0x1050  :    0 - 0x0 -- Background 0x5
    "00000000", -- 4177 - 0x1051  :    0 - 0x0
    "00000000", -- 4178 - 0x1052  :    0 - 0x0
    "00000000", -- 4179 - 0x1053  :    0 - 0x0
    "00000000", -- 4180 - 0x1054  :    0 - 0x0
    "00000000", -- 4181 - 0x1055  :    0 - 0x0
    "00000000", -- 4182 - 0x1056  :    0 - 0x0
    "00000000", -- 4183 - 0x1057  :    0 - 0x0
    "00001111", -- 4184 - 0x1058  :   15 - 0xf
    "00001111", -- 4185 - 0x1059  :   15 - 0xf
    "00001111", -- 4186 - 0x105a  :   15 - 0xf
    "00001111", -- 4187 - 0x105b  :   15 - 0xf
    "00001111", -- 4188 - 0x105c  :   15 - 0xf
    "00001111", -- 4189 - 0x105d  :   15 - 0xf
    "00001111", -- 4190 - 0x105e  :   15 - 0xf
    "00001111", -- 4191 - 0x105f  :   15 - 0xf
    "00000000", -- 4192 - 0x1060  :    0 - 0x0 -- Background 0x6
    "00000000", -- 4193 - 0x1061  :    0 - 0x0
    "00000000", -- 4194 - 0x1062  :    0 - 0x0
    "00000000", -- 4195 - 0x1063  :    0 - 0x0
    "00000000", -- 4196 - 0x1064  :    0 - 0x0
    "00000000", -- 4197 - 0x1065  :    0 - 0x0
    "00000000", -- 4198 - 0x1066  :    0 - 0x0
    "00000000", -- 4199 - 0x1067  :    0 - 0x0
    "11110000", -- 4200 - 0x1068  :  240 - 0xf0
    "11110000", -- 4201 - 0x1069  :  240 - 0xf0
    "11110000", -- 4202 - 0x106a  :  240 - 0xf0
    "11110000", -- 4203 - 0x106b  :  240 - 0xf0
    "11110000", -- 4204 - 0x106c  :  240 - 0xf0
    "11110000", -- 4205 - 0x106d  :  240 - 0xf0
    "11110000", -- 4206 - 0x106e  :  240 - 0xf0
    "11110000", -- 4207 - 0x106f  :  240 - 0xf0
    "00000000", -- 4208 - 0x1070  :    0 - 0x0 -- Background 0x7
    "00000000", -- 4209 - 0x1071  :    0 - 0x0
    "00000000", -- 4210 - 0x1072  :    0 - 0x0
    "00000000", -- 4211 - 0x1073  :    0 - 0x0
    "00000000", -- 4212 - 0x1074  :    0 - 0x0
    "00000000", -- 4213 - 0x1075  :    0 - 0x0
    "00000000", -- 4214 - 0x1076  :    0 - 0x0
    "00000000", -- 4215 - 0x1077  :    0 - 0x0
    "00000000", -- 4216 - 0x1078  :    0 - 0x0
    "00000000", -- 4217 - 0x1079  :    0 - 0x0
    "00000000", -- 4218 - 0x107a  :    0 - 0x0
    "00000000", -- 4219 - 0x107b  :    0 - 0x0
    "00000000", -- 4220 - 0x107c  :    0 - 0x0
    "00000000", -- 4221 - 0x107d  :    0 - 0x0
    "00000000", -- 4222 - 0x107e  :    0 - 0x0
    "00000000", -- 4223 - 0x107f  :    0 - 0x0
    "00000000", -- 4224 - 0x1080  :    0 - 0x0 -- Background 0x8
    "00000000", -- 4225 - 0x1081  :    0 - 0x0
    "00000000", -- 4226 - 0x1082  :    0 - 0x0
    "00000000", -- 4227 - 0x1083  :    0 - 0x0
    "00000000", -- 4228 - 0x1084  :    0 - 0x0
    "00000000", -- 4229 - 0x1085  :    0 - 0x0
    "00000000", -- 4230 - 0x1086  :    0 - 0x0
    "00000000", -- 4231 - 0x1087  :    0 - 0x0
    "00000000", -- 4232 - 0x1088  :    0 - 0x0
    "00000000", -- 4233 - 0x1089  :    0 - 0x0
    "00000000", -- 4234 - 0x108a  :    0 - 0x0
    "00000000", -- 4235 - 0x108b  :    0 - 0x0
    "00000000", -- 4236 - 0x108c  :    0 - 0x0
    "00000000", -- 4237 - 0x108d  :    0 - 0x0
    "00000000", -- 4238 - 0x108e  :    0 - 0x0
    "00000000", -- 4239 - 0x108f  :    0 - 0x0
    "00000000", -- 4240 - 0x1090  :    0 - 0x0 -- Background 0x9
    "00000000", -- 4241 - 0x1091  :    0 - 0x0
    "00000000", -- 4242 - 0x1092  :    0 - 0x0
    "00011000", -- 4243 - 0x1093  :   24 - 0x18
    "00011000", -- 4244 - 0x1094  :   24 - 0x18
    "00000000", -- 4245 - 0x1095  :    0 - 0x0
    "00000000", -- 4246 - 0x1096  :    0 - 0x0
    "00000000", -- 4247 - 0x1097  :    0 - 0x0
    "00000000", -- 4248 - 0x1098  :    0 - 0x0
    "00000000", -- 4249 - 0x1099  :    0 - 0x0
    "00000000", -- 4250 - 0x109a  :    0 - 0x0
    "00011000", -- 4251 - 0x109b  :   24 - 0x18
    "00011000", -- 4252 - 0x109c  :   24 - 0x18
    "00000000", -- 4253 - 0x109d  :    0 - 0x0
    "00000000", -- 4254 - 0x109e  :    0 - 0x0
    "00000000", -- 4255 - 0x109f  :    0 - 0x0
    "00000000", -- 4256 - 0x10a0  :    0 - 0x0 -- Background 0xa
    "00000000", -- 4257 - 0x10a1  :    0 - 0x0
    "00000000", -- 4258 - 0x10a2  :    0 - 0x0
    "00000000", -- 4259 - 0x10a3  :    0 - 0x0
    "00000000", -- 4260 - 0x10a4  :    0 - 0x0
    "00000000", -- 4261 - 0x10a5  :    0 - 0x0
    "00000000", -- 4262 - 0x10a6  :    0 - 0x0
    "00000000", -- 4263 - 0x10a7  :    0 - 0x0
    "00000000", -- 4264 - 0x10a8  :    0 - 0x0
    "00000000", -- 4265 - 0x10a9  :    0 - 0x0
    "00000000", -- 4266 - 0x10aa  :    0 - 0x0
    "00000000", -- 4267 - 0x10ab  :    0 - 0x0
    "00000000", -- 4268 - 0x10ac  :    0 - 0x0
    "00000000", -- 4269 - 0x10ad  :    0 - 0x0
    "00000000", -- 4270 - 0x10ae  :    0 - 0x0
    "00000000", -- 4271 - 0x10af  :    0 - 0x0
    "00000000", -- 4272 - 0x10b0  :    0 - 0x0 -- Background 0xb
    "00000000", -- 4273 - 0x10b1  :    0 - 0x0
    "00000000", -- 4274 - 0x10b2  :    0 - 0x0
    "00000000", -- 4275 - 0x10b3  :    0 - 0x0
    "00000000", -- 4276 - 0x10b4  :    0 - 0x0
    "00000000", -- 4277 - 0x10b5  :    0 - 0x0
    "00000000", -- 4278 - 0x10b6  :    0 - 0x0
    "00000000", -- 4279 - 0x10b7  :    0 - 0x0
    "00000000", -- 4280 - 0x10b8  :    0 - 0x0
    "00000000", -- 4281 - 0x10b9  :    0 - 0x0
    "00000000", -- 4282 - 0x10ba  :    0 - 0x0
    "00000000", -- 4283 - 0x10bb  :    0 - 0x0
    "00000000", -- 4284 - 0x10bc  :    0 - 0x0
    "00000000", -- 4285 - 0x10bd  :    0 - 0x0
    "00000000", -- 4286 - 0x10be  :    0 - 0x0
    "00000000", -- 4287 - 0x10bf  :    0 - 0x0
    "00000000", -- 4288 - 0x10c0  :    0 - 0x0 -- Background 0xc
    "00000000", -- 4289 - 0x10c1  :    0 - 0x0
    "00000000", -- 4290 - 0x10c2  :    0 - 0x0
    "00000000", -- 4291 - 0x10c3  :    0 - 0x0
    "00000000", -- 4292 - 0x10c4  :    0 - 0x0
    "00000000", -- 4293 - 0x10c5  :    0 - 0x0
    "00000000", -- 4294 - 0x10c6  :    0 - 0x0
    "00000000", -- 4295 - 0x10c7  :    0 - 0x0
    "00000000", -- 4296 - 0x10c8  :    0 - 0x0
    "00000000", -- 4297 - 0x10c9  :    0 - 0x0
    "00000000", -- 4298 - 0x10ca  :    0 - 0x0
    "00000000", -- 4299 - 0x10cb  :    0 - 0x0
    "00000000", -- 4300 - 0x10cc  :    0 - 0x0
    "00000000", -- 4301 - 0x10cd  :    0 - 0x0
    "00000000", -- 4302 - 0x10ce  :    0 - 0x0
    "00000000", -- 4303 - 0x10cf  :    0 - 0x0
    "00000000", -- 4304 - 0x10d0  :    0 - 0x0 -- Background 0xd
    "00000000", -- 4305 - 0x10d1  :    0 - 0x0
    "00000000", -- 4306 - 0x10d2  :    0 - 0x0
    "00000000", -- 4307 - 0x10d3  :    0 - 0x0
    "00000000", -- 4308 - 0x10d4  :    0 - 0x0
    "00000000", -- 4309 - 0x10d5  :    0 - 0x0
    "00000000", -- 4310 - 0x10d6  :    0 - 0x0
    "00000000", -- 4311 - 0x10d7  :    0 - 0x0
    "00000000", -- 4312 - 0x10d8  :    0 - 0x0
    "00000000", -- 4313 - 0x10d9  :    0 - 0x0
    "00000000", -- 4314 - 0x10da  :    0 - 0x0
    "00000000", -- 4315 - 0x10db  :    0 - 0x0
    "00000000", -- 4316 - 0x10dc  :    0 - 0x0
    "00000000", -- 4317 - 0x10dd  :    0 - 0x0
    "00000000", -- 4318 - 0x10de  :    0 - 0x0
    "00000000", -- 4319 - 0x10df  :    0 - 0x0
    "00000000", -- 4320 - 0x10e0  :    0 - 0x0 -- Background 0xe
    "00000000", -- 4321 - 0x10e1  :    0 - 0x0
    "00000000", -- 4322 - 0x10e2  :    0 - 0x0
    "00000000", -- 4323 - 0x10e3  :    0 - 0x0
    "00000000", -- 4324 - 0x10e4  :    0 - 0x0
    "00000000", -- 4325 - 0x10e5  :    0 - 0x0
    "00000000", -- 4326 - 0x10e6  :    0 - 0x0
    "00000000", -- 4327 - 0x10e7  :    0 - 0x0
    "00000000", -- 4328 - 0x10e8  :    0 - 0x0
    "00000000", -- 4329 - 0x10e9  :    0 - 0x0
    "00000000", -- 4330 - 0x10ea  :    0 - 0x0
    "00000000", -- 4331 - 0x10eb  :    0 - 0x0
    "00000000", -- 4332 - 0x10ec  :    0 - 0x0
    "00000000", -- 4333 - 0x10ed  :    0 - 0x0
    "00000000", -- 4334 - 0x10ee  :    0 - 0x0
    "00000000", -- 4335 - 0x10ef  :    0 - 0x0
    "00000000", -- 4336 - 0x10f0  :    0 - 0x0 -- Background 0xf
    "00000000", -- 4337 - 0x10f1  :    0 - 0x0
    "00000000", -- 4338 - 0x10f2  :    0 - 0x0
    "00000000", -- 4339 - 0x10f3  :    0 - 0x0
    "00000000", -- 4340 - 0x10f4  :    0 - 0x0
    "00000000", -- 4341 - 0x10f5  :    0 - 0x0
    "00000000", -- 4342 - 0x10f6  :    0 - 0x0
    "00000000", -- 4343 - 0x10f7  :    0 - 0x0
    "00000000", -- 4344 - 0x10f8  :    0 - 0x0
    "00000000", -- 4345 - 0x10f9  :    0 - 0x0
    "00000000", -- 4346 - 0x10fa  :    0 - 0x0
    "00000000", -- 4347 - 0x10fb  :    0 - 0x0
    "00000000", -- 4348 - 0x10fc  :    0 - 0x0
    "00000000", -- 4349 - 0x10fd  :    0 - 0x0
    "00000000", -- 4350 - 0x10fe  :    0 - 0x0
    "00000000", -- 4351 - 0x10ff  :    0 - 0x0
    "00000000", -- 4352 - 0x1100  :    0 - 0x0 -- Background 0x10
    "00000000", -- 4353 - 0x1101  :    0 - 0x0
    "11111111", -- 4354 - 0x1102  :  255 - 0xff
    "00000000", -- 4355 - 0x1103  :    0 - 0x0
    "00000000", -- 4356 - 0x1104  :    0 - 0x0
    "11111111", -- 4357 - 0x1105  :  255 - 0xff
    "00000000", -- 4358 - 0x1106  :    0 - 0x0
    "00000000", -- 4359 - 0x1107  :    0 - 0x0
    "00000000", -- 4360 - 0x1108  :    0 - 0x0
    "00000000", -- 4361 - 0x1109  :    0 - 0x0
    "00000000", -- 4362 - 0x110a  :    0 - 0x0
    "00000000", -- 4363 - 0x110b  :    0 - 0x0
    "00000000", -- 4364 - 0x110c  :    0 - 0x0
    "00000000", -- 4365 - 0x110d  :    0 - 0x0
    "00000000", -- 4366 - 0x110e  :    0 - 0x0
    "00000000", -- 4367 - 0x110f  :    0 - 0x0
    "00100100", -- 4368 - 0x1110  :   36 - 0x24 -- Background 0x11
    "00100100", -- 4369 - 0x1111  :   36 - 0x24
    "00100100", -- 4370 - 0x1112  :   36 - 0x24
    "00100100", -- 4371 - 0x1113  :   36 - 0x24
    "00100100", -- 4372 - 0x1114  :   36 - 0x24
    "00100100", -- 4373 - 0x1115  :   36 - 0x24
    "00100100", -- 4374 - 0x1116  :   36 - 0x24
    "00100100", -- 4375 - 0x1117  :   36 - 0x24
    "00000000", -- 4376 - 0x1118  :    0 - 0x0
    "00000000", -- 4377 - 0x1119  :    0 - 0x0
    "00000000", -- 4378 - 0x111a  :    0 - 0x0
    "00000000", -- 4379 - 0x111b  :    0 - 0x0
    "00000000", -- 4380 - 0x111c  :    0 - 0x0
    "00000000", -- 4381 - 0x111d  :    0 - 0x0
    "00000000", -- 4382 - 0x111e  :    0 - 0x0
    "00000000", -- 4383 - 0x111f  :    0 - 0x0
    "00100100", -- 4384 - 0x1120  :   36 - 0x24 -- Background 0x12
    "00100100", -- 4385 - 0x1121  :   36 - 0x24
    "11000011", -- 4386 - 0x1122  :  195 - 0xc3
    "00000000", -- 4387 - 0x1123  :    0 - 0x0
    "00000000", -- 4388 - 0x1124  :    0 - 0x0
    "11111111", -- 4389 - 0x1125  :  255 - 0xff
    "00000000", -- 4390 - 0x1126  :    0 - 0x0
    "00000000", -- 4391 - 0x1127  :    0 - 0x0
    "00000000", -- 4392 - 0x1128  :    0 - 0x0
    "00000000", -- 4393 - 0x1129  :    0 - 0x0
    "00000000", -- 4394 - 0x112a  :    0 - 0x0
    "00000000", -- 4395 - 0x112b  :    0 - 0x0
    "00000000", -- 4396 - 0x112c  :    0 - 0x0
    "00000000", -- 4397 - 0x112d  :    0 - 0x0
    "00000000", -- 4398 - 0x112e  :    0 - 0x0
    "00000000", -- 4399 - 0x112f  :    0 - 0x0
    "00000000", -- 4400 - 0x1130  :    0 - 0x0 -- Background 0x13
    "00000000", -- 4401 - 0x1131  :    0 - 0x0
    "11111111", -- 4402 - 0x1132  :  255 - 0xff
    "00000000", -- 4403 - 0x1133  :    0 - 0x0
    "00000000", -- 4404 - 0x1134  :    0 - 0x0
    "11000011", -- 4405 - 0x1135  :  195 - 0xc3
    "00100100", -- 4406 - 0x1136  :   36 - 0x24
    "00100100", -- 4407 - 0x1137  :   36 - 0x24
    "00000000", -- 4408 - 0x1138  :    0 - 0x0
    "00000000", -- 4409 - 0x1139  :    0 - 0x0
    "00000000", -- 4410 - 0x113a  :    0 - 0x0
    "00000000", -- 4411 - 0x113b  :    0 - 0x0
    "00000000", -- 4412 - 0x113c  :    0 - 0x0
    "00000000", -- 4413 - 0x113d  :    0 - 0x0
    "00000000", -- 4414 - 0x113e  :    0 - 0x0
    "00000000", -- 4415 - 0x113f  :    0 - 0x0
    "00100100", -- 4416 - 0x1140  :   36 - 0x24 -- Background 0x14
    "00100100", -- 4417 - 0x1141  :   36 - 0x24
    "11000100", -- 4418 - 0x1142  :  196 - 0xc4
    "00000100", -- 4419 - 0x1143  :    4 - 0x4
    "00000100", -- 4420 - 0x1144  :    4 - 0x4
    "11000100", -- 4421 - 0x1145  :  196 - 0xc4
    "00100100", -- 4422 - 0x1146  :   36 - 0x24
    "00100100", -- 4423 - 0x1147  :   36 - 0x24
    "00000000", -- 4424 - 0x1148  :    0 - 0x0
    "00000000", -- 4425 - 0x1149  :    0 - 0x0
    "00000000", -- 4426 - 0x114a  :    0 - 0x0
    "00000000", -- 4427 - 0x114b  :    0 - 0x0
    "00000000", -- 4428 - 0x114c  :    0 - 0x0
    "00000000", -- 4429 - 0x114d  :    0 - 0x0
    "00000000", -- 4430 - 0x114e  :    0 - 0x0
    "00000000", -- 4431 - 0x114f  :    0 - 0x0
    "00100100", -- 4432 - 0x1150  :   36 - 0x24 -- Background 0x15
    "00100100", -- 4433 - 0x1151  :   36 - 0x24
    "00100011", -- 4434 - 0x1152  :   35 - 0x23
    "00100000", -- 4435 - 0x1153  :   32 - 0x20
    "00100000", -- 4436 - 0x1154  :   32 - 0x20
    "00100011", -- 4437 - 0x1155  :   35 - 0x23
    "00100100", -- 4438 - 0x1156  :   36 - 0x24
    "00100100", -- 4439 - 0x1157  :   36 - 0x24
    "00000000", -- 4440 - 0x1158  :    0 - 0x0
    "00000000", -- 4441 - 0x1159  :    0 - 0x0
    "00000000", -- 4442 - 0x115a  :    0 - 0x0
    "00000000", -- 4443 - 0x115b  :    0 - 0x0
    "00000000", -- 4444 - 0x115c  :    0 - 0x0
    "00000000", -- 4445 - 0x115d  :    0 - 0x0
    "00000000", -- 4446 - 0x115e  :    0 - 0x0
    "00000000", -- 4447 - 0x115f  :    0 - 0x0
    "00000000", -- 4448 - 0x1160  :    0 - 0x0 -- Background 0x16
    "00000000", -- 4449 - 0x1161  :    0 - 0x0
    "00001111", -- 4450 - 0x1162  :   15 - 0xf
    "00010000", -- 4451 - 0x1163  :   16 - 0x10
    "11110000", -- 4452 - 0x1164  :  240 - 0xf0
    "00001111", -- 4453 - 0x1165  :   15 - 0xf
    "00000000", -- 4454 - 0x1166  :    0 - 0x0
    "00000000", -- 4455 - 0x1167  :    0 - 0x0
    "00000000", -- 4456 - 0x1168  :    0 - 0x0
    "00000000", -- 4457 - 0x1169  :    0 - 0x0
    "00000000", -- 4458 - 0x116a  :    0 - 0x0
    "00000000", -- 4459 - 0x116b  :    0 - 0x0
    "00000000", -- 4460 - 0x116c  :    0 - 0x0
    "00000000", -- 4461 - 0x116d  :    0 - 0x0
    "00000000", -- 4462 - 0x116e  :    0 - 0x0
    "00000000", -- 4463 - 0x116f  :    0 - 0x0
    "00000000", -- 4464 - 0x1170  :    0 - 0x0 -- Background 0x17
    "00000000", -- 4465 - 0x1171  :    0 - 0x0
    "11110000", -- 4466 - 0x1172  :  240 - 0xf0
    "00001000", -- 4467 - 0x1173  :    8 - 0x8
    "00001111", -- 4468 - 0x1174  :   15 - 0xf
    "11110000", -- 4469 - 0x1175  :  240 - 0xf0
    "00000000", -- 4470 - 0x1176  :    0 - 0x0
    "00000000", -- 4471 - 0x1177  :    0 - 0x0
    "00000000", -- 4472 - 0x1178  :    0 - 0x0
    "00000000", -- 4473 - 0x1179  :    0 - 0x0
    "00000000", -- 4474 - 0x117a  :    0 - 0x0
    "00000000", -- 4475 - 0x117b  :    0 - 0x0
    "00000000", -- 4476 - 0x117c  :    0 - 0x0
    "00000000", -- 4477 - 0x117d  :    0 - 0x0
    "00000000", -- 4478 - 0x117e  :    0 - 0x0
    "00000000", -- 4479 - 0x117f  :    0 - 0x0
    "00000000", -- 4480 - 0x1180  :    0 - 0x0 -- Background 0x18
    "00000000", -- 4481 - 0x1181  :    0 - 0x0
    "11110000", -- 4482 - 0x1182  :  240 - 0xf0
    "00001000", -- 4483 - 0x1183  :    8 - 0x8
    "00001000", -- 4484 - 0x1184  :    8 - 0x8
    "11110000", -- 4485 - 0x1185  :  240 - 0xf0
    "00000000", -- 4486 - 0x1186  :    0 - 0x0
    "00000000", -- 4487 - 0x1187  :    0 - 0x0
    "00000000", -- 4488 - 0x1188  :    0 - 0x0
    "00000000", -- 4489 - 0x1189  :    0 - 0x0
    "00000000", -- 4490 - 0x118a  :    0 - 0x0
    "00000000", -- 4491 - 0x118b  :    0 - 0x0
    "00000000", -- 4492 - 0x118c  :    0 - 0x0
    "00000000", -- 4493 - 0x118d  :    0 - 0x0
    "00000000", -- 4494 - 0x118e  :    0 - 0x0
    "00000000", -- 4495 - 0x118f  :    0 - 0x0
    "00000000", -- 4496 - 0x1190  :    0 - 0x0 -- Background 0x19
    "00000000", -- 4497 - 0x1191  :    0 - 0x0
    "00001111", -- 4498 - 0x1192  :   15 - 0xf
    "00010000", -- 4499 - 0x1193  :   16 - 0x10
    "00010000", -- 4500 - 0x1194  :   16 - 0x10
    "00001111", -- 4501 - 0x1195  :   15 - 0xf
    "00000000", -- 4502 - 0x1196  :    0 - 0x0
    "00000000", -- 4503 - 0x1197  :    0 - 0x0
    "00000000", -- 4504 - 0x1198  :    0 - 0x0
    "00000000", -- 4505 - 0x1199  :    0 - 0x0
    "00000000", -- 4506 - 0x119a  :    0 - 0x0
    "00000000", -- 4507 - 0x119b  :    0 - 0x0
    "00000000", -- 4508 - 0x119c  :    0 - 0x0
    "00000000", -- 4509 - 0x119d  :    0 - 0x0
    "00000000", -- 4510 - 0x119e  :    0 - 0x0
    "00000000", -- 4511 - 0x119f  :    0 - 0x0
    "00100100", -- 4512 - 0x11a0  :   36 - 0x24 -- Background 0x1a
    "00100100", -- 4513 - 0x11a1  :   36 - 0x24
    "00100100", -- 4514 - 0x11a2  :   36 - 0x24
    "00100100", -- 4515 - 0x11a3  :   36 - 0x24
    "00011000", -- 4516 - 0x11a4  :   24 - 0x18
    "00000000", -- 4517 - 0x11a5  :    0 - 0x0
    "00000000", -- 4518 - 0x11a6  :    0 - 0x0
    "00000000", -- 4519 - 0x11a7  :    0 - 0x0
    "00000000", -- 4520 - 0x11a8  :    0 - 0x0
    "00000000", -- 4521 - 0x11a9  :    0 - 0x0
    "00000000", -- 4522 - 0x11aa  :    0 - 0x0
    "00000000", -- 4523 - 0x11ab  :    0 - 0x0
    "00000000", -- 4524 - 0x11ac  :    0 - 0x0
    "00000000", -- 4525 - 0x11ad  :    0 - 0x0
    "00000000", -- 4526 - 0x11ae  :    0 - 0x0
    "00000000", -- 4527 - 0x11af  :    0 - 0x0
    "00000000", -- 4528 - 0x11b0  :    0 - 0x0 -- Background 0x1b
    "00000000", -- 4529 - 0x11b1  :    0 - 0x0
    "00000000", -- 4530 - 0x11b2  :    0 - 0x0
    "00011000", -- 4531 - 0x11b3  :   24 - 0x18
    "00100100", -- 4532 - 0x11b4  :   36 - 0x24
    "00100100", -- 4533 - 0x11b5  :   36 - 0x24
    "00100100", -- 4534 - 0x11b6  :   36 - 0x24
    "00100100", -- 4535 - 0x11b7  :   36 - 0x24
    "00000000", -- 4536 - 0x11b8  :    0 - 0x0
    "00000000", -- 4537 - 0x11b9  :    0 - 0x0
    "00000000", -- 4538 - 0x11ba  :    0 - 0x0
    "00000000", -- 4539 - 0x11bb  :    0 - 0x0
    "00000000", -- 4540 - 0x11bc  :    0 - 0x0
    "00000000", -- 4541 - 0x11bd  :    0 - 0x0
    "00000000", -- 4542 - 0x11be  :    0 - 0x0
    "00000000", -- 4543 - 0x11bf  :    0 - 0x0
    "00100100", -- 4544 - 0x11c0  :   36 - 0x24 -- Background 0x1c
    "00100100", -- 4545 - 0x11c1  :   36 - 0x24
    "11000100", -- 4546 - 0x11c2  :  196 - 0xc4
    "00000100", -- 4547 - 0x11c3  :    4 - 0x4
    "00001000", -- 4548 - 0x11c4  :    8 - 0x8
    "11110000", -- 4549 - 0x11c5  :  240 - 0xf0
    "00000000", -- 4550 - 0x11c6  :    0 - 0x0
    "00000000", -- 4551 - 0x11c7  :    0 - 0x0
    "00000000", -- 4552 - 0x11c8  :    0 - 0x0
    "00000000", -- 4553 - 0x11c9  :    0 - 0x0
    "00000000", -- 4554 - 0x11ca  :    0 - 0x0
    "00000000", -- 4555 - 0x11cb  :    0 - 0x0
    "00000000", -- 4556 - 0x11cc  :    0 - 0x0
    "00000000", -- 4557 - 0x11cd  :    0 - 0x0
    "00000000", -- 4558 - 0x11ce  :    0 - 0x0
    "00000000", -- 4559 - 0x11cf  :    0 - 0x0
    "00000000", -- 4560 - 0x11d0  :    0 - 0x0 -- Background 0x1d
    "00000000", -- 4561 - 0x11d1  :    0 - 0x0
    "11110000", -- 4562 - 0x11d2  :  240 - 0xf0
    "00001000", -- 4563 - 0x11d3  :    8 - 0x8
    "00000100", -- 4564 - 0x11d4  :    4 - 0x4
    "11000100", -- 4565 - 0x11d5  :  196 - 0xc4
    "00100100", -- 4566 - 0x11d6  :   36 - 0x24
    "00100100", -- 4567 - 0x11d7  :   36 - 0x24
    "00000000", -- 4568 - 0x11d8  :    0 - 0x0
    "00000000", -- 4569 - 0x11d9  :    0 - 0x0
    "00000000", -- 4570 - 0x11da  :    0 - 0x0
    "00000000", -- 4571 - 0x11db  :    0 - 0x0
    "00000000", -- 4572 - 0x11dc  :    0 - 0x0
    "00000000", -- 4573 - 0x11dd  :    0 - 0x0
    "00000000", -- 4574 - 0x11de  :    0 - 0x0
    "00000000", -- 4575 - 0x11df  :    0 - 0x0
    "00100100", -- 4576 - 0x11e0  :   36 - 0x24 -- Background 0x1e
    "00100100", -- 4577 - 0x11e1  :   36 - 0x24
    "00100011", -- 4578 - 0x11e2  :   35 - 0x23
    "00100000", -- 4579 - 0x11e3  :   32 - 0x20
    "00010000", -- 4580 - 0x11e4  :   16 - 0x10
    "00001111", -- 4581 - 0x11e5  :   15 - 0xf
    "00000000", -- 4582 - 0x11e6  :    0 - 0x0
    "00000000", -- 4583 - 0x11e7  :    0 - 0x0
    "00000000", -- 4584 - 0x11e8  :    0 - 0x0
    "00000000", -- 4585 - 0x11e9  :    0 - 0x0
    "00000000", -- 4586 - 0x11ea  :    0 - 0x0
    "00000000", -- 4587 - 0x11eb  :    0 - 0x0
    "00000000", -- 4588 - 0x11ec  :    0 - 0x0
    "00000000", -- 4589 - 0x11ed  :    0 - 0x0
    "00000000", -- 4590 - 0x11ee  :    0 - 0x0
    "00000000", -- 4591 - 0x11ef  :    0 - 0x0
    "00000000", -- 4592 - 0x11f0  :    0 - 0x0 -- Background 0x1f
    "00000000", -- 4593 - 0x11f1  :    0 - 0x0
    "00001111", -- 4594 - 0x11f2  :   15 - 0xf
    "00010000", -- 4595 - 0x11f3  :   16 - 0x10
    "00100000", -- 4596 - 0x11f4  :   32 - 0x20
    "00100011", -- 4597 - 0x11f5  :   35 - 0x23
    "00100100", -- 4598 - 0x11f6  :   36 - 0x24
    "00100100", -- 4599 - 0x11f7  :   36 - 0x24
    "00000000", -- 4600 - 0x11f8  :    0 - 0x0
    "00000000", -- 4601 - 0x11f9  :    0 - 0x0
    "00000000", -- 4602 - 0x11fa  :    0 - 0x0
    "00000000", -- 4603 - 0x11fb  :    0 - 0x0
    "00000000", -- 4604 - 0x11fc  :    0 - 0x0
    "00000000", -- 4605 - 0x11fd  :    0 - 0x0
    "00000000", -- 4606 - 0x11fe  :    0 - 0x0
    "00000000", -- 4607 - 0x11ff  :    0 - 0x0
    "00000000", -- 4608 - 0x1200  :    0 - 0x0 -- Background 0x20
    "00000000", -- 4609 - 0x1201  :    0 - 0x0
    "00000000", -- 4610 - 0x1202  :    0 - 0x0
    "00000000", -- 4611 - 0x1203  :    0 - 0x0
    "00000000", -- 4612 - 0x1204  :    0 - 0x0
    "00000000", -- 4613 - 0x1205  :    0 - 0x0
    "00000000", -- 4614 - 0x1206  :    0 - 0x0
    "00000000", -- 4615 - 0x1207  :    0 - 0x0
    "00000000", -- 4616 - 0x1208  :    0 - 0x0
    "00000000", -- 4617 - 0x1209  :    0 - 0x0
    "00000000", -- 4618 - 0x120a  :    0 - 0x0
    "00000000", -- 4619 - 0x120b  :    0 - 0x0
    "00000000", -- 4620 - 0x120c  :    0 - 0x0
    "00000000", -- 4621 - 0x120d  :    0 - 0x0
    "00000000", -- 4622 - 0x120e  :    0 - 0x0
    "00000000", -- 4623 - 0x120f  :    0 - 0x0
    "00000000", -- 4624 - 0x1210  :    0 - 0x0 -- Background 0x21
    "00000000", -- 4625 - 0x1211  :    0 - 0x0
    "11110000", -- 4626 - 0x1212  :  240 - 0xf0
    "00001000", -- 4627 - 0x1213  :    8 - 0x8
    "00001000", -- 4628 - 0x1214  :    8 - 0x8
    "11110000", -- 4629 - 0x1215  :  240 - 0xf0
    "00000000", -- 4630 - 0x1216  :    0 - 0x0
    "00000000", -- 4631 - 0x1217  :    0 - 0x0
    "00001111", -- 4632 - 0x1218  :   15 - 0xf
    "00001111", -- 4633 - 0x1219  :   15 - 0xf
    "00001111", -- 4634 - 0x121a  :   15 - 0xf
    "00000111", -- 4635 - 0x121b  :    7 - 0x7
    "00000111", -- 4636 - 0x121c  :    7 - 0x7
    "00001111", -- 4637 - 0x121d  :   15 - 0xf
    "00001111", -- 4638 - 0x121e  :   15 - 0xf
    "00001111", -- 4639 - 0x121f  :   15 - 0xf
    "00000000", -- 4640 - 0x1220  :    0 - 0x0 -- Background 0x22
    "00000000", -- 4641 - 0x1221  :    0 - 0x0
    "00001111", -- 4642 - 0x1222  :   15 - 0xf
    "00010000", -- 4643 - 0x1223  :   16 - 0x10
    "00010000", -- 4644 - 0x1224  :   16 - 0x10
    "00001111", -- 4645 - 0x1225  :   15 - 0xf
    "00000000", -- 4646 - 0x1226  :    0 - 0x0
    "00000000", -- 4647 - 0x1227  :    0 - 0x0
    "11110000", -- 4648 - 0x1228  :  240 - 0xf0
    "11110000", -- 4649 - 0x1229  :  240 - 0xf0
    "11110000", -- 4650 - 0x122a  :  240 - 0xf0
    "11100000", -- 4651 - 0x122b  :  224 - 0xe0
    "11100000", -- 4652 - 0x122c  :  224 - 0xe0
    "11110000", -- 4653 - 0x122d  :  240 - 0xf0
    "11110000", -- 4654 - 0x122e  :  240 - 0xf0
    "11110000", -- 4655 - 0x122f  :  240 - 0xf0
    "11111111", -- 4656 - 0x1230  :  255 - 0xff -- Background 0x23
    "11111111", -- 4657 - 0x1231  :  255 - 0xff
    "11100001", -- 4658 - 0x1232  :  225 - 0xe1
    "11100001", -- 4659 - 0x1233  :  225 - 0xe1
    "11100001", -- 4660 - 0x1234  :  225 - 0xe1
    "11100001", -- 4661 - 0x1235  :  225 - 0xe1
    "11100001", -- 4662 - 0x1236  :  225 - 0xe1
    "11100001", -- 4663 - 0x1237  :  225 - 0xe1
    "11111111", -- 4664 - 0x1238  :  255 - 0xff
    "11111111", -- 4665 - 0x1239  :  255 - 0xff
    "11100001", -- 4666 - 0x123a  :  225 - 0xe1
    "11100001", -- 4667 - 0x123b  :  225 - 0xe1
    "11100001", -- 4668 - 0x123c  :  225 - 0xe1
    "11100001", -- 4669 - 0x123d  :  225 - 0xe1
    "11100001", -- 4670 - 0x123e  :  225 - 0xe1
    "11100001", -- 4671 - 0x123f  :  225 - 0xe1
    "10000111", -- 4672 - 0x1240  :  135 - 0x87 -- Background 0x24
    "11000111", -- 4673 - 0x1241  :  199 - 0xc7
    "11000000", -- 4674 - 0x1242  :  192 - 0xc0
    "11000111", -- 4675 - 0x1243  :  199 - 0xc7
    "11001111", -- 4676 - 0x1244  :  207 - 0xcf
    "11001110", -- 4677 - 0x1245  :  206 - 0xce
    "11001111", -- 4678 - 0x1246  :  207 - 0xcf
    "11000111", -- 4679 - 0x1247  :  199 - 0xc7
    "10000111", -- 4680 - 0x1248  :  135 - 0x87
    "11000111", -- 4681 - 0x1249  :  199 - 0xc7
    "11000000", -- 4682 - 0x124a  :  192 - 0xc0
    "11000111", -- 4683 - 0x124b  :  199 - 0xc7
    "11001111", -- 4684 - 0x124c  :  207 - 0xcf
    "11001110", -- 4685 - 0x124d  :  206 - 0xce
    "11001111", -- 4686 - 0x124e  :  207 - 0xcf
    "11000111", -- 4687 - 0x124f  :  199 - 0xc7
    "11111000", -- 4688 - 0x1250  :  248 - 0xf8 -- Background 0x25
    "11111100", -- 4689 - 0x1251  :  252 - 0xfc
    "00011100", -- 4690 - 0x1252  :   28 - 0x1c
    "11111100", -- 4691 - 0x1253  :  252 - 0xfc
    "11111100", -- 4692 - 0x1254  :  252 - 0xfc
    "00011100", -- 4693 - 0x1255  :   28 - 0x1c
    "11111100", -- 4694 - 0x1256  :  252 - 0xfc
    "11111100", -- 4695 - 0x1257  :  252 - 0xfc
    "11111000", -- 4696 - 0x1258  :  248 - 0xf8
    "11111100", -- 4697 - 0x1259  :  252 - 0xfc
    "00011100", -- 4698 - 0x125a  :   28 - 0x1c
    "11111100", -- 4699 - 0x125b  :  252 - 0xfc
    "11111100", -- 4700 - 0x125c  :  252 - 0xfc
    "00011100", -- 4701 - 0x125d  :   28 - 0x1c
    "11111100", -- 4702 - 0x125e  :  252 - 0xfc
    "11111100", -- 4703 - 0x125f  :  252 - 0xfc
    "11111111", -- 4704 - 0x1260  :  255 - 0xff -- Background 0x26
    "11111111", -- 4705 - 0x1261  :  255 - 0xff
    "11100111", -- 4706 - 0x1262  :  231 - 0xe7
    "11100111", -- 4707 - 0x1263  :  231 - 0xe7
    "11100111", -- 4708 - 0x1264  :  231 - 0xe7
    "11100111", -- 4709 - 0x1265  :  231 - 0xe7
    "11100111", -- 4710 - 0x1266  :  231 - 0xe7
    "11100111", -- 4711 - 0x1267  :  231 - 0xe7
    "11111111", -- 4712 - 0x1268  :  255 - 0xff
    "11111111", -- 4713 - 0x1269  :  255 - 0xff
    "11100111", -- 4714 - 0x126a  :  231 - 0xe7
    "11100111", -- 4715 - 0x126b  :  231 - 0xe7
    "11100111", -- 4716 - 0x126c  :  231 - 0xe7
    "11100111", -- 4717 - 0x126d  :  231 - 0xe7
    "11100111", -- 4718 - 0x126e  :  231 - 0xe7
    "11100111", -- 4719 - 0x126f  :  231 - 0xe7
    "11110000", -- 4720 - 0x1270  :  240 - 0xf0 -- Background 0x27
    "11111001", -- 4721 - 0x1271  :  249 - 0xf9
    "00111001", -- 4722 - 0x1272  :   57 - 0x39
    "00111001", -- 4723 - 0x1273  :   57 - 0x39
    "00111001", -- 4724 - 0x1274  :   57 - 0x39
    "00111001", -- 4725 - 0x1275  :   57 - 0x39
    "00111001", -- 4726 - 0x1276  :   57 - 0x39
    "00111000", -- 4727 - 0x1277  :   56 - 0x38
    "11110000", -- 4728 - 0x1278  :  240 - 0xf0
    "11111001", -- 4729 - 0x1279  :  249 - 0xf9
    "00111001", -- 4730 - 0x127a  :   57 - 0x39
    "00111001", -- 4731 - 0x127b  :   57 - 0x39
    "00111001", -- 4732 - 0x127c  :   57 - 0x39
    "00111001", -- 4733 - 0x127d  :   57 - 0x39
    "00111001", -- 4734 - 0x127e  :   57 - 0x39
    "00111000", -- 4735 - 0x127f  :   56 - 0x38
    "11111111", -- 4736 - 0x1280  :  255 - 0xff -- Background 0x28
    "11111111", -- 4737 - 0x1281  :  255 - 0xff
    "11000000", -- 4738 - 0x1282  :  192 - 0xc0
    "11000000", -- 4739 - 0x1283  :  192 - 0xc0
    "11000000", -- 4740 - 0x1284  :  192 - 0xc0
    "11000000", -- 4741 - 0x1285  :  192 - 0xc0
    "11111111", -- 4742 - 0x1286  :  255 - 0xff
    "11111111", -- 4743 - 0x1287  :  255 - 0xff
    "11111111", -- 4744 - 0x1288  :  255 - 0xff
    "11111111", -- 4745 - 0x1289  :  255 - 0xff
    "11000000", -- 4746 - 0x128a  :  192 - 0xc0
    "11000000", -- 4747 - 0x128b  :  192 - 0xc0
    "11000000", -- 4748 - 0x128c  :  192 - 0xc0
    "11000000", -- 4749 - 0x128d  :  192 - 0xc0
    "11111111", -- 4750 - 0x128e  :  255 - 0xff
    "11111111", -- 4751 - 0x128f  :  255 - 0xff
    "00011111", -- 4752 - 0x1290  :   31 - 0x1f -- Background 0x29
    "00111111", -- 4753 - 0x1291  :   63 - 0x3f
    "00110000", -- 4754 - 0x1292  :   48 - 0x30
    "00110000", -- 4755 - 0x1293  :   48 - 0x30
    "00110000", -- 4756 - 0x1294  :   48 - 0x30
    "00110000", -- 4757 - 0x1295  :   48 - 0x30
    "00111111", -- 4758 - 0x1296  :   63 - 0x3f
    "00011111", -- 4759 - 0x1297  :   31 - 0x1f
    "00011111", -- 4760 - 0x1298  :   31 - 0x1f
    "00111111", -- 4761 - 0x1299  :   63 - 0x3f
    "00110000", -- 4762 - 0x129a  :   48 - 0x30
    "00110000", -- 4763 - 0x129b  :   48 - 0x30
    "00110000", -- 4764 - 0x129c  :   48 - 0x30
    "00110000", -- 4765 - 0x129d  :   48 - 0x30
    "00111111", -- 4766 - 0x129e  :   63 - 0x3f
    "00011111", -- 4767 - 0x129f  :   31 - 0x1f
    "11100011", -- 4768 - 0x12a0  :  227 - 0xe3 -- Background 0x2a
    "11110011", -- 4769 - 0x12a1  :  243 - 0xf3
    "01110000", -- 4770 - 0x12a2  :  112 - 0x70
    "01110000", -- 4771 - 0x12a3  :  112 - 0x70
    "01110000", -- 4772 - 0x12a4  :  112 - 0x70
    "01110000", -- 4773 - 0x12a5  :  112 - 0x70
    "11110000", -- 4774 - 0x12a6  :  240 - 0xf0
    "11100000", -- 4775 - 0x12a7  :  224 - 0xe0
    "11100011", -- 4776 - 0x12a8  :  227 - 0xe3
    "11110011", -- 4777 - 0x12a9  :  243 - 0xf3
    "01110000", -- 4778 - 0x12aa  :  112 - 0x70
    "01110000", -- 4779 - 0x12ab  :  112 - 0x70
    "01110000", -- 4780 - 0x12ac  :  112 - 0x70
    "01110000", -- 4781 - 0x12ad  :  112 - 0x70
    "11110000", -- 4782 - 0x12ae  :  240 - 0xf0
    "11100000", -- 4783 - 0x12af  :  224 - 0xe0
    "11111110", -- 4784 - 0x12b0  :  254 - 0xfe -- Background 0x2b
    "11111110", -- 4785 - 0x12b1  :  254 - 0xfe
    "01110000", -- 4786 - 0x12b2  :  112 - 0x70
    "01110000", -- 4787 - 0x12b3  :  112 - 0x70
    "01110000", -- 4788 - 0x12b4  :  112 - 0x70
    "01110000", -- 4789 - 0x12b5  :  112 - 0x70
    "01110000", -- 4790 - 0x12b6  :  112 - 0x70
    "01110000", -- 4791 - 0x12b7  :  112 - 0x70
    "11111110", -- 4792 - 0x12b8  :  254 - 0xfe
    "11111110", -- 4793 - 0x12b9  :  254 - 0xfe
    "01110000", -- 4794 - 0x12ba  :  112 - 0x70
    "01110000", -- 4795 - 0x12bb  :  112 - 0x70
    "01110000", -- 4796 - 0x12bc  :  112 - 0x70
    "01110000", -- 4797 - 0x12bd  :  112 - 0x70
    "01110000", -- 4798 - 0x12be  :  112 - 0x70
    "01110000", -- 4799 - 0x12bf  :  112 - 0x70
    "00000000", -- 4800 - 0x12c0  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 4801 - 0x12c1  :    0 - 0x0
    "00000000", -- 4802 - 0x12c2  :    0 - 0x0
    "00000000", -- 4803 - 0x12c3  :    0 - 0x0
    "11111111", -- 4804 - 0x12c4  :  255 - 0xff
    "00000000", -- 4805 - 0x12c5  :    0 - 0x0
    "00000000", -- 4806 - 0x12c6  :    0 - 0x0
    "00000000", -- 4807 - 0x12c7  :    0 - 0x0
    "00000000", -- 4808 - 0x12c8  :    0 - 0x0
    "00000000", -- 4809 - 0x12c9  :    0 - 0x0
    "00000000", -- 4810 - 0x12ca  :    0 - 0x0
    "00000000", -- 4811 - 0x12cb  :    0 - 0x0
    "00000000", -- 4812 - 0x12cc  :    0 - 0x0
    "00000000", -- 4813 - 0x12cd  :    0 - 0x0
    "00000000", -- 4814 - 0x12ce  :    0 - 0x0
    "00000000", -- 4815 - 0x12cf  :    0 - 0x0
    "00000000", -- 4816 - 0x12d0  :    0 - 0x0 -- Background 0x2d
    "00000000", -- 4817 - 0x12d1  :    0 - 0x0
    "00000000", -- 4818 - 0x12d2  :    0 - 0x0
    "00000000", -- 4819 - 0x12d3  :    0 - 0x0
    "00000000", -- 4820 - 0x12d4  :    0 - 0x0
    "00000000", -- 4821 - 0x12d5  :    0 - 0x0
    "00000000", -- 4822 - 0x12d6  :    0 - 0x0
    "00000000", -- 4823 - 0x12d7  :    0 - 0x0
    "11111111", -- 4824 - 0x12d8  :  255 - 0xff
    "11111111", -- 4825 - 0x12d9  :  255 - 0xff
    "11111111", -- 4826 - 0x12da  :  255 - 0xff
    "11111111", -- 4827 - 0x12db  :  255 - 0xff
    "11111111", -- 4828 - 0x12dc  :  255 - 0xff
    "11111111", -- 4829 - 0x12dd  :  255 - 0xff
    "11111111", -- 4830 - 0x12de  :  255 - 0xff
    "11111111", -- 4831 - 0x12df  :  255 - 0xff
    "00000000", -- 4832 - 0x12e0  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 4833 - 0x12e1  :    0 - 0x0
    "00000000", -- 4834 - 0x12e2  :    0 - 0x0
    "00011000", -- 4835 - 0x12e3  :   24 - 0x18
    "00011000", -- 4836 - 0x12e4  :   24 - 0x18
    "00000000", -- 4837 - 0x12e5  :    0 - 0x0
    "00000000", -- 4838 - 0x12e6  :    0 - 0x0
    "00000000", -- 4839 - 0x12e7  :    0 - 0x0
    "00000000", -- 4840 - 0x12e8  :    0 - 0x0
    "00000000", -- 4841 - 0x12e9  :    0 - 0x0
    "00000000", -- 4842 - 0x12ea  :    0 - 0x0
    "00000000", -- 4843 - 0x12eb  :    0 - 0x0
    "00000000", -- 4844 - 0x12ec  :    0 - 0x0
    "00000000", -- 4845 - 0x12ed  :    0 - 0x0
    "00000000", -- 4846 - 0x12ee  :    0 - 0x0
    "00000000", -- 4847 - 0x12ef  :    0 - 0x0
    "00000000", -- 4848 - 0x12f0  :    0 - 0x0 -- Background 0x2f
    "00000000", -- 4849 - 0x12f1  :    0 - 0x0
    "00000000", -- 4850 - 0x12f2  :    0 - 0x0
    "00000000", -- 4851 - 0x12f3  :    0 - 0x0
    "00000000", -- 4852 - 0x12f4  :    0 - 0x0
    "00000000", -- 4853 - 0x12f5  :    0 - 0x0
    "00000000", -- 4854 - 0x12f6  :    0 - 0x0
    "00000000", -- 4855 - 0x12f7  :    0 - 0x0
    "00000000", -- 4856 - 0x12f8  :    0 - 0x0
    "00000000", -- 4857 - 0x12f9  :    0 - 0x0
    "00000000", -- 4858 - 0x12fa  :    0 - 0x0
    "00011000", -- 4859 - 0x12fb  :   24 - 0x18
    "00011000", -- 4860 - 0x12fc  :   24 - 0x18
    "00000000", -- 4861 - 0x12fd  :    0 - 0x0
    "00000000", -- 4862 - 0x12fe  :    0 - 0x0
    "00000000", -- 4863 - 0x12ff  :    0 - 0x0
    "00011100", -- 4864 - 0x1300  :   28 - 0x1c -- Background 0x30
    "00100110", -- 4865 - 0x1301  :   38 - 0x26
    "01100011", -- 4866 - 0x1302  :   99 - 0x63
    "01100011", -- 4867 - 0x1303  :   99 - 0x63
    "01100011", -- 4868 - 0x1304  :   99 - 0x63
    "00110010", -- 4869 - 0x1305  :   50 - 0x32
    "00011100", -- 4870 - 0x1306  :   28 - 0x1c
    "00000000", -- 4871 - 0x1307  :    0 - 0x0
    "00000000", -- 4872 - 0x1308  :    0 - 0x0
    "00000000", -- 4873 - 0x1309  :    0 - 0x0
    "00000000", -- 4874 - 0x130a  :    0 - 0x0
    "00000000", -- 4875 - 0x130b  :    0 - 0x0
    "00000000", -- 4876 - 0x130c  :    0 - 0x0
    "00000000", -- 4877 - 0x130d  :    0 - 0x0
    "00000000", -- 4878 - 0x130e  :    0 - 0x0
    "00000000", -- 4879 - 0x130f  :    0 - 0x0
    "00001100", -- 4880 - 0x1310  :   12 - 0xc -- Background 0x31
    "00011100", -- 4881 - 0x1311  :   28 - 0x1c
    "00001100", -- 4882 - 0x1312  :   12 - 0xc
    "00001100", -- 4883 - 0x1313  :   12 - 0xc
    "00001100", -- 4884 - 0x1314  :   12 - 0xc
    "00001100", -- 4885 - 0x1315  :   12 - 0xc
    "00111111", -- 4886 - 0x1316  :   63 - 0x3f
    "00000000", -- 4887 - 0x1317  :    0 - 0x0
    "00000000", -- 4888 - 0x1318  :    0 - 0x0
    "00000000", -- 4889 - 0x1319  :    0 - 0x0
    "00000000", -- 4890 - 0x131a  :    0 - 0x0
    "00000000", -- 4891 - 0x131b  :    0 - 0x0
    "00000000", -- 4892 - 0x131c  :    0 - 0x0
    "00000000", -- 4893 - 0x131d  :    0 - 0x0
    "00000000", -- 4894 - 0x131e  :    0 - 0x0
    "00000000", -- 4895 - 0x131f  :    0 - 0x0
    "00111110", -- 4896 - 0x1320  :   62 - 0x3e -- Background 0x32
    "01100011", -- 4897 - 0x1321  :   99 - 0x63
    "00000111", -- 4898 - 0x1322  :    7 - 0x7
    "00011110", -- 4899 - 0x1323  :   30 - 0x1e
    "00111100", -- 4900 - 0x1324  :   60 - 0x3c
    "01110000", -- 4901 - 0x1325  :  112 - 0x70
    "01111111", -- 4902 - 0x1326  :  127 - 0x7f
    "00000000", -- 4903 - 0x1327  :    0 - 0x0
    "00000000", -- 4904 - 0x1328  :    0 - 0x0
    "00000000", -- 4905 - 0x1329  :    0 - 0x0
    "00000000", -- 4906 - 0x132a  :    0 - 0x0
    "00000000", -- 4907 - 0x132b  :    0 - 0x0
    "00000000", -- 4908 - 0x132c  :    0 - 0x0
    "00000000", -- 4909 - 0x132d  :    0 - 0x0
    "00000000", -- 4910 - 0x132e  :    0 - 0x0
    "00000000", -- 4911 - 0x132f  :    0 - 0x0
    "00111111", -- 4912 - 0x1330  :   63 - 0x3f -- Background 0x33
    "00000110", -- 4913 - 0x1331  :    6 - 0x6
    "00001100", -- 4914 - 0x1332  :   12 - 0xc
    "00011110", -- 4915 - 0x1333  :   30 - 0x1e
    "00000011", -- 4916 - 0x1334  :    3 - 0x3
    "01100011", -- 4917 - 0x1335  :   99 - 0x63
    "00111110", -- 4918 - 0x1336  :   62 - 0x3e
    "00000000", -- 4919 - 0x1337  :    0 - 0x0
    "00000000", -- 4920 - 0x1338  :    0 - 0x0
    "00000000", -- 4921 - 0x1339  :    0 - 0x0
    "00000000", -- 4922 - 0x133a  :    0 - 0x0
    "00000000", -- 4923 - 0x133b  :    0 - 0x0
    "00000000", -- 4924 - 0x133c  :    0 - 0x0
    "00000000", -- 4925 - 0x133d  :    0 - 0x0
    "00000000", -- 4926 - 0x133e  :    0 - 0x0
    "00000000", -- 4927 - 0x133f  :    0 - 0x0
    "00001110", -- 4928 - 0x1340  :   14 - 0xe -- Background 0x34
    "00011110", -- 4929 - 0x1341  :   30 - 0x1e
    "00110110", -- 4930 - 0x1342  :   54 - 0x36
    "01100110", -- 4931 - 0x1343  :  102 - 0x66
    "01111111", -- 4932 - 0x1344  :  127 - 0x7f
    "00000110", -- 4933 - 0x1345  :    6 - 0x6
    "00000110", -- 4934 - 0x1346  :    6 - 0x6
    "00000000", -- 4935 - 0x1347  :    0 - 0x0
    "00000000", -- 4936 - 0x1348  :    0 - 0x0
    "00000000", -- 4937 - 0x1349  :    0 - 0x0
    "00000000", -- 4938 - 0x134a  :    0 - 0x0
    "00000000", -- 4939 - 0x134b  :    0 - 0x0
    "00000000", -- 4940 - 0x134c  :    0 - 0x0
    "00000000", -- 4941 - 0x134d  :    0 - 0x0
    "00000000", -- 4942 - 0x134e  :    0 - 0x0
    "00000000", -- 4943 - 0x134f  :    0 - 0x0
    "01111110", -- 4944 - 0x1350  :  126 - 0x7e -- Background 0x35
    "01100000", -- 4945 - 0x1351  :   96 - 0x60
    "01111110", -- 4946 - 0x1352  :  126 - 0x7e
    "00000011", -- 4947 - 0x1353  :    3 - 0x3
    "00000011", -- 4948 - 0x1354  :    3 - 0x3
    "01100011", -- 4949 - 0x1355  :   99 - 0x63
    "00111110", -- 4950 - 0x1356  :   62 - 0x3e
    "00000000", -- 4951 - 0x1357  :    0 - 0x0
    "00000000", -- 4952 - 0x1358  :    0 - 0x0
    "00000000", -- 4953 - 0x1359  :    0 - 0x0
    "00000000", -- 4954 - 0x135a  :    0 - 0x0
    "00000000", -- 4955 - 0x135b  :    0 - 0x0
    "00000000", -- 4956 - 0x135c  :    0 - 0x0
    "00000000", -- 4957 - 0x135d  :    0 - 0x0
    "00000000", -- 4958 - 0x135e  :    0 - 0x0
    "00000000", -- 4959 - 0x135f  :    0 - 0x0
    "00011110", -- 4960 - 0x1360  :   30 - 0x1e -- Background 0x36
    "00110000", -- 4961 - 0x1361  :   48 - 0x30
    "01100000", -- 4962 - 0x1362  :   96 - 0x60
    "01111110", -- 4963 - 0x1363  :  126 - 0x7e
    "01100011", -- 4964 - 0x1364  :   99 - 0x63
    "01100011", -- 4965 - 0x1365  :   99 - 0x63
    "00111110", -- 4966 - 0x1366  :   62 - 0x3e
    "00000000", -- 4967 - 0x1367  :    0 - 0x0
    "00000000", -- 4968 - 0x1368  :    0 - 0x0
    "00000000", -- 4969 - 0x1369  :    0 - 0x0
    "00000000", -- 4970 - 0x136a  :    0 - 0x0
    "00000000", -- 4971 - 0x136b  :    0 - 0x0
    "00000000", -- 4972 - 0x136c  :    0 - 0x0
    "00000000", -- 4973 - 0x136d  :    0 - 0x0
    "00000000", -- 4974 - 0x136e  :    0 - 0x0
    "00000000", -- 4975 - 0x136f  :    0 - 0x0
    "01111111", -- 4976 - 0x1370  :  127 - 0x7f -- Background 0x37
    "01100011", -- 4977 - 0x1371  :   99 - 0x63
    "00000110", -- 4978 - 0x1372  :    6 - 0x6
    "00001100", -- 4979 - 0x1373  :   12 - 0xc
    "00011000", -- 4980 - 0x1374  :   24 - 0x18
    "00011000", -- 4981 - 0x1375  :   24 - 0x18
    "00011000", -- 4982 - 0x1376  :   24 - 0x18
    "00000000", -- 4983 - 0x1377  :    0 - 0x0
    "00000000", -- 4984 - 0x1378  :    0 - 0x0
    "00000000", -- 4985 - 0x1379  :    0 - 0x0
    "00000000", -- 4986 - 0x137a  :    0 - 0x0
    "00000000", -- 4987 - 0x137b  :    0 - 0x0
    "00000000", -- 4988 - 0x137c  :    0 - 0x0
    "00000000", -- 4989 - 0x137d  :    0 - 0x0
    "00000000", -- 4990 - 0x137e  :    0 - 0x0
    "00000000", -- 4991 - 0x137f  :    0 - 0x0
    "00111100", -- 4992 - 0x1380  :   60 - 0x3c -- Background 0x38
    "01100010", -- 4993 - 0x1381  :   98 - 0x62
    "01110010", -- 4994 - 0x1382  :  114 - 0x72
    "00111100", -- 4995 - 0x1383  :   60 - 0x3c
    "01001111", -- 4996 - 0x1384  :   79 - 0x4f
    "01000011", -- 4997 - 0x1385  :   67 - 0x43
    "00111110", -- 4998 - 0x1386  :   62 - 0x3e
    "00000000", -- 4999 - 0x1387  :    0 - 0x0
    "00000000", -- 5000 - 0x1388  :    0 - 0x0
    "00000000", -- 5001 - 0x1389  :    0 - 0x0
    "00000000", -- 5002 - 0x138a  :    0 - 0x0
    "00000000", -- 5003 - 0x138b  :    0 - 0x0
    "00000000", -- 5004 - 0x138c  :    0 - 0x0
    "00000000", -- 5005 - 0x138d  :    0 - 0x0
    "00000000", -- 5006 - 0x138e  :    0 - 0x0
    "00000000", -- 5007 - 0x138f  :    0 - 0x0
    "00111110", -- 5008 - 0x1390  :   62 - 0x3e -- Background 0x39
    "01100011", -- 5009 - 0x1391  :   99 - 0x63
    "01100011", -- 5010 - 0x1392  :   99 - 0x63
    "00111111", -- 5011 - 0x1393  :   63 - 0x3f
    "00000011", -- 5012 - 0x1394  :    3 - 0x3
    "00000110", -- 5013 - 0x1395  :    6 - 0x6
    "00111100", -- 5014 - 0x1396  :   60 - 0x3c
    "00000000", -- 5015 - 0x1397  :    0 - 0x0
    "00000000", -- 5016 - 0x1398  :    0 - 0x0
    "00000000", -- 5017 - 0x1399  :    0 - 0x0
    "00000000", -- 5018 - 0x139a  :    0 - 0x0
    "00000000", -- 5019 - 0x139b  :    0 - 0x0
    "00000000", -- 5020 - 0x139c  :    0 - 0x0
    "00000000", -- 5021 - 0x139d  :    0 - 0x0
    "00000000", -- 5022 - 0x139e  :    0 - 0x0
    "00000000", -- 5023 - 0x139f  :    0 - 0x0
    "00000000", -- 5024 - 0x13a0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 5025 - 0x13a1  :    0 - 0x0
    "00000000", -- 5026 - 0x13a2  :    0 - 0x0
    "01111110", -- 5027 - 0x13a3  :  126 - 0x7e
    "00000000", -- 5028 - 0x13a4  :    0 - 0x0
    "00000000", -- 5029 - 0x13a5  :    0 - 0x0
    "00000000", -- 5030 - 0x13a6  :    0 - 0x0
    "00000000", -- 5031 - 0x13a7  :    0 - 0x0
    "00000000", -- 5032 - 0x13a8  :    0 - 0x0
    "00000000", -- 5033 - 0x13a9  :    0 - 0x0
    "00000000", -- 5034 - 0x13aa  :    0 - 0x0
    "00000000", -- 5035 - 0x13ab  :    0 - 0x0
    "00000000", -- 5036 - 0x13ac  :    0 - 0x0
    "00000000", -- 5037 - 0x13ad  :    0 - 0x0
    "00000000", -- 5038 - 0x13ae  :    0 - 0x0
    "00000000", -- 5039 - 0x13af  :    0 - 0x0
    "00000000", -- 5040 - 0x13b0  :    0 - 0x0 -- Background 0x3b
    "00000010", -- 5041 - 0x13b1  :    2 - 0x2
    "00000100", -- 5042 - 0x13b2  :    4 - 0x4
    "00001000", -- 5043 - 0x13b3  :    8 - 0x8
    "00010000", -- 5044 - 0x13b4  :   16 - 0x10
    "00100000", -- 5045 - 0x13b5  :   32 - 0x20
    "00000000", -- 5046 - 0x13b6  :    0 - 0x0
    "00000000", -- 5047 - 0x13b7  :    0 - 0x0
    "00000000", -- 5048 - 0x13b8  :    0 - 0x0
    "00000000", -- 5049 - 0x13b9  :    0 - 0x0
    "00000000", -- 5050 - 0x13ba  :    0 - 0x0
    "00000000", -- 5051 - 0x13bb  :    0 - 0x0
    "00000000", -- 5052 - 0x13bc  :    0 - 0x0
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "00000000", -- 5054 - 0x13be  :    0 - 0x0
    "00000000", -- 5055 - 0x13bf  :    0 - 0x0
    "00000000", -- 5056 - 0x13c0  :    0 - 0x0 -- Background 0x3c
    "00000111", -- 5057 - 0x13c1  :    7 - 0x7
    "00011111", -- 5058 - 0x13c2  :   31 - 0x1f
    "00111111", -- 5059 - 0x13c3  :   63 - 0x3f
    "00111111", -- 5060 - 0x13c4  :   63 - 0x3f
    "00001111", -- 5061 - 0x13c5  :   15 - 0xf
    "00000011", -- 5062 - 0x13c6  :    3 - 0x3
    "00000000", -- 5063 - 0x13c7  :    0 - 0x0
    "00000000", -- 5064 - 0x13c8  :    0 - 0x0
    "00000111", -- 5065 - 0x13c9  :    7 - 0x7
    "00011111", -- 5066 - 0x13ca  :   31 - 0x1f
    "00111111", -- 5067 - 0x13cb  :   63 - 0x3f
    "00111111", -- 5068 - 0x13cc  :   63 - 0x3f
    "00001111", -- 5069 - 0x13cd  :   15 - 0xf
    "00000011", -- 5070 - 0x13ce  :    3 - 0x3
    "00000000", -- 5071 - 0x13cf  :    0 - 0x0
    "00000000", -- 5072 - 0x13d0  :    0 - 0x0 -- Background 0x3d
    "11000000", -- 5073 - 0x13d1  :  192 - 0xc0
    "11110000", -- 5074 - 0x13d2  :  240 - 0xf0
    "11111000", -- 5075 - 0x13d3  :  248 - 0xf8
    "11111000", -- 5076 - 0x13d4  :  248 - 0xf8
    "11111100", -- 5077 - 0x13d5  :  252 - 0xfc
    "11111100", -- 5078 - 0x13d6  :  252 - 0xfc
    "11111100", -- 5079 - 0x13d7  :  252 - 0xfc
    "00000000", -- 5080 - 0x13d8  :    0 - 0x0
    "11000000", -- 5081 - 0x13d9  :  192 - 0xc0
    "11110000", -- 5082 - 0x13da  :  240 - 0xf0
    "11111000", -- 5083 - 0x13db  :  248 - 0xf8
    "11111000", -- 5084 - 0x13dc  :  248 - 0xf8
    "11111100", -- 5085 - 0x13dd  :  252 - 0xfc
    "11111100", -- 5086 - 0x13de  :  252 - 0xfc
    "11111100", -- 5087 - 0x13df  :  252 - 0xfc
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0 -- Background 0x3e
    "00000011", -- 5089 - 0x13e1  :    3 - 0x3
    "00001111", -- 5090 - 0x13e2  :   15 - 0xf
    "00111111", -- 5091 - 0x13e3  :   63 - 0x3f
    "00111111", -- 5092 - 0x13e4  :   63 - 0x3f
    "00011111", -- 5093 - 0x13e5  :   31 - 0x1f
    "00000111", -- 5094 - 0x13e6  :    7 - 0x7
    "00000000", -- 5095 - 0x13e7  :    0 - 0x0
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000011", -- 5097 - 0x13e9  :    3 - 0x3
    "00001111", -- 5098 - 0x13ea  :   15 - 0xf
    "00111111", -- 5099 - 0x13eb  :   63 - 0x3f
    "00111111", -- 5100 - 0x13ec  :   63 - 0x3f
    "00011111", -- 5101 - 0x13ed  :   31 - 0x1f
    "00000111", -- 5102 - 0x13ee  :    7 - 0x7
    "00000000", -- 5103 - 0x13ef  :    0 - 0x0
    "11111100", -- 5104 - 0x13f0  :  252 - 0xfc -- Background 0x3f
    "11111100", -- 5105 - 0x13f1  :  252 - 0xfc
    "11111100", -- 5106 - 0x13f2  :  252 - 0xfc
    "11111000", -- 5107 - 0x13f3  :  248 - 0xf8
    "11111000", -- 5108 - 0x13f4  :  248 - 0xf8
    "11110000", -- 5109 - 0x13f5  :  240 - 0xf0
    "11000000", -- 5110 - 0x13f6  :  192 - 0xc0
    "00000000", -- 5111 - 0x13f7  :    0 - 0x0
    "11111100", -- 5112 - 0x13f8  :  252 - 0xfc
    "11111100", -- 5113 - 0x13f9  :  252 - 0xfc
    "11111100", -- 5114 - 0x13fa  :  252 - 0xfc
    "11111000", -- 5115 - 0x13fb  :  248 - 0xf8
    "11111000", -- 5116 - 0x13fc  :  248 - 0xf8
    "11110000", -- 5117 - 0x13fd  :  240 - 0xf0
    "11000000", -- 5118 - 0x13fe  :  192 - 0xc0
    "00000000", -- 5119 - 0x13ff  :    0 - 0x0
    "00000000", -- 5120 - 0x1400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 5121 - 0x1401  :    0 - 0x0
    "00000000", -- 5122 - 0x1402  :    0 - 0x0
    "00000000", -- 5123 - 0x1403  :    0 - 0x0
    "00000000", -- 5124 - 0x1404  :    0 - 0x0
    "00000000", -- 5125 - 0x1405  :    0 - 0x0
    "00000000", -- 5126 - 0x1406  :    0 - 0x0
    "00000000", -- 5127 - 0x1407  :    0 - 0x0
    "00000000", -- 5128 - 0x1408  :    0 - 0x0
    "00000000", -- 5129 - 0x1409  :    0 - 0x0
    "00000000", -- 5130 - 0x140a  :    0 - 0x0
    "00000000", -- 5131 - 0x140b  :    0 - 0x0
    "00000000", -- 5132 - 0x140c  :    0 - 0x0
    "00000000", -- 5133 - 0x140d  :    0 - 0x0
    "00000000", -- 5134 - 0x140e  :    0 - 0x0
    "00000000", -- 5135 - 0x140f  :    0 - 0x0
    "00011100", -- 5136 - 0x1410  :   28 - 0x1c -- Background 0x41
    "00110110", -- 5137 - 0x1411  :   54 - 0x36
    "01100011", -- 5138 - 0x1412  :   99 - 0x63
    "01100011", -- 5139 - 0x1413  :   99 - 0x63
    "01111111", -- 5140 - 0x1414  :  127 - 0x7f
    "01100011", -- 5141 - 0x1415  :   99 - 0x63
    "01100011", -- 5142 - 0x1416  :   99 - 0x63
    "00000000", -- 5143 - 0x1417  :    0 - 0x0
    "00000000", -- 5144 - 0x1418  :    0 - 0x0
    "00000000", -- 5145 - 0x1419  :    0 - 0x0
    "00000000", -- 5146 - 0x141a  :    0 - 0x0
    "00000000", -- 5147 - 0x141b  :    0 - 0x0
    "00000000", -- 5148 - 0x141c  :    0 - 0x0
    "00000000", -- 5149 - 0x141d  :    0 - 0x0
    "00000000", -- 5150 - 0x141e  :    0 - 0x0
    "00000000", -- 5151 - 0x141f  :    0 - 0x0
    "01111110", -- 5152 - 0x1420  :  126 - 0x7e -- Background 0x42
    "01100011", -- 5153 - 0x1421  :   99 - 0x63
    "01100011", -- 5154 - 0x1422  :   99 - 0x63
    "01111110", -- 5155 - 0x1423  :  126 - 0x7e
    "01100011", -- 5156 - 0x1424  :   99 - 0x63
    "01100011", -- 5157 - 0x1425  :   99 - 0x63
    "01111110", -- 5158 - 0x1426  :  126 - 0x7e
    "00000000", -- 5159 - 0x1427  :    0 - 0x0
    "00000000", -- 5160 - 0x1428  :    0 - 0x0
    "00000000", -- 5161 - 0x1429  :    0 - 0x0
    "00000000", -- 5162 - 0x142a  :    0 - 0x0
    "00000000", -- 5163 - 0x142b  :    0 - 0x0
    "00000000", -- 5164 - 0x142c  :    0 - 0x0
    "00000000", -- 5165 - 0x142d  :    0 - 0x0
    "00000000", -- 5166 - 0x142e  :    0 - 0x0
    "00000000", -- 5167 - 0x142f  :    0 - 0x0
    "00011110", -- 5168 - 0x1430  :   30 - 0x1e -- Background 0x43
    "00110011", -- 5169 - 0x1431  :   51 - 0x33
    "01100000", -- 5170 - 0x1432  :   96 - 0x60
    "01100000", -- 5171 - 0x1433  :   96 - 0x60
    "01100000", -- 5172 - 0x1434  :   96 - 0x60
    "00110011", -- 5173 - 0x1435  :   51 - 0x33
    "00011110", -- 5174 - 0x1436  :   30 - 0x1e
    "00000000", -- 5175 - 0x1437  :    0 - 0x0
    "00000000", -- 5176 - 0x1438  :    0 - 0x0
    "00000000", -- 5177 - 0x1439  :    0 - 0x0
    "00000000", -- 5178 - 0x143a  :    0 - 0x0
    "00000000", -- 5179 - 0x143b  :    0 - 0x0
    "00000000", -- 5180 - 0x143c  :    0 - 0x0
    "00000000", -- 5181 - 0x143d  :    0 - 0x0
    "00000000", -- 5182 - 0x143e  :    0 - 0x0
    "00000000", -- 5183 - 0x143f  :    0 - 0x0
    "01111100", -- 5184 - 0x1440  :  124 - 0x7c -- Background 0x44
    "01100110", -- 5185 - 0x1441  :  102 - 0x66
    "01100011", -- 5186 - 0x1442  :   99 - 0x63
    "01100011", -- 5187 - 0x1443  :   99 - 0x63
    "01100011", -- 5188 - 0x1444  :   99 - 0x63
    "01100110", -- 5189 - 0x1445  :  102 - 0x66
    "01111100", -- 5190 - 0x1446  :  124 - 0x7c
    "00000000", -- 5191 - 0x1447  :    0 - 0x0
    "00000000", -- 5192 - 0x1448  :    0 - 0x0
    "00000000", -- 5193 - 0x1449  :    0 - 0x0
    "00000000", -- 5194 - 0x144a  :    0 - 0x0
    "00000000", -- 5195 - 0x144b  :    0 - 0x0
    "00000000", -- 5196 - 0x144c  :    0 - 0x0
    "00000000", -- 5197 - 0x144d  :    0 - 0x0
    "00000000", -- 5198 - 0x144e  :    0 - 0x0
    "00000000", -- 5199 - 0x144f  :    0 - 0x0
    "01111111", -- 5200 - 0x1450  :  127 - 0x7f -- Background 0x45
    "01100000", -- 5201 - 0x1451  :   96 - 0x60
    "01100000", -- 5202 - 0x1452  :   96 - 0x60
    "01111110", -- 5203 - 0x1453  :  126 - 0x7e
    "01100000", -- 5204 - 0x1454  :   96 - 0x60
    "01100000", -- 5205 - 0x1455  :   96 - 0x60
    "01111111", -- 5206 - 0x1456  :  127 - 0x7f
    "00000000", -- 5207 - 0x1457  :    0 - 0x0
    "00000000", -- 5208 - 0x1458  :    0 - 0x0
    "00000000", -- 5209 - 0x1459  :    0 - 0x0
    "00000000", -- 5210 - 0x145a  :    0 - 0x0
    "00000000", -- 5211 - 0x145b  :    0 - 0x0
    "00000000", -- 5212 - 0x145c  :    0 - 0x0
    "00000000", -- 5213 - 0x145d  :    0 - 0x0
    "00000000", -- 5214 - 0x145e  :    0 - 0x0
    "00000000", -- 5215 - 0x145f  :    0 - 0x0
    "01111111", -- 5216 - 0x1460  :  127 - 0x7f -- Background 0x46
    "01100000", -- 5217 - 0x1461  :   96 - 0x60
    "01100000", -- 5218 - 0x1462  :   96 - 0x60
    "01111110", -- 5219 - 0x1463  :  126 - 0x7e
    "01100000", -- 5220 - 0x1464  :   96 - 0x60
    "01100000", -- 5221 - 0x1465  :   96 - 0x60
    "01100000", -- 5222 - 0x1466  :   96 - 0x60
    "00000000", -- 5223 - 0x1467  :    0 - 0x0
    "00000000", -- 5224 - 0x1468  :    0 - 0x0
    "00000000", -- 5225 - 0x1469  :    0 - 0x0
    "00000000", -- 5226 - 0x146a  :    0 - 0x0
    "00000000", -- 5227 - 0x146b  :    0 - 0x0
    "00000000", -- 5228 - 0x146c  :    0 - 0x0
    "00000000", -- 5229 - 0x146d  :    0 - 0x0
    "00000000", -- 5230 - 0x146e  :    0 - 0x0
    "00000000", -- 5231 - 0x146f  :    0 - 0x0
    "00011111", -- 5232 - 0x1470  :   31 - 0x1f -- Background 0x47
    "00110000", -- 5233 - 0x1471  :   48 - 0x30
    "01100000", -- 5234 - 0x1472  :   96 - 0x60
    "01100111", -- 5235 - 0x1473  :  103 - 0x67
    "01100011", -- 5236 - 0x1474  :   99 - 0x63
    "00110011", -- 5237 - 0x1475  :   51 - 0x33
    "00011111", -- 5238 - 0x1476  :   31 - 0x1f
    "00000000", -- 5239 - 0x1477  :    0 - 0x0
    "00000000", -- 5240 - 0x1478  :    0 - 0x0
    "00000000", -- 5241 - 0x1479  :    0 - 0x0
    "00000000", -- 5242 - 0x147a  :    0 - 0x0
    "00000000", -- 5243 - 0x147b  :    0 - 0x0
    "00000000", -- 5244 - 0x147c  :    0 - 0x0
    "00000000", -- 5245 - 0x147d  :    0 - 0x0
    "00000000", -- 5246 - 0x147e  :    0 - 0x0
    "00000000", -- 5247 - 0x147f  :    0 - 0x0
    "01100011", -- 5248 - 0x1480  :   99 - 0x63 -- Background 0x48
    "01100011", -- 5249 - 0x1481  :   99 - 0x63
    "01100011", -- 5250 - 0x1482  :   99 - 0x63
    "01111111", -- 5251 - 0x1483  :  127 - 0x7f
    "01100011", -- 5252 - 0x1484  :   99 - 0x63
    "01100011", -- 5253 - 0x1485  :   99 - 0x63
    "01100011", -- 5254 - 0x1486  :   99 - 0x63
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "00000000", -- 5257 - 0x1489  :    0 - 0x0
    "00000000", -- 5258 - 0x148a  :    0 - 0x0
    "00000000", -- 5259 - 0x148b  :    0 - 0x0
    "00000000", -- 5260 - 0x148c  :    0 - 0x0
    "00000000", -- 5261 - 0x148d  :    0 - 0x0
    "00000000", -- 5262 - 0x148e  :    0 - 0x0
    "00000000", -- 5263 - 0x148f  :    0 - 0x0
    "00111111", -- 5264 - 0x1490  :   63 - 0x3f -- Background 0x49
    "00001100", -- 5265 - 0x1491  :   12 - 0xc
    "00001100", -- 5266 - 0x1492  :   12 - 0xc
    "00001100", -- 5267 - 0x1493  :   12 - 0xc
    "00001100", -- 5268 - 0x1494  :   12 - 0xc
    "00001100", -- 5269 - 0x1495  :   12 - 0xc
    "00111111", -- 5270 - 0x1496  :   63 - 0x3f
    "00000000", -- 5271 - 0x1497  :    0 - 0x0
    "00000000", -- 5272 - 0x1498  :    0 - 0x0
    "00000000", -- 5273 - 0x1499  :    0 - 0x0
    "00000000", -- 5274 - 0x149a  :    0 - 0x0
    "00000000", -- 5275 - 0x149b  :    0 - 0x0
    "00000000", -- 5276 - 0x149c  :    0 - 0x0
    "00000000", -- 5277 - 0x149d  :    0 - 0x0
    "00000000", -- 5278 - 0x149e  :    0 - 0x0
    "00000000", -- 5279 - 0x149f  :    0 - 0x0
    "00000011", -- 5280 - 0x14a0  :    3 - 0x3 -- Background 0x4a
    "00000011", -- 5281 - 0x14a1  :    3 - 0x3
    "00000011", -- 5282 - 0x14a2  :    3 - 0x3
    "00000011", -- 5283 - 0x14a3  :    3 - 0x3
    "00000011", -- 5284 - 0x14a4  :    3 - 0x3
    "01100011", -- 5285 - 0x14a5  :   99 - 0x63
    "00111110", -- 5286 - 0x14a6  :   62 - 0x3e
    "00000000", -- 5287 - 0x14a7  :    0 - 0x0
    "00000000", -- 5288 - 0x14a8  :    0 - 0x0
    "00000000", -- 5289 - 0x14a9  :    0 - 0x0
    "00000000", -- 5290 - 0x14aa  :    0 - 0x0
    "00000000", -- 5291 - 0x14ab  :    0 - 0x0
    "00000000", -- 5292 - 0x14ac  :    0 - 0x0
    "00000000", -- 5293 - 0x14ad  :    0 - 0x0
    "00000000", -- 5294 - 0x14ae  :    0 - 0x0
    "00000000", -- 5295 - 0x14af  :    0 - 0x0
    "01100011", -- 5296 - 0x14b0  :   99 - 0x63 -- Background 0x4b
    "01100110", -- 5297 - 0x14b1  :  102 - 0x66
    "01101100", -- 5298 - 0x14b2  :  108 - 0x6c
    "01111000", -- 5299 - 0x14b3  :  120 - 0x78
    "01111100", -- 5300 - 0x14b4  :  124 - 0x7c
    "01100110", -- 5301 - 0x14b5  :  102 - 0x66
    "01100011", -- 5302 - 0x14b6  :   99 - 0x63
    "00000000", -- 5303 - 0x14b7  :    0 - 0x0
    "00000000", -- 5304 - 0x14b8  :    0 - 0x0
    "00000000", -- 5305 - 0x14b9  :    0 - 0x0
    "00000000", -- 5306 - 0x14ba  :    0 - 0x0
    "00000000", -- 5307 - 0x14bb  :    0 - 0x0
    "00000000", -- 5308 - 0x14bc  :    0 - 0x0
    "00000000", -- 5309 - 0x14bd  :    0 - 0x0
    "00000000", -- 5310 - 0x14be  :    0 - 0x0
    "00000000", -- 5311 - 0x14bf  :    0 - 0x0
    "01100000", -- 5312 - 0x14c0  :   96 - 0x60 -- Background 0x4c
    "01100000", -- 5313 - 0x14c1  :   96 - 0x60
    "01100000", -- 5314 - 0x14c2  :   96 - 0x60
    "01100000", -- 5315 - 0x14c3  :   96 - 0x60
    "01100000", -- 5316 - 0x14c4  :   96 - 0x60
    "01100000", -- 5317 - 0x14c5  :   96 - 0x60
    "01111111", -- 5318 - 0x14c6  :  127 - 0x7f
    "00000000", -- 5319 - 0x14c7  :    0 - 0x0
    "00000000", -- 5320 - 0x14c8  :    0 - 0x0
    "00000000", -- 5321 - 0x14c9  :    0 - 0x0
    "00000000", -- 5322 - 0x14ca  :    0 - 0x0
    "00000000", -- 5323 - 0x14cb  :    0 - 0x0
    "00000000", -- 5324 - 0x14cc  :    0 - 0x0
    "00000000", -- 5325 - 0x14cd  :    0 - 0x0
    "00000000", -- 5326 - 0x14ce  :    0 - 0x0
    "00000000", -- 5327 - 0x14cf  :    0 - 0x0
    "01100011", -- 5328 - 0x14d0  :   99 - 0x63 -- Background 0x4d
    "01110111", -- 5329 - 0x14d1  :  119 - 0x77
    "01111111", -- 5330 - 0x14d2  :  127 - 0x7f
    "01111111", -- 5331 - 0x14d3  :  127 - 0x7f
    "01101011", -- 5332 - 0x14d4  :  107 - 0x6b
    "01100011", -- 5333 - 0x14d5  :   99 - 0x63
    "01100011", -- 5334 - 0x14d6  :   99 - 0x63
    "00000000", -- 5335 - 0x14d7  :    0 - 0x0
    "00000000", -- 5336 - 0x14d8  :    0 - 0x0
    "00000000", -- 5337 - 0x14d9  :    0 - 0x0
    "00000000", -- 5338 - 0x14da  :    0 - 0x0
    "00000000", -- 5339 - 0x14db  :    0 - 0x0
    "00000000", -- 5340 - 0x14dc  :    0 - 0x0
    "00000000", -- 5341 - 0x14dd  :    0 - 0x0
    "00000000", -- 5342 - 0x14de  :    0 - 0x0
    "00000000", -- 5343 - 0x14df  :    0 - 0x0
    "01100011", -- 5344 - 0x14e0  :   99 - 0x63 -- Background 0x4e
    "01110011", -- 5345 - 0x14e1  :  115 - 0x73
    "01111011", -- 5346 - 0x14e2  :  123 - 0x7b
    "01111111", -- 5347 - 0x14e3  :  127 - 0x7f
    "01101111", -- 5348 - 0x14e4  :  111 - 0x6f
    "01100111", -- 5349 - 0x14e5  :  103 - 0x67
    "01100011", -- 5350 - 0x14e6  :   99 - 0x63
    "00000000", -- 5351 - 0x14e7  :    0 - 0x0
    "00000000", -- 5352 - 0x14e8  :    0 - 0x0
    "00000000", -- 5353 - 0x14e9  :    0 - 0x0
    "00000000", -- 5354 - 0x14ea  :    0 - 0x0
    "00000000", -- 5355 - 0x14eb  :    0 - 0x0
    "00000000", -- 5356 - 0x14ec  :    0 - 0x0
    "00000000", -- 5357 - 0x14ed  :    0 - 0x0
    "00000000", -- 5358 - 0x14ee  :    0 - 0x0
    "00000000", -- 5359 - 0x14ef  :    0 - 0x0
    "00111110", -- 5360 - 0x14f0  :   62 - 0x3e -- Background 0x4f
    "01100011", -- 5361 - 0x14f1  :   99 - 0x63
    "01100011", -- 5362 - 0x14f2  :   99 - 0x63
    "01100011", -- 5363 - 0x14f3  :   99 - 0x63
    "01100011", -- 5364 - 0x14f4  :   99 - 0x63
    "01100011", -- 5365 - 0x14f5  :   99 - 0x63
    "00111110", -- 5366 - 0x14f6  :   62 - 0x3e
    "00000000", -- 5367 - 0x14f7  :    0 - 0x0
    "00000000", -- 5368 - 0x14f8  :    0 - 0x0
    "00000000", -- 5369 - 0x14f9  :    0 - 0x0
    "00000000", -- 5370 - 0x14fa  :    0 - 0x0
    "00000000", -- 5371 - 0x14fb  :    0 - 0x0
    "00000000", -- 5372 - 0x14fc  :    0 - 0x0
    "00000000", -- 5373 - 0x14fd  :    0 - 0x0
    "00000000", -- 5374 - 0x14fe  :    0 - 0x0
    "00000000", -- 5375 - 0x14ff  :    0 - 0x0
    "01111110", -- 5376 - 0x1500  :  126 - 0x7e -- Background 0x50
    "01100011", -- 5377 - 0x1501  :   99 - 0x63
    "01100011", -- 5378 - 0x1502  :   99 - 0x63
    "01100011", -- 5379 - 0x1503  :   99 - 0x63
    "01111110", -- 5380 - 0x1504  :  126 - 0x7e
    "01100000", -- 5381 - 0x1505  :   96 - 0x60
    "01100000", -- 5382 - 0x1506  :   96 - 0x60
    "00000000", -- 5383 - 0x1507  :    0 - 0x0
    "00000000", -- 5384 - 0x1508  :    0 - 0x0
    "00000000", -- 5385 - 0x1509  :    0 - 0x0
    "00000000", -- 5386 - 0x150a  :    0 - 0x0
    "00000000", -- 5387 - 0x150b  :    0 - 0x0
    "00000000", -- 5388 - 0x150c  :    0 - 0x0
    "00000000", -- 5389 - 0x150d  :    0 - 0x0
    "00000000", -- 5390 - 0x150e  :    0 - 0x0
    "00000000", -- 5391 - 0x150f  :    0 - 0x0
    "00111110", -- 5392 - 0x1510  :   62 - 0x3e -- Background 0x51
    "01100011", -- 5393 - 0x1511  :   99 - 0x63
    "01100011", -- 5394 - 0x1512  :   99 - 0x63
    "01100011", -- 5395 - 0x1513  :   99 - 0x63
    "01101111", -- 5396 - 0x1514  :  111 - 0x6f
    "01100110", -- 5397 - 0x1515  :  102 - 0x66
    "00111101", -- 5398 - 0x1516  :   61 - 0x3d
    "00000000", -- 5399 - 0x1517  :    0 - 0x0
    "00000000", -- 5400 - 0x1518  :    0 - 0x0
    "00000000", -- 5401 - 0x1519  :    0 - 0x0
    "00000000", -- 5402 - 0x151a  :    0 - 0x0
    "00000000", -- 5403 - 0x151b  :    0 - 0x0
    "00000000", -- 5404 - 0x151c  :    0 - 0x0
    "00000000", -- 5405 - 0x151d  :    0 - 0x0
    "00000000", -- 5406 - 0x151e  :    0 - 0x0
    "00000000", -- 5407 - 0x151f  :    0 - 0x0
    "01111110", -- 5408 - 0x1520  :  126 - 0x7e -- Background 0x52
    "01100011", -- 5409 - 0x1521  :   99 - 0x63
    "01100011", -- 5410 - 0x1522  :   99 - 0x63
    "01100111", -- 5411 - 0x1523  :  103 - 0x67
    "01111100", -- 5412 - 0x1524  :  124 - 0x7c
    "01101110", -- 5413 - 0x1525  :  110 - 0x6e
    "01100111", -- 5414 - 0x1526  :  103 - 0x67
    "00000000", -- 5415 - 0x1527  :    0 - 0x0
    "00000000", -- 5416 - 0x1528  :    0 - 0x0
    "00000000", -- 5417 - 0x1529  :    0 - 0x0
    "00000000", -- 5418 - 0x152a  :    0 - 0x0
    "00000000", -- 5419 - 0x152b  :    0 - 0x0
    "00000000", -- 5420 - 0x152c  :    0 - 0x0
    "00000000", -- 5421 - 0x152d  :    0 - 0x0
    "00000000", -- 5422 - 0x152e  :    0 - 0x0
    "00000000", -- 5423 - 0x152f  :    0 - 0x0
    "00111100", -- 5424 - 0x1530  :   60 - 0x3c -- Background 0x53
    "01100110", -- 5425 - 0x1531  :  102 - 0x66
    "01100000", -- 5426 - 0x1532  :   96 - 0x60
    "00111110", -- 5427 - 0x1533  :   62 - 0x3e
    "00000011", -- 5428 - 0x1534  :    3 - 0x3
    "01100011", -- 5429 - 0x1535  :   99 - 0x63
    "00111110", -- 5430 - 0x1536  :   62 - 0x3e
    "00000000", -- 5431 - 0x1537  :    0 - 0x0
    "00000000", -- 5432 - 0x1538  :    0 - 0x0
    "00000000", -- 5433 - 0x1539  :    0 - 0x0
    "00000000", -- 5434 - 0x153a  :    0 - 0x0
    "00000000", -- 5435 - 0x153b  :    0 - 0x0
    "00000000", -- 5436 - 0x153c  :    0 - 0x0
    "00000000", -- 5437 - 0x153d  :    0 - 0x0
    "00000000", -- 5438 - 0x153e  :    0 - 0x0
    "00000000", -- 5439 - 0x153f  :    0 - 0x0
    "00111111", -- 5440 - 0x1540  :   63 - 0x3f -- Background 0x54
    "00001100", -- 5441 - 0x1541  :   12 - 0xc
    "00001100", -- 5442 - 0x1542  :   12 - 0xc
    "00001100", -- 5443 - 0x1543  :   12 - 0xc
    "00001100", -- 5444 - 0x1544  :   12 - 0xc
    "00001100", -- 5445 - 0x1545  :   12 - 0xc
    "00001100", -- 5446 - 0x1546  :   12 - 0xc
    "00000000", -- 5447 - 0x1547  :    0 - 0x0
    "00000000", -- 5448 - 0x1548  :    0 - 0x0
    "00000000", -- 5449 - 0x1549  :    0 - 0x0
    "00000000", -- 5450 - 0x154a  :    0 - 0x0
    "00000000", -- 5451 - 0x154b  :    0 - 0x0
    "00000000", -- 5452 - 0x154c  :    0 - 0x0
    "00000000", -- 5453 - 0x154d  :    0 - 0x0
    "00000000", -- 5454 - 0x154e  :    0 - 0x0
    "00000000", -- 5455 - 0x154f  :    0 - 0x0
    "01100011", -- 5456 - 0x1550  :   99 - 0x63 -- Background 0x55
    "01100011", -- 5457 - 0x1551  :   99 - 0x63
    "01100011", -- 5458 - 0x1552  :   99 - 0x63
    "01100011", -- 5459 - 0x1553  :   99 - 0x63
    "01100011", -- 5460 - 0x1554  :   99 - 0x63
    "01100011", -- 5461 - 0x1555  :   99 - 0x63
    "00111110", -- 5462 - 0x1556  :   62 - 0x3e
    "00000000", -- 5463 - 0x1557  :    0 - 0x0
    "00000000", -- 5464 - 0x1558  :    0 - 0x0
    "00000000", -- 5465 - 0x1559  :    0 - 0x0
    "00000000", -- 5466 - 0x155a  :    0 - 0x0
    "00000000", -- 5467 - 0x155b  :    0 - 0x0
    "00000000", -- 5468 - 0x155c  :    0 - 0x0
    "00000000", -- 5469 - 0x155d  :    0 - 0x0
    "00000000", -- 5470 - 0x155e  :    0 - 0x0
    "00000000", -- 5471 - 0x155f  :    0 - 0x0
    "01100011", -- 5472 - 0x1560  :   99 - 0x63 -- Background 0x56
    "01100011", -- 5473 - 0x1561  :   99 - 0x63
    "01100011", -- 5474 - 0x1562  :   99 - 0x63
    "01110111", -- 5475 - 0x1563  :  119 - 0x77
    "00111110", -- 5476 - 0x1564  :   62 - 0x3e
    "00011100", -- 5477 - 0x1565  :   28 - 0x1c
    "00001000", -- 5478 - 0x1566  :    8 - 0x8
    "00000000", -- 5479 - 0x1567  :    0 - 0x0
    "00000000", -- 5480 - 0x1568  :    0 - 0x0
    "00000000", -- 5481 - 0x1569  :    0 - 0x0
    "00000000", -- 5482 - 0x156a  :    0 - 0x0
    "00000000", -- 5483 - 0x156b  :    0 - 0x0
    "00000000", -- 5484 - 0x156c  :    0 - 0x0
    "00000000", -- 5485 - 0x156d  :    0 - 0x0
    "00000000", -- 5486 - 0x156e  :    0 - 0x0
    "00000000", -- 5487 - 0x156f  :    0 - 0x0
    "01100011", -- 5488 - 0x1570  :   99 - 0x63 -- Background 0x57
    "01100011", -- 5489 - 0x1571  :   99 - 0x63
    "01101011", -- 5490 - 0x1572  :  107 - 0x6b
    "01111111", -- 5491 - 0x1573  :  127 - 0x7f
    "01111111", -- 5492 - 0x1574  :  127 - 0x7f
    "01110111", -- 5493 - 0x1575  :  119 - 0x77
    "01100011", -- 5494 - 0x1576  :   99 - 0x63
    "00000000", -- 5495 - 0x1577  :    0 - 0x0
    "00000000", -- 5496 - 0x1578  :    0 - 0x0
    "00000000", -- 5497 - 0x1579  :    0 - 0x0
    "00000000", -- 5498 - 0x157a  :    0 - 0x0
    "00000000", -- 5499 - 0x157b  :    0 - 0x0
    "00000000", -- 5500 - 0x157c  :    0 - 0x0
    "00000000", -- 5501 - 0x157d  :    0 - 0x0
    "00000000", -- 5502 - 0x157e  :    0 - 0x0
    "00000000", -- 5503 - 0x157f  :    0 - 0x0
    "01100011", -- 5504 - 0x1580  :   99 - 0x63 -- Background 0x58
    "01110111", -- 5505 - 0x1581  :  119 - 0x77
    "00111110", -- 5506 - 0x1582  :   62 - 0x3e
    "00011100", -- 5507 - 0x1583  :   28 - 0x1c
    "00111110", -- 5508 - 0x1584  :   62 - 0x3e
    "01110111", -- 5509 - 0x1585  :  119 - 0x77
    "01100011", -- 5510 - 0x1586  :   99 - 0x63
    "00000000", -- 5511 - 0x1587  :    0 - 0x0
    "00000000", -- 5512 - 0x1588  :    0 - 0x0
    "00000000", -- 5513 - 0x1589  :    0 - 0x0
    "00000000", -- 5514 - 0x158a  :    0 - 0x0
    "00000000", -- 5515 - 0x158b  :    0 - 0x0
    "00000000", -- 5516 - 0x158c  :    0 - 0x0
    "00000000", -- 5517 - 0x158d  :    0 - 0x0
    "00000000", -- 5518 - 0x158e  :    0 - 0x0
    "00000000", -- 5519 - 0x158f  :    0 - 0x0
    "00110011", -- 5520 - 0x1590  :   51 - 0x33 -- Background 0x59
    "00110011", -- 5521 - 0x1591  :   51 - 0x33
    "00110011", -- 5522 - 0x1592  :   51 - 0x33
    "00011110", -- 5523 - 0x1593  :   30 - 0x1e
    "00001100", -- 5524 - 0x1594  :   12 - 0xc
    "00001100", -- 5525 - 0x1595  :   12 - 0xc
    "00001100", -- 5526 - 0x1596  :   12 - 0xc
    "00000000", -- 5527 - 0x1597  :    0 - 0x0
    "00000000", -- 5528 - 0x1598  :    0 - 0x0
    "00000000", -- 5529 - 0x1599  :    0 - 0x0
    "00000000", -- 5530 - 0x159a  :    0 - 0x0
    "00000000", -- 5531 - 0x159b  :    0 - 0x0
    "00000000", -- 5532 - 0x159c  :    0 - 0x0
    "00000000", -- 5533 - 0x159d  :    0 - 0x0
    "00000000", -- 5534 - 0x159e  :    0 - 0x0
    "00000000", -- 5535 - 0x159f  :    0 - 0x0
    "01111111", -- 5536 - 0x15a0  :  127 - 0x7f -- Background 0x5a
    "00000111", -- 5537 - 0x15a1  :    7 - 0x7
    "00001110", -- 5538 - 0x15a2  :   14 - 0xe
    "00011100", -- 5539 - 0x15a3  :   28 - 0x1c
    "00111000", -- 5540 - 0x15a4  :   56 - 0x38
    "01110000", -- 5541 - 0x15a5  :  112 - 0x70
    "01111111", -- 5542 - 0x15a6  :  127 - 0x7f
    "00000000", -- 5543 - 0x15a7  :    0 - 0x0
    "00000000", -- 5544 - 0x15a8  :    0 - 0x0
    "00000000", -- 5545 - 0x15a9  :    0 - 0x0
    "00000000", -- 5546 - 0x15aa  :    0 - 0x0
    "00000000", -- 5547 - 0x15ab  :    0 - 0x0
    "00000000", -- 5548 - 0x15ac  :    0 - 0x0
    "00000000", -- 5549 - 0x15ad  :    0 - 0x0
    "00000000", -- 5550 - 0x15ae  :    0 - 0x0
    "00000000", -- 5551 - 0x15af  :    0 - 0x0
    "00000000", -- 5552 - 0x15b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 5553 - 0x15b1  :    0 - 0x0
    "00000000", -- 5554 - 0x15b2  :    0 - 0x0
    "00000000", -- 5555 - 0x15b3  :    0 - 0x0
    "00000000", -- 5556 - 0x15b4  :    0 - 0x0
    "00110000", -- 5557 - 0x15b5  :   48 - 0x30
    "00110000", -- 5558 - 0x15b6  :   48 - 0x30
    "00000000", -- 5559 - 0x15b7  :    0 - 0x0
    "00000000", -- 5560 - 0x15b8  :    0 - 0x0
    "00000000", -- 5561 - 0x15b9  :    0 - 0x0
    "00000000", -- 5562 - 0x15ba  :    0 - 0x0
    "00000000", -- 5563 - 0x15bb  :    0 - 0x0
    "00000000", -- 5564 - 0x15bc  :    0 - 0x0
    "00000000", -- 5565 - 0x15bd  :    0 - 0x0
    "00000000", -- 5566 - 0x15be  :    0 - 0x0
    "00000000", -- 5567 - 0x15bf  :    0 - 0x0
    "11000000", -- 5568 - 0x15c0  :  192 - 0xc0 -- Background 0x5c
    "11110000", -- 5569 - 0x15c1  :  240 - 0xf0
    "11111100", -- 5570 - 0x15c2  :  252 - 0xfc
    "11111111", -- 5571 - 0x15c3  :  255 - 0xff
    "11111100", -- 5572 - 0x15c4  :  252 - 0xfc
    "11110000", -- 5573 - 0x15c5  :  240 - 0xf0
    "11000000", -- 5574 - 0x15c6  :  192 - 0xc0
    "00000000", -- 5575 - 0x15c7  :    0 - 0x0
    "00000000", -- 5576 - 0x15c8  :    0 - 0x0
    "00000000", -- 5577 - 0x15c9  :    0 - 0x0
    "00000000", -- 5578 - 0x15ca  :    0 - 0x0
    "00000000", -- 5579 - 0x15cb  :    0 - 0x0
    "00000000", -- 5580 - 0x15cc  :    0 - 0x0
    "00000000", -- 5581 - 0x15cd  :    0 - 0x0
    "00000000", -- 5582 - 0x15ce  :    0 - 0x0
    "00000000", -- 5583 - 0x15cf  :    0 - 0x0
    "00111100", -- 5584 - 0x15d0  :   60 - 0x3c -- Background 0x5d
    "01000010", -- 5585 - 0x15d1  :   66 - 0x42
    "10011001", -- 5586 - 0x15d2  :  153 - 0x99
    "10100001", -- 5587 - 0x15d3  :  161 - 0xa1
    "10100001", -- 5588 - 0x15d4  :  161 - 0xa1
    "10011001", -- 5589 - 0x15d5  :  153 - 0x99
    "01000010", -- 5590 - 0x15d6  :   66 - 0x42
    "00111100", -- 5591 - 0x15d7  :   60 - 0x3c
    "00000000", -- 5592 - 0x15d8  :    0 - 0x0
    "00000000", -- 5593 - 0x15d9  :    0 - 0x0
    "00000000", -- 5594 - 0x15da  :    0 - 0x0
    "00000000", -- 5595 - 0x15db  :    0 - 0x0
    "00000000", -- 5596 - 0x15dc  :    0 - 0x0
    "00000000", -- 5597 - 0x15dd  :    0 - 0x0
    "00000000", -- 5598 - 0x15de  :    0 - 0x0
    "00000000", -- 5599 - 0x15df  :    0 - 0x0
    "00000000", -- 5600 - 0x15e0  :    0 - 0x0 -- Background 0x5e
    "00000000", -- 5601 - 0x15e1  :    0 - 0x0
    "00010000", -- 5602 - 0x15e2  :   16 - 0x10
    "00010000", -- 5603 - 0x15e3  :   16 - 0x10
    "00010000", -- 5604 - 0x15e4  :   16 - 0x10
    "00010000", -- 5605 - 0x15e5  :   16 - 0x10
    "00000000", -- 5606 - 0x15e6  :    0 - 0x0
    "00000000", -- 5607 - 0x15e7  :    0 - 0x0
    "00000000", -- 5608 - 0x15e8  :    0 - 0x0
    "00000000", -- 5609 - 0x15e9  :    0 - 0x0
    "00010000", -- 5610 - 0x15ea  :   16 - 0x10
    "00010000", -- 5611 - 0x15eb  :   16 - 0x10
    "00010000", -- 5612 - 0x15ec  :   16 - 0x10
    "00010000", -- 5613 - 0x15ed  :   16 - 0x10
    "00000000", -- 5614 - 0x15ee  :    0 - 0x0
    "00000000", -- 5615 - 0x15ef  :    0 - 0x0
    "00110110", -- 5616 - 0x15f0  :   54 - 0x36 -- Background 0x5f
    "00110110", -- 5617 - 0x15f1  :   54 - 0x36
    "00010010", -- 5618 - 0x15f2  :   18 - 0x12
    "00000000", -- 5619 - 0x15f3  :    0 - 0x0
    "00000000", -- 5620 - 0x15f4  :    0 - 0x0
    "00000000", -- 5621 - 0x15f5  :    0 - 0x0
    "00000000", -- 5622 - 0x15f6  :    0 - 0x0
    "00000000", -- 5623 - 0x15f7  :    0 - 0x0
    "00000000", -- 5624 - 0x15f8  :    0 - 0x0
    "00000000", -- 5625 - 0x15f9  :    0 - 0x0
    "00000000", -- 5626 - 0x15fa  :    0 - 0x0
    "00000000", -- 5627 - 0x15fb  :    0 - 0x0
    "00000000", -- 5628 - 0x15fc  :    0 - 0x0
    "00000000", -- 5629 - 0x15fd  :    0 - 0x0
    "00000000", -- 5630 - 0x15fe  :    0 - 0x0
    "00000000", -- 5631 - 0x15ff  :    0 - 0x0
    "00000000", -- 5632 - 0x1600  :    0 - 0x0 -- Background 0x60
    "00000000", -- 5633 - 0x1601  :    0 - 0x0
    "00000000", -- 5634 - 0x1602  :    0 - 0x0
    "00000000", -- 5635 - 0x1603  :    0 - 0x0
    "00000000", -- 5636 - 0x1604  :    0 - 0x0
    "00000001", -- 5637 - 0x1605  :    1 - 0x1
    "00011110", -- 5638 - 0x1606  :   30 - 0x1e
    "00111011", -- 5639 - 0x1607  :   59 - 0x3b
    "00000000", -- 5640 - 0x1608  :    0 - 0x0
    "00000000", -- 5641 - 0x1609  :    0 - 0x0
    "00000000", -- 5642 - 0x160a  :    0 - 0x0
    "00000000", -- 5643 - 0x160b  :    0 - 0x0
    "00000000", -- 5644 - 0x160c  :    0 - 0x0
    "00000000", -- 5645 - 0x160d  :    0 - 0x0
    "00000000", -- 5646 - 0x160e  :    0 - 0x0
    "00000000", -- 5647 - 0x160f  :    0 - 0x0
    "00000000", -- 5648 - 0x1610  :    0 - 0x0 -- Background 0x61
    "00000000", -- 5649 - 0x1611  :    0 - 0x0
    "00001100", -- 5650 - 0x1612  :   12 - 0xc
    "00111100", -- 5651 - 0x1613  :   60 - 0x3c
    "11010000", -- 5652 - 0x1614  :  208 - 0xd0
    "00010000", -- 5653 - 0x1615  :   16 - 0x10
    "00100000", -- 5654 - 0x1616  :   32 - 0x20
    "01000000", -- 5655 - 0x1617  :   64 - 0x40
    "00000000", -- 5656 - 0x1618  :    0 - 0x0
    "00000000", -- 5657 - 0x1619  :    0 - 0x0
    "00000000", -- 5658 - 0x161a  :    0 - 0x0
    "00000000", -- 5659 - 0x161b  :    0 - 0x0
    "00000000", -- 5660 - 0x161c  :    0 - 0x0
    "00000000", -- 5661 - 0x161d  :    0 - 0x0
    "00000000", -- 5662 - 0x161e  :    0 - 0x0
    "00000000", -- 5663 - 0x161f  :    0 - 0x0
    "00111110", -- 5664 - 0x1620  :   62 - 0x3e -- Background 0x62
    "00101101", -- 5665 - 0x1621  :   45 - 0x2d
    "00110101", -- 5666 - 0x1622  :   53 - 0x35
    "00011101", -- 5667 - 0x1623  :   29 - 0x1d
    "00000001", -- 5668 - 0x1624  :    1 - 0x1
    "00000000", -- 5669 - 0x1625  :    0 - 0x0
    "00000000", -- 5670 - 0x1626  :    0 - 0x0
    "00000000", -- 5671 - 0x1627  :    0 - 0x0
    "00000000", -- 5672 - 0x1628  :    0 - 0x0
    "00000000", -- 5673 - 0x1629  :    0 - 0x0
    "00000000", -- 5674 - 0x162a  :    0 - 0x0
    "00000000", -- 5675 - 0x162b  :    0 - 0x0
    "00000000", -- 5676 - 0x162c  :    0 - 0x0
    "00000000", -- 5677 - 0x162d  :    0 - 0x0
    "00000000", -- 5678 - 0x162e  :    0 - 0x0
    "00000000", -- 5679 - 0x162f  :    0 - 0x0
    "10110000", -- 5680 - 0x1630  :  176 - 0xb0 -- Background 0x63
    "10111000", -- 5681 - 0x1631  :  184 - 0xb8
    "11111000", -- 5682 - 0x1632  :  248 - 0xf8
    "01111000", -- 5683 - 0x1633  :  120 - 0x78
    "10011000", -- 5684 - 0x1634  :  152 - 0x98
    "11110000", -- 5685 - 0x1635  :  240 - 0xf0
    "00000000", -- 5686 - 0x1636  :    0 - 0x0
    "00000000", -- 5687 - 0x1637  :    0 - 0x0
    "00000000", -- 5688 - 0x1638  :    0 - 0x0
    "00000000", -- 5689 - 0x1639  :    0 - 0x0
    "00000000", -- 5690 - 0x163a  :    0 - 0x0
    "00000000", -- 5691 - 0x163b  :    0 - 0x0
    "00000000", -- 5692 - 0x163c  :    0 - 0x0
    "00000000", -- 5693 - 0x163d  :    0 - 0x0
    "00000000", -- 5694 - 0x163e  :    0 - 0x0
    "00000000", -- 5695 - 0x163f  :    0 - 0x0
    "00000000", -- 5696 - 0x1640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 5697 - 0x1641  :    0 - 0x0
    "00000111", -- 5698 - 0x1642  :    7 - 0x7
    "00000011", -- 5699 - 0x1643  :    3 - 0x3
    "00001101", -- 5700 - 0x1644  :   13 - 0xd
    "00011110", -- 5701 - 0x1645  :   30 - 0x1e
    "00010111", -- 5702 - 0x1646  :   23 - 0x17
    "00011101", -- 5703 - 0x1647  :   29 - 0x1d
    "00000000", -- 5704 - 0x1648  :    0 - 0x0
    "00000000", -- 5705 - 0x1649  :    0 - 0x0
    "00000000", -- 5706 - 0x164a  :    0 - 0x0
    "00000000", -- 5707 - 0x164b  :    0 - 0x0
    "00000000", -- 5708 - 0x164c  :    0 - 0x0
    "00000000", -- 5709 - 0x164d  :    0 - 0x0
    "00000000", -- 5710 - 0x164e  :    0 - 0x0
    "00000000", -- 5711 - 0x164f  :    0 - 0x0
    "00000000", -- 5712 - 0x1650  :    0 - 0x0 -- Background 0x65
    "10000000", -- 5713 - 0x1651  :  128 - 0x80
    "01110000", -- 5714 - 0x1652  :  112 - 0x70
    "11100000", -- 5715 - 0x1653  :  224 - 0xe0
    "11011000", -- 5716 - 0x1654  :  216 - 0xd8
    "10111100", -- 5717 - 0x1655  :  188 - 0xbc
    "01110100", -- 5718 - 0x1656  :  116 - 0x74
    "11011100", -- 5719 - 0x1657  :  220 - 0xdc
    "00000000", -- 5720 - 0x1658  :    0 - 0x0
    "00000000", -- 5721 - 0x1659  :    0 - 0x0
    "00000000", -- 5722 - 0x165a  :    0 - 0x0
    "00000000", -- 5723 - 0x165b  :    0 - 0x0
    "00000000", -- 5724 - 0x165c  :    0 - 0x0
    "00000000", -- 5725 - 0x165d  :    0 - 0x0
    "00000000", -- 5726 - 0x165e  :    0 - 0x0
    "00000000", -- 5727 - 0x165f  :    0 - 0x0
    "00011111", -- 5728 - 0x1660  :   31 - 0x1f -- Background 0x66
    "00001011", -- 5729 - 0x1661  :   11 - 0xb
    "00001111", -- 5730 - 0x1662  :   15 - 0xf
    "00000101", -- 5731 - 0x1663  :    5 - 0x5
    "00000011", -- 5732 - 0x1664  :    3 - 0x3
    "00000001", -- 5733 - 0x1665  :    1 - 0x1
    "00000000", -- 5734 - 0x1666  :    0 - 0x0
    "00000000", -- 5735 - 0x1667  :    0 - 0x0
    "00000000", -- 5736 - 0x1668  :    0 - 0x0
    "00000000", -- 5737 - 0x1669  :    0 - 0x0
    "00000000", -- 5738 - 0x166a  :    0 - 0x0
    "00000000", -- 5739 - 0x166b  :    0 - 0x0
    "00000000", -- 5740 - 0x166c  :    0 - 0x0
    "00000000", -- 5741 - 0x166d  :    0 - 0x0
    "00000000", -- 5742 - 0x166e  :    0 - 0x0
    "00000000", -- 5743 - 0x166f  :    0 - 0x0
    "11111100", -- 5744 - 0x1670  :  252 - 0xfc -- Background 0x67
    "01101000", -- 5745 - 0x1671  :  104 - 0x68
    "11111000", -- 5746 - 0x1672  :  248 - 0xf8
    "10110000", -- 5747 - 0x1673  :  176 - 0xb0
    "11100000", -- 5748 - 0x1674  :  224 - 0xe0
    "10000000", -- 5749 - 0x1675  :  128 - 0x80
    "00000000", -- 5750 - 0x1676  :    0 - 0x0
    "00000000", -- 5751 - 0x1677  :    0 - 0x0
    "00000000", -- 5752 - 0x1678  :    0 - 0x0
    "00000000", -- 5753 - 0x1679  :    0 - 0x0
    "00000000", -- 5754 - 0x167a  :    0 - 0x0
    "00000000", -- 5755 - 0x167b  :    0 - 0x0
    "00000000", -- 5756 - 0x167c  :    0 - 0x0
    "00000000", -- 5757 - 0x167d  :    0 - 0x0
    "00000000", -- 5758 - 0x167e  :    0 - 0x0
    "00000000", -- 5759 - 0x167f  :    0 - 0x0
    "00000000", -- 5760 - 0x1680  :    0 - 0x0 -- Background 0x68
    "00000000", -- 5761 - 0x1681  :    0 - 0x0
    "00000000", -- 5762 - 0x1682  :    0 - 0x0
    "00000000", -- 5763 - 0x1683  :    0 - 0x0
    "00000000", -- 5764 - 0x1684  :    0 - 0x0
    "00000000", -- 5765 - 0x1685  :    0 - 0x0
    "00000000", -- 5766 - 0x1686  :    0 - 0x0
    "00000000", -- 5767 - 0x1687  :    0 - 0x0
    "00000000", -- 5768 - 0x1688  :    0 - 0x0
    "00000000", -- 5769 - 0x1689  :    0 - 0x0
    "00000000", -- 5770 - 0x168a  :    0 - 0x0
    "00000001", -- 5771 - 0x168b  :    1 - 0x1
    "00000001", -- 5772 - 0x168c  :    1 - 0x1
    "00001011", -- 5773 - 0x168d  :   11 - 0xb
    "00011100", -- 5774 - 0x168e  :   28 - 0x1c
    "00111111", -- 5775 - 0x168f  :   63 - 0x3f
    "00000000", -- 5776 - 0x1690  :    0 - 0x0 -- Background 0x69
    "00000000", -- 5777 - 0x1691  :    0 - 0x0
    "00000000", -- 5778 - 0x1692  :    0 - 0x0
    "00000000", -- 5779 - 0x1693  :    0 - 0x0
    "00000000", -- 5780 - 0x1694  :    0 - 0x0
    "00000000", -- 5781 - 0x1695  :    0 - 0x0
    "00000000", -- 5782 - 0x1696  :    0 - 0x0
    "00000000", -- 5783 - 0x1697  :    0 - 0x0
    "00000000", -- 5784 - 0x1698  :    0 - 0x0
    "00000000", -- 5785 - 0x1699  :    0 - 0x0
    "00110000", -- 5786 - 0x169a  :   48 - 0x30
    "01111000", -- 5787 - 0x169b  :  120 - 0x78
    "10000000", -- 5788 - 0x169c  :  128 - 0x80
    "11110000", -- 5789 - 0x169d  :  240 - 0xf0
    "11111000", -- 5790 - 0x169e  :  248 - 0xf8
    "11111100", -- 5791 - 0x169f  :  252 - 0xfc
    "00000000", -- 5792 - 0x16a0  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 5793 - 0x16a1  :    0 - 0x0
    "00000000", -- 5794 - 0x16a2  :    0 - 0x0
    "00000000", -- 5795 - 0x16a3  :    0 - 0x0
    "00000000", -- 5796 - 0x16a4  :    0 - 0x0
    "00000000", -- 5797 - 0x16a5  :    0 - 0x0
    "00000000", -- 5798 - 0x16a6  :    0 - 0x0
    "00000000", -- 5799 - 0x16a7  :    0 - 0x0
    "00111111", -- 5800 - 0x16a8  :   63 - 0x3f
    "00111111", -- 5801 - 0x16a9  :   63 - 0x3f
    "00111111", -- 5802 - 0x16aa  :   63 - 0x3f
    "00011111", -- 5803 - 0x16ab  :   31 - 0x1f
    "00011111", -- 5804 - 0x16ac  :   31 - 0x1f
    "00000111", -- 5805 - 0x16ad  :    7 - 0x7
    "00000000", -- 5806 - 0x16ae  :    0 - 0x0
    "00000000", -- 5807 - 0x16af  :    0 - 0x0
    "00000000", -- 5808 - 0x16b0  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 5809 - 0x16b1  :    0 - 0x0
    "00000000", -- 5810 - 0x16b2  :    0 - 0x0
    "00000000", -- 5811 - 0x16b3  :    0 - 0x0
    "00000000", -- 5812 - 0x16b4  :    0 - 0x0
    "00000000", -- 5813 - 0x16b5  :    0 - 0x0
    "00000000", -- 5814 - 0x16b6  :    0 - 0x0
    "00000000", -- 5815 - 0x16b7  :    0 - 0x0
    "11111100", -- 5816 - 0x16b8  :  252 - 0xfc
    "11101100", -- 5817 - 0x16b9  :  236 - 0xec
    "11101100", -- 5818 - 0x16ba  :  236 - 0xec
    "11011000", -- 5819 - 0x16bb  :  216 - 0xd8
    "11111000", -- 5820 - 0x16bc  :  248 - 0xf8
    "11100000", -- 5821 - 0x16bd  :  224 - 0xe0
    "00000000", -- 5822 - 0x16be  :    0 - 0x0
    "00000000", -- 5823 - 0x16bf  :    0 - 0x0
    "00000000", -- 5824 - 0x16c0  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 5825 - 0x16c1  :    0 - 0x0
    "00000001", -- 5826 - 0x16c2  :    1 - 0x1
    "00011101", -- 5827 - 0x16c3  :   29 - 0x1d
    "00111110", -- 5828 - 0x16c4  :   62 - 0x3e
    "00111111", -- 5829 - 0x16c5  :   63 - 0x3f
    "00111111", -- 5830 - 0x16c6  :   63 - 0x3f
    "00111111", -- 5831 - 0x16c7  :   63 - 0x3f
    "00000000", -- 5832 - 0x16c8  :    0 - 0x0
    "00000000", -- 5833 - 0x16c9  :    0 - 0x0
    "00000001", -- 5834 - 0x16ca  :    1 - 0x1
    "00011101", -- 5835 - 0x16cb  :   29 - 0x1d
    "00111110", -- 5836 - 0x16cc  :   62 - 0x3e
    "00111111", -- 5837 - 0x16cd  :   63 - 0x3f
    "00111111", -- 5838 - 0x16ce  :   63 - 0x3f
    "00111111", -- 5839 - 0x16cf  :   63 - 0x3f
    "00000000", -- 5840 - 0x16d0  :    0 - 0x0 -- Background 0x6d
    "10000000", -- 5841 - 0x16d1  :  128 - 0x80
    "00000000", -- 5842 - 0x16d2  :    0 - 0x0
    "01110000", -- 5843 - 0x16d3  :  112 - 0x70
    "11111000", -- 5844 - 0x16d4  :  248 - 0xf8
    "11111100", -- 5845 - 0x16d5  :  252 - 0xfc
    "11111100", -- 5846 - 0x16d6  :  252 - 0xfc
    "11111100", -- 5847 - 0x16d7  :  252 - 0xfc
    "00000000", -- 5848 - 0x16d8  :    0 - 0x0
    "10000000", -- 5849 - 0x16d9  :  128 - 0x80
    "00000000", -- 5850 - 0x16da  :    0 - 0x0
    "01110000", -- 5851 - 0x16db  :  112 - 0x70
    "11111000", -- 5852 - 0x16dc  :  248 - 0xf8
    "11111100", -- 5853 - 0x16dd  :  252 - 0xfc
    "11111100", -- 5854 - 0x16de  :  252 - 0xfc
    "11111100", -- 5855 - 0x16df  :  252 - 0xfc
    "00111111", -- 5856 - 0x16e0  :   63 - 0x3f -- Background 0x6e
    "00111111", -- 5857 - 0x16e1  :   63 - 0x3f
    "00011111", -- 5858 - 0x16e2  :   31 - 0x1f
    "00011111", -- 5859 - 0x16e3  :   31 - 0x1f
    "00001111", -- 5860 - 0x16e4  :   15 - 0xf
    "00000110", -- 5861 - 0x16e5  :    6 - 0x6
    "00000000", -- 5862 - 0x16e6  :    0 - 0x0
    "00000000", -- 5863 - 0x16e7  :    0 - 0x0
    "00111111", -- 5864 - 0x16e8  :   63 - 0x3f
    "00111111", -- 5865 - 0x16e9  :   63 - 0x3f
    "00011111", -- 5866 - 0x16ea  :   31 - 0x1f
    "00011111", -- 5867 - 0x16eb  :   31 - 0x1f
    "00001111", -- 5868 - 0x16ec  :   15 - 0xf
    "00000110", -- 5869 - 0x16ed  :    6 - 0x6
    "00000000", -- 5870 - 0x16ee  :    0 - 0x0
    "00000000", -- 5871 - 0x16ef  :    0 - 0x0
    "11101100", -- 5872 - 0x16f0  :  236 - 0xec -- Background 0x6f
    "11101100", -- 5873 - 0x16f1  :  236 - 0xec
    "11011000", -- 5874 - 0x16f2  :  216 - 0xd8
    "11111000", -- 5875 - 0x16f3  :  248 - 0xf8
    "11110000", -- 5876 - 0x16f4  :  240 - 0xf0
    "11100000", -- 5877 - 0x16f5  :  224 - 0xe0
    "00000000", -- 5878 - 0x16f6  :    0 - 0x0
    "00000000", -- 5879 - 0x16f7  :    0 - 0x0
    "11101100", -- 5880 - 0x16f8  :  236 - 0xec
    "11101100", -- 5881 - 0x16f9  :  236 - 0xec
    "11011000", -- 5882 - 0x16fa  :  216 - 0xd8
    "11111000", -- 5883 - 0x16fb  :  248 - 0xf8
    "11110000", -- 5884 - 0x16fc  :  240 - 0xf0
    "11100000", -- 5885 - 0x16fd  :  224 - 0xe0
    "00000000", -- 5886 - 0x16fe  :    0 - 0x0
    "00000000", -- 5887 - 0x16ff  :    0 - 0x0
    "00000000", -- 5888 - 0x1700  :    0 - 0x0 -- Background 0x70
    "00000100", -- 5889 - 0x1701  :    4 - 0x4
    "00000011", -- 5890 - 0x1702  :    3 - 0x3
    "00000000", -- 5891 - 0x1703  :    0 - 0x0
    "00000001", -- 5892 - 0x1704  :    1 - 0x1
    "00000111", -- 5893 - 0x1705  :    7 - 0x7
    "00001111", -- 5894 - 0x1706  :   15 - 0xf
    "00001100", -- 5895 - 0x1707  :   12 - 0xc
    "00000000", -- 5896 - 0x1708  :    0 - 0x0
    "00000000", -- 5897 - 0x1709  :    0 - 0x0
    "00000000", -- 5898 - 0x170a  :    0 - 0x0
    "00000000", -- 5899 - 0x170b  :    0 - 0x0
    "00000000", -- 5900 - 0x170c  :    0 - 0x0
    "00000000", -- 5901 - 0x170d  :    0 - 0x0
    "00000000", -- 5902 - 0x170e  :    0 - 0x0
    "00000000", -- 5903 - 0x170f  :    0 - 0x0
    "00000000", -- 5904 - 0x1710  :    0 - 0x0 -- Background 0x71
    "00000000", -- 5905 - 0x1711  :    0 - 0x0
    "11100000", -- 5906 - 0x1712  :  224 - 0xe0
    "10000000", -- 5907 - 0x1713  :  128 - 0x80
    "01000000", -- 5908 - 0x1714  :   64 - 0x40
    "11110000", -- 5909 - 0x1715  :  240 - 0xf0
    "10011000", -- 5910 - 0x1716  :  152 - 0x98
    "11111000", -- 5911 - 0x1717  :  248 - 0xf8
    "00000000", -- 5912 - 0x1718  :    0 - 0x0
    "00000000", -- 5913 - 0x1719  :    0 - 0x0
    "00000000", -- 5914 - 0x171a  :    0 - 0x0
    "00000000", -- 5915 - 0x171b  :    0 - 0x0
    "00000000", -- 5916 - 0x171c  :    0 - 0x0
    "00000000", -- 5917 - 0x171d  :    0 - 0x0
    "00000000", -- 5918 - 0x171e  :    0 - 0x0
    "00000000", -- 5919 - 0x171f  :    0 - 0x0
    "00011111", -- 5920 - 0x1720  :   31 - 0x1f -- Background 0x72
    "00010011", -- 5921 - 0x1721  :   19 - 0x13
    "00011111", -- 5922 - 0x1722  :   31 - 0x1f
    "00001111", -- 5923 - 0x1723  :   15 - 0xf
    "00001001", -- 5924 - 0x1724  :    9 - 0x9
    "00000111", -- 5925 - 0x1725  :    7 - 0x7
    "00000001", -- 5926 - 0x1726  :    1 - 0x1
    "00000000", -- 5927 - 0x1727  :    0 - 0x0
    "00000000", -- 5928 - 0x1728  :    0 - 0x0
    "00000000", -- 5929 - 0x1729  :    0 - 0x0
    "00000000", -- 5930 - 0x172a  :    0 - 0x0
    "00000000", -- 5931 - 0x172b  :    0 - 0x0
    "00000000", -- 5932 - 0x172c  :    0 - 0x0
    "00000000", -- 5933 - 0x172d  :    0 - 0x0
    "00000000", -- 5934 - 0x172e  :    0 - 0x0
    "00000000", -- 5935 - 0x172f  :    0 - 0x0
    "11100100", -- 5936 - 0x1730  :  228 - 0xe4 -- Background 0x73
    "00111100", -- 5937 - 0x1731  :   60 - 0x3c
    "11100100", -- 5938 - 0x1732  :  228 - 0xe4
    "00111000", -- 5939 - 0x1733  :   56 - 0x38
    "11111000", -- 5940 - 0x1734  :  248 - 0xf8
    "11110000", -- 5941 - 0x1735  :  240 - 0xf0
    "11000000", -- 5942 - 0x1736  :  192 - 0xc0
    "00000000", -- 5943 - 0x1737  :    0 - 0x0
    "00000000", -- 5944 - 0x1738  :    0 - 0x0
    "00000000", -- 5945 - 0x1739  :    0 - 0x0
    "00000000", -- 5946 - 0x173a  :    0 - 0x0
    "00000000", -- 5947 - 0x173b  :    0 - 0x0
    "00000000", -- 5948 - 0x173c  :    0 - 0x0
    "00000000", -- 5949 - 0x173d  :    0 - 0x0
    "00000000", -- 5950 - 0x173e  :    0 - 0x0
    "00000000", -- 5951 - 0x173f  :    0 - 0x0
    "00000000", -- 5952 - 0x1740  :    0 - 0x0 -- Background 0x74
    "00000000", -- 5953 - 0x1741  :    0 - 0x0
    "00000000", -- 5954 - 0x1742  :    0 - 0x0
    "00000000", -- 5955 - 0x1743  :    0 - 0x0
    "00000000", -- 5956 - 0x1744  :    0 - 0x0
    "00000000", -- 5957 - 0x1745  :    0 - 0x0
    "00000000", -- 5958 - 0x1746  :    0 - 0x0
    "00000000", -- 5959 - 0x1747  :    0 - 0x0
    "00000000", -- 5960 - 0x1748  :    0 - 0x0
    "00000000", -- 5961 - 0x1749  :    0 - 0x0
    "00000000", -- 5962 - 0x174a  :    0 - 0x0
    "00000000", -- 5963 - 0x174b  :    0 - 0x0
    "00010001", -- 5964 - 0x174c  :   17 - 0x11
    "00010011", -- 5965 - 0x174d  :   19 - 0x13
    "00011111", -- 5966 - 0x174e  :   31 - 0x1f
    "00011111", -- 5967 - 0x174f  :   31 - 0x1f
    "00000000", -- 5968 - 0x1750  :    0 - 0x0 -- Background 0x75
    "00000000", -- 5969 - 0x1751  :    0 - 0x0
    "00000000", -- 5970 - 0x1752  :    0 - 0x0
    "00000000", -- 5971 - 0x1753  :    0 - 0x0
    "00000000", -- 5972 - 0x1754  :    0 - 0x0
    "00000000", -- 5973 - 0x1755  :    0 - 0x0
    "00000000", -- 5974 - 0x1756  :    0 - 0x0
    "00000000", -- 5975 - 0x1757  :    0 - 0x0
    "00000000", -- 5976 - 0x1758  :    0 - 0x0
    "00000000", -- 5977 - 0x1759  :    0 - 0x0
    "00000000", -- 5978 - 0x175a  :    0 - 0x0
    "10000000", -- 5979 - 0x175b  :  128 - 0x80
    "11000100", -- 5980 - 0x175c  :  196 - 0xc4
    "11100100", -- 5981 - 0x175d  :  228 - 0xe4
    "11111100", -- 5982 - 0x175e  :  252 - 0xfc
    "11111100", -- 5983 - 0x175f  :  252 - 0xfc
    "00000000", -- 5984 - 0x1760  :    0 - 0x0 -- Background 0x76
    "00000000", -- 5985 - 0x1761  :    0 - 0x0
    "00000000", -- 5986 - 0x1762  :    0 - 0x0
    "00000000", -- 5987 - 0x1763  :    0 - 0x0
    "00000000", -- 5988 - 0x1764  :    0 - 0x0
    "00000000", -- 5989 - 0x1765  :    0 - 0x0
    "00000000", -- 5990 - 0x1766  :    0 - 0x0
    "00000000", -- 5991 - 0x1767  :    0 - 0x0
    "00011111", -- 5992 - 0x1768  :   31 - 0x1f
    "00001110", -- 5993 - 0x1769  :   14 - 0xe
    "00000110", -- 5994 - 0x176a  :    6 - 0x6
    "00000010", -- 5995 - 0x176b  :    2 - 0x2
    "00000000", -- 5996 - 0x176c  :    0 - 0x0
    "00000000", -- 5997 - 0x176d  :    0 - 0x0
    "00000000", -- 5998 - 0x176e  :    0 - 0x0
    "00000000", -- 5999 - 0x176f  :    0 - 0x0
    "00000000", -- 6000 - 0x1770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 6001 - 0x1771  :    0 - 0x0
    "00000000", -- 6002 - 0x1772  :    0 - 0x0
    "00000000", -- 6003 - 0x1773  :    0 - 0x0
    "00000000", -- 6004 - 0x1774  :    0 - 0x0
    "00000000", -- 6005 - 0x1775  :    0 - 0x0
    "00000000", -- 6006 - 0x1776  :    0 - 0x0
    "00000000", -- 6007 - 0x1777  :    0 - 0x0
    "11111100", -- 6008 - 0x1778  :  252 - 0xfc
    "10111000", -- 6009 - 0x1779  :  184 - 0xb8
    "10110000", -- 6010 - 0x177a  :  176 - 0xb0
    "10100000", -- 6011 - 0x177b  :  160 - 0xa0
    "10000000", -- 6012 - 0x177c  :  128 - 0x80
    "00000000", -- 6013 - 0x177d  :    0 - 0x0
    "00000000", -- 6014 - 0x177e  :    0 - 0x0
    "00000000", -- 6015 - 0x177f  :    0 - 0x0
    "00000000", -- 6016 - 0x1780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 6017 - 0x1781  :    0 - 0x0
    "00000000", -- 6018 - 0x1782  :    0 - 0x0
    "00000000", -- 6019 - 0x1783  :    0 - 0x0
    "00000000", -- 6020 - 0x1784  :    0 - 0x0
    "00000000", -- 6021 - 0x1785  :    0 - 0x0
    "00000000", -- 6022 - 0x1786  :    0 - 0x0
    "00000000", -- 6023 - 0x1787  :    0 - 0x0
    "00000000", -- 6024 - 0x1788  :    0 - 0x0
    "00000000", -- 6025 - 0x1789  :    0 - 0x0
    "00000000", -- 6026 - 0x178a  :    0 - 0x0
    "00000001", -- 6027 - 0x178b  :    1 - 0x1
    "00000011", -- 6028 - 0x178c  :    3 - 0x3
    "00000110", -- 6029 - 0x178d  :    6 - 0x6
    "00000110", -- 6030 - 0x178e  :    6 - 0x6
    "00001111", -- 6031 - 0x178f  :   15 - 0xf
    "00000000", -- 6032 - 0x1790  :    0 - 0x0 -- Background 0x79
    "00000000", -- 6033 - 0x1791  :    0 - 0x0
    "00000000", -- 6034 - 0x1792  :    0 - 0x0
    "00000000", -- 6035 - 0x1793  :    0 - 0x0
    "00000000", -- 6036 - 0x1794  :    0 - 0x0
    "00000000", -- 6037 - 0x1795  :    0 - 0x0
    "00000000", -- 6038 - 0x1796  :    0 - 0x0
    "00000000", -- 6039 - 0x1797  :    0 - 0x0
    "00000000", -- 6040 - 0x1798  :    0 - 0x0
    "00011000", -- 6041 - 0x1799  :   24 - 0x18
    "11110100", -- 6042 - 0x179a  :  244 - 0xf4
    "11111000", -- 6043 - 0x179b  :  248 - 0xf8
    "00111000", -- 6044 - 0x179c  :   56 - 0x38
    "01111100", -- 6045 - 0x179d  :  124 - 0x7c
    "11111100", -- 6046 - 0x179e  :  252 - 0xfc
    "11111100", -- 6047 - 0x179f  :  252 - 0xfc
    "00000000", -- 6048 - 0x17a0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 6049 - 0x17a1  :    0 - 0x0
    "00000000", -- 6050 - 0x17a2  :    0 - 0x0
    "00000000", -- 6051 - 0x17a3  :    0 - 0x0
    "00000000", -- 6052 - 0x17a4  :    0 - 0x0
    "00000000", -- 6053 - 0x17a5  :    0 - 0x0
    "00000000", -- 6054 - 0x17a6  :    0 - 0x0
    "00000000", -- 6055 - 0x17a7  :    0 - 0x0
    "00001111", -- 6056 - 0x17a8  :   15 - 0xf
    "00011111", -- 6057 - 0x17a9  :   31 - 0x1f
    "00110000", -- 6058 - 0x17aa  :   48 - 0x30
    "00111000", -- 6059 - 0x17ab  :   56 - 0x38
    "00011101", -- 6060 - 0x17ac  :   29 - 0x1d
    "00000011", -- 6061 - 0x17ad  :    3 - 0x3
    "00000011", -- 6062 - 0x17ae  :    3 - 0x3
    "00000000", -- 6063 - 0x17af  :    0 - 0x0
    "00000000", -- 6064 - 0x17b0  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 6065 - 0x17b1  :    0 - 0x0
    "00000000", -- 6066 - 0x17b2  :    0 - 0x0
    "00000000", -- 6067 - 0x17b3  :    0 - 0x0
    "00000000", -- 6068 - 0x17b4  :    0 - 0x0
    "00000000", -- 6069 - 0x17b5  :    0 - 0x0
    "00000000", -- 6070 - 0x17b6  :    0 - 0x0
    "00000000", -- 6071 - 0x17b7  :    0 - 0x0
    "11111100", -- 6072 - 0x17b8  :  252 - 0xfc
    "11111100", -- 6073 - 0x17b9  :  252 - 0xfc
    "01111100", -- 6074 - 0x17ba  :  124 - 0x7c
    "10001110", -- 6075 - 0x17bb  :  142 - 0x8e
    "10000110", -- 6076 - 0x17bc  :  134 - 0x86
    "10011100", -- 6077 - 0x17bd  :  156 - 0x9c
    "01111000", -- 6078 - 0x17be  :  120 - 0x78
    "00000000", -- 6079 - 0x17bf  :    0 - 0x0
    "00000000", -- 6080 - 0x17c0  :    0 - 0x0 -- Background 0x7c
    "00000001", -- 6081 - 0x17c1  :    1 - 0x1
    "00000110", -- 6082 - 0x17c2  :    6 - 0x6
    "00000111", -- 6083 - 0x17c3  :    7 - 0x7
    "00000111", -- 6084 - 0x17c4  :    7 - 0x7
    "00000111", -- 6085 - 0x17c5  :    7 - 0x7
    "00000001", -- 6086 - 0x17c6  :    1 - 0x1
    "00000011", -- 6087 - 0x17c7  :    3 - 0x3
    "00000000", -- 6088 - 0x17c8  :    0 - 0x0
    "00000001", -- 6089 - 0x17c9  :    1 - 0x1
    "00000110", -- 6090 - 0x17ca  :    6 - 0x6
    "00000111", -- 6091 - 0x17cb  :    7 - 0x7
    "00000111", -- 6092 - 0x17cc  :    7 - 0x7
    "00000111", -- 6093 - 0x17cd  :    7 - 0x7
    "00000001", -- 6094 - 0x17ce  :    1 - 0x1
    "00000011", -- 6095 - 0x17cf  :    3 - 0x3
    "00000000", -- 6096 - 0x17d0  :    0 - 0x0 -- Background 0x7d
    "11000000", -- 6097 - 0x17d1  :  192 - 0xc0
    "00110000", -- 6098 - 0x17d2  :   48 - 0x30
    "11110000", -- 6099 - 0x17d3  :  240 - 0xf0
    "11110000", -- 6100 - 0x17d4  :  240 - 0xf0
    "11110000", -- 6101 - 0x17d5  :  240 - 0xf0
    "01000000", -- 6102 - 0x17d6  :   64 - 0x40
    "01000000", -- 6103 - 0x17d7  :   64 - 0x40
    "00000000", -- 6104 - 0x17d8  :    0 - 0x0
    "11000000", -- 6105 - 0x17d9  :  192 - 0xc0
    "00110000", -- 6106 - 0x17da  :   48 - 0x30
    "11110000", -- 6107 - 0x17db  :  240 - 0xf0
    "11110000", -- 6108 - 0x17dc  :  240 - 0xf0
    "11110000", -- 6109 - 0x17dd  :  240 - 0xf0
    "01000000", -- 6110 - 0x17de  :   64 - 0x40
    "01000000", -- 6111 - 0x17df  :   64 - 0x40
    "00000001", -- 6112 - 0x17e0  :    1 - 0x1 -- Background 0x7e
    "00000000", -- 6113 - 0x17e1  :    0 - 0x0
    "00000001", -- 6114 - 0x17e2  :    1 - 0x1
    "00000011", -- 6115 - 0x17e3  :    3 - 0x3
    "00000001", -- 6116 - 0x17e4  :    1 - 0x1
    "00000000", -- 6117 - 0x17e5  :    0 - 0x0
    "00000000", -- 6118 - 0x17e6  :    0 - 0x0
    "00000000", -- 6119 - 0x17e7  :    0 - 0x0
    "00000001", -- 6120 - 0x17e8  :    1 - 0x1
    "00000000", -- 6121 - 0x17e9  :    0 - 0x0
    "00000001", -- 6122 - 0x17ea  :    1 - 0x1
    "00000011", -- 6123 - 0x17eb  :    3 - 0x3
    "00000001", -- 6124 - 0x17ec  :    1 - 0x1
    "00000000", -- 6125 - 0x17ed  :    0 - 0x0
    "00000000", -- 6126 - 0x17ee  :    0 - 0x0
    "00000000", -- 6127 - 0x17ef  :    0 - 0x0
    "01000000", -- 6128 - 0x17f0  :   64 - 0x40 -- Background 0x7f
    "01000000", -- 6129 - 0x17f1  :   64 - 0x40
    "01000000", -- 6130 - 0x17f2  :   64 - 0x40
    "01000000", -- 6131 - 0x17f3  :   64 - 0x40
    "01000000", -- 6132 - 0x17f4  :   64 - 0x40
    "10000000", -- 6133 - 0x17f5  :  128 - 0x80
    "00000000", -- 6134 - 0x17f6  :    0 - 0x0
    "00000000", -- 6135 - 0x17f7  :    0 - 0x0
    "01000000", -- 6136 - 0x17f8  :   64 - 0x40
    "01000000", -- 6137 - 0x17f9  :   64 - 0x40
    "01000000", -- 6138 - 0x17fa  :   64 - 0x40
    "01000000", -- 6139 - 0x17fb  :   64 - 0x40
    "01000000", -- 6140 - 0x17fc  :   64 - 0x40
    "10000000", -- 6141 - 0x17fd  :  128 - 0x80
    "00000000", -- 6142 - 0x17fe  :    0 - 0x0
    "00000000", -- 6143 - 0x17ff  :    0 - 0x0
    "11111111", -- 6144 - 0x1800  :  255 - 0xff -- Background 0x80
    "11111111", -- 6145 - 0x1801  :  255 - 0xff
    "11111111", -- 6146 - 0x1802  :  255 - 0xff
    "11111111", -- 6147 - 0x1803  :  255 - 0xff
    "11000000", -- 6148 - 0x1804  :  192 - 0xc0
    "11000000", -- 6149 - 0x1805  :  192 - 0xc0
    "11000000", -- 6150 - 0x1806  :  192 - 0xc0
    "11000111", -- 6151 - 0x1807  :  199 - 0xc7
    "00000000", -- 6152 - 0x1808  :    0 - 0x0
    "00000000", -- 6153 - 0x1809  :    0 - 0x0
    "00000000", -- 6154 - 0x180a  :    0 - 0x0
    "00000000", -- 6155 - 0x180b  :    0 - 0x0
    "00000000", -- 6156 - 0x180c  :    0 - 0x0
    "00011111", -- 6157 - 0x180d  :   31 - 0x1f
    "00010000", -- 6158 - 0x180e  :   16 - 0x10
    "00010111", -- 6159 - 0x180f  :   23 - 0x17
    "11111111", -- 6160 - 0x1810  :  255 - 0xff -- Background 0x81
    "11111111", -- 6161 - 0x1811  :  255 - 0xff
    "11111111", -- 6162 - 0x1812  :  255 - 0xff
    "11111111", -- 6163 - 0x1813  :  255 - 0xff
    "00000000", -- 6164 - 0x1814  :    0 - 0x0
    "00000000", -- 6165 - 0x1815  :    0 - 0x0
    "00000000", -- 6166 - 0x1816  :    0 - 0x0
    "11111111", -- 6167 - 0x1817  :  255 - 0xff
    "00000000", -- 6168 - 0x1818  :    0 - 0x0
    "00000000", -- 6169 - 0x1819  :    0 - 0x0
    "00000000", -- 6170 - 0x181a  :    0 - 0x0
    "00000000", -- 6171 - 0x181b  :    0 - 0x0
    "00000000", -- 6172 - 0x181c  :    0 - 0x0
    "11111111", -- 6173 - 0x181d  :  255 - 0xff
    "00000000", -- 6174 - 0x181e  :    0 - 0x0
    "11111111", -- 6175 - 0x181f  :  255 - 0xff
    "11111111", -- 6176 - 0x1820  :  255 - 0xff -- Background 0x82
    "11111111", -- 6177 - 0x1821  :  255 - 0xff
    "11111111", -- 6178 - 0x1822  :  255 - 0xff
    "11111111", -- 6179 - 0x1823  :  255 - 0xff
    "01111111", -- 6180 - 0x1824  :  127 - 0x7f
    "00111111", -- 6181 - 0x1825  :   63 - 0x3f
    "00011111", -- 6182 - 0x1826  :   31 - 0x1f
    "11001111", -- 6183 - 0x1827  :  207 - 0xcf
    "00000000", -- 6184 - 0x1828  :    0 - 0x0
    "00000000", -- 6185 - 0x1829  :    0 - 0x0
    "00000000", -- 6186 - 0x182a  :    0 - 0x0
    "00000000", -- 6187 - 0x182b  :    0 - 0x0
    "00000000", -- 6188 - 0x182c  :    0 - 0x0
    "10000000", -- 6189 - 0x182d  :  128 - 0x80
    "00000000", -- 6190 - 0x182e  :    0 - 0x0
    "11000000", -- 6191 - 0x182f  :  192 - 0xc0
    "11111111", -- 6192 - 0x1830  :  255 - 0xff -- Background 0x83
    "11111111", -- 6193 - 0x1831  :  255 - 0xff
    "11111111", -- 6194 - 0x1832  :  255 - 0xff
    "11110111", -- 6195 - 0x1833  :  247 - 0xf7
    "11110111", -- 6196 - 0x1834  :  247 - 0xf7
    "11100010", -- 6197 - 0x1835  :  226 - 0xe2
    "11100000", -- 6198 - 0x1836  :  224 - 0xe0
    "11000110", -- 6199 - 0x1837  :  198 - 0xc6
    "00000000", -- 6200 - 0x1838  :    0 - 0x0
    "00000000", -- 6201 - 0x1839  :    0 - 0x0
    "00000000", -- 6202 - 0x183a  :    0 - 0x0
    "00000000", -- 6203 - 0x183b  :    0 - 0x0
    "00000000", -- 6204 - 0x183c  :    0 - 0x0
    "00001000", -- 6205 - 0x183d  :    8 - 0x8
    "00001000", -- 6206 - 0x183e  :    8 - 0x8
    "00010110", -- 6207 - 0x183f  :   22 - 0x16
    "11111111", -- 6208 - 0x1840  :  255 - 0xff -- Background 0x84
    "11111111", -- 6209 - 0x1841  :  255 - 0xff
    "11111111", -- 6210 - 0x1842  :  255 - 0xff
    "11111111", -- 6211 - 0x1843  :  255 - 0xff
    "10111111", -- 6212 - 0x1844  :  191 - 0xbf
    "10111111", -- 6213 - 0x1845  :  191 - 0xbf
    "00011111", -- 6214 - 0x1846  :   31 - 0x1f
    "00011111", -- 6215 - 0x1847  :   31 - 0x1f
    "00000000", -- 6216 - 0x1848  :    0 - 0x0
    "00000000", -- 6217 - 0x1849  :    0 - 0x0
    "00000000", -- 6218 - 0x184a  :    0 - 0x0
    "00000000", -- 6219 - 0x184b  :    0 - 0x0
    "00000000", -- 6220 - 0x184c  :    0 - 0x0
    "00000000", -- 6221 - 0x184d  :    0 - 0x0
    "01000000", -- 6222 - 0x184e  :   64 - 0x40
    "11000000", -- 6223 - 0x184f  :  192 - 0xc0
    "11111111", -- 6224 - 0x1850  :  255 - 0xff -- Background 0x85
    "11111111", -- 6225 - 0x1851  :  255 - 0xff
    "11111111", -- 6226 - 0x1852  :  255 - 0xff
    "11111111", -- 6227 - 0x1853  :  255 - 0xff
    "11111110", -- 6228 - 0x1854  :  254 - 0xfe
    "11111000", -- 6229 - 0x1855  :  248 - 0xf8
    "11100000", -- 6230 - 0x1856  :  224 - 0xe0
    "11000000", -- 6231 - 0x1857  :  192 - 0xc0
    "00000000", -- 6232 - 0x1858  :    0 - 0x0
    "00000000", -- 6233 - 0x1859  :    0 - 0x0
    "00000000", -- 6234 - 0x185a  :    0 - 0x0
    "00000000", -- 6235 - 0x185b  :    0 - 0x0
    "00000000", -- 6236 - 0x185c  :    0 - 0x0
    "00000001", -- 6237 - 0x185d  :    1 - 0x1
    "00000111", -- 6238 - 0x185e  :    7 - 0x7
    "00001100", -- 6239 - 0x185f  :   12 - 0xc
    "11111111", -- 6240 - 0x1860  :  255 - 0xff -- Background 0x86
    "11111111", -- 6241 - 0x1861  :  255 - 0xff
    "11111111", -- 6242 - 0x1862  :  255 - 0xff
    "11111111", -- 6243 - 0x1863  :  255 - 0xff
    "00000111", -- 6244 - 0x1864  :    7 - 0x7
    "00000000", -- 6245 - 0x1865  :    0 - 0x0
    "00111111", -- 6246 - 0x1866  :   63 - 0x3f
    "11111111", -- 6247 - 0x1867  :  255 - 0xff
    "00000000", -- 6248 - 0x1868  :    0 - 0x0
    "00000000", -- 6249 - 0x1869  :    0 - 0x0
    "00000000", -- 6250 - 0x186a  :    0 - 0x0
    "00000000", -- 6251 - 0x186b  :    0 - 0x0
    "00000000", -- 6252 - 0x186c  :    0 - 0x0
    "11000000", -- 6253 - 0x186d  :  192 - 0xc0
    "00111111", -- 6254 - 0x186e  :   63 - 0x3f
    "11111111", -- 6255 - 0x186f  :  255 - 0xff
    "11111111", -- 6256 - 0x1870  :  255 - 0xff -- Background 0x87
    "11111111", -- 6257 - 0x1871  :  255 - 0xff
    "11111111", -- 6258 - 0x1872  :  255 - 0xff
    "11111111", -- 6259 - 0x1873  :  255 - 0xff
    "11111111", -- 6260 - 0x1874  :  255 - 0xff
    "11111111", -- 6261 - 0x1875  :  255 - 0xff
    "00111111", -- 6262 - 0x1876  :   63 - 0x3f
    "11001111", -- 6263 - 0x1877  :  207 - 0xcf
    "00000000", -- 6264 - 0x1878  :    0 - 0x0
    "00000000", -- 6265 - 0x1879  :    0 - 0x0
    "00000000", -- 6266 - 0x187a  :    0 - 0x0
    "00000000", -- 6267 - 0x187b  :    0 - 0x0
    "00000000", -- 6268 - 0x187c  :    0 - 0x0
    "00000000", -- 6269 - 0x187d  :    0 - 0x0
    "00000000", -- 6270 - 0x187e  :    0 - 0x0
    "11000000", -- 6271 - 0x187f  :  192 - 0xc0
    "11111111", -- 6272 - 0x1880  :  255 - 0xff -- Background 0x88
    "11111111", -- 6273 - 0x1881  :  255 - 0xff
    "11111111", -- 6274 - 0x1882  :  255 - 0xff
    "11111111", -- 6275 - 0x1883  :  255 - 0xff
    "11111111", -- 6276 - 0x1884  :  255 - 0xff
    "11111111", -- 6277 - 0x1885  :  255 - 0xff
    "11111111", -- 6278 - 0x1886  :  255 - 0xff
    "11111111", -- 6279 - 0x1887  :  255 - 0xff
    "00000000", -- 6280 - 0x1888  :    0 - 0x0
    "00000000", -- 6281 - 0x1889  :    0 - 0x0
    "00000000", -- 6282 - 0x188a  :    0 - 0x0
    "00000000", -- 6283 - 0x188b  :    0 - 0x0
    "00000000", -- 6284 - 0x188c  :    0 - 0x0
    "00000000", -- 6285 - 0x188d  :    0 - 0x0
    "00000000", -- 6286 - 0x188e  :    0 - 0x0
    "00000000", -- 6287 - 0x188f  :    0 - 0x0
    "11111111", -- 6288 - 0x1890  :  255 - 0xff -- Background 0x89
    "11111111", -- 6289 - 0x1891  :  255 - 0xff
    "11111111", -- 6290 - 0x1892  :  255 - 0xff
    "01110111", -- 6291 - 0x1893  :  119 - 0x77
    "00010011", -- 6292 - 0x1894  :   19 - 0x13
    "00000001", -- 6293 - 0x1895  :    1 - 0x1
    "00010000", -- 6294 - 0x1896  :   16 - 0x10
    "00011000", -- 6295 - 0x1897  :   24 - 0x18
    "00000000", -- 6296 - 0x1898  :    0 - 0x0
    "00000000", -- 6297 - 0x1899  :    0 - 0x0
    "00000000", -- 6298 - 0x189a  :    0 - 0x0
    "00000000", -- 6299 - 0x189b  :    0 - 0x0
    "00000000", -- 6300 - 0x189c  :    0 - 0x0
    "01000100", -- 6301 - 0x189d  :   68 - 0x44
    "01010110", -- 6302 - 0x189e  :   86 - 0x56
    "01011011", -- 6303 - 0x189f  :   91 - 0x5b
    "11111111", -- 6304 - 0x18a0  :  255 - 0xff -- Background 0x8a
    "11111111", -- 6305 - 0x18a1  :  255 - 0xff
    "11111111", -- 6306 - 0x18a2  :  255 - 0xff
    "11111111", -- 6307 - 0x18a3  :  255 - 0xff
    "11111111", -- 6308 - 0x18a4  :  255 - 0xff
    "11111111", -- 6309 - 0x18a5  :  255 - 0xff
    "11111111", -- 6310 - 0x18a6  :  255 - 0xff
    "01111111", -- 6311 - 0x18a7  :  127 - 0x7f
    "00000000", -- 6312 - 0x18a8  :    0 - 0x0
    "00000000", -- 6313 - 0x18a9  :    0 - 0x0
    "00000000", -- 6314 - 0x18aa  :    0 - 0x0
    "00000000", -- 6315 - 0x18ab  :    0 - 0x0
    "00000000", -- 6316 - 0x18ac  :    0 - 0x0
    "00000000", -- 6317 - 0x18ad  :    0 - 0x0
    "00000000", -- 6318 - 0x18ae  :    0 - 0x0
    "00000000", -- 6319 - 0x18af  :    0 - 0x0
    "11111111", -- 6320 - 0x18b0  :  255 - 0xff -- Background 0x8b
    "11111111", -- 6321 - 0x18b1  :  255 - 0xff
    "11111111", -- 6322 - 0x18b2  :  255 - 0xff
    "11110111", -- 6323 - 0x18b3  :  247 - 0xf7
    "11100101", -- 6324 - 0x18b4  :  229 - 0xe5
    "11000001", -- 6325 - 0x18b5  :  193 - 0xc1
    "10000100", -- 6326 - 0x18b6  :  132 - 0x84
    "00001100", -- 6327 - 0x18b7  :   12 - 0xc
    "00000000", -- 6328 - 0x18b8  :    0 - 0x0
    "00000000", -- 6329 - 0x18b9  :    0 - 0x0
    "00000000", -- 6330 - 0x18ba  :    0 - 0x0
    "00000000", -- 6331 - 0x18bb  :    0 - 0x0
    "00000000", -- 6332 - 0x18bc  :    0 - 0x0
    "00010000", -- 6333 - 0x18bd  :   16 - 0x10
    "00110100", -- 6334 - 0x18be  :   52 - 0x34
    "01101101", -- 6335 - 0x18bf  :  109 - 0x6d
    "11111111", -- 6336 - 0x18c0  :  255 - 0xff -- Background 0x8c
    "11111111", -- 6337 - 0x18c1  :  255 - 0xff
    "11111111", -- 6338 - 0x18c2  :  255 - 0xff
    "11111111", -- 6339 - 0x18c3  :  255 - 0xff
    "11111111", -- 6340 - 0x18c4  :  255 - 0xff
    "01111111", -- 6341 - 0x18c5  :  127 - 0x7f
    "01111110", -- 6342 - 0x18c6  :  126 - 0x7e
    "01111110", -- 6343 - 0x18c7  :  126 - 0x7e
    "00000000", -- 6344 - 0x18c8  :    0 - 0x0
    "00000000", -- 6345 - 0x18c9  :    0 - 0x0
    "00000000", -- 6346 - 0x18ca  :    0 - 0x0
    "00000000", -- 6347 - 0x18cb  :    0 - 0x0
    "00000000", -- 6348 - 0x18cc  :    0 - 0x0
    "00000000", -- 6349 - 0x18cd  :    0 - 0x0
    "00000000", -- 6350 - 0x18ce  :    0 - 0x0
    "00000000", -- 6351 - 0x18cf  :    0 - 0x0
    "11111111", -- 6352 - 0x18d0  :  255 - 0xff -- Background 0x8d
    "11111111", -- 6353 - 0x18d1  :  255 - 0xff
    "10111111", -- 6354 - 0x18d2  :  191 - 0xbf
    "10110111", -- 6355 - 0x18d3  :  183 - 0xb7
    "00010111", -- 6356 - 0x18d4  :   23 - 0x17
    "00000011", -- 6357 - 0x18d5  :    3 - 0x3
    "00100011", -- 6358 - 0x18d6  :   35 - 0x23
    "00100001", -- 6359 - 0x18d7  :   33 - 0x21
    "00000000", -- 6360 - 0x18d8  :    0 - 0x0
    "00000000", -- 6361 - 0x18d9  :    0 - 0x0
    "00000000", -- 6362 - 0x18da  :    0 - 0x0
    "00000000", -- 6363 - 0x18db  :    0 - 0x0
    "01000000", -- 6364 - 0x18dc  :   64 - 0x40
    "01001000", -- 6365 - 0x18dd  :   72 - 0x48
    "10101000", -- 6366 - 0x18de  :  168 - 0xa8
    "10101100", -- 6367 - 0x18df  :  172 - 0xac
    "11111111", -- 6368 - 0x18e0  :  255 - 0xff -- Background 0x8e
    "11111111", -- 6369 - 0x18e1  :  255 - 0xff
    "11111011", -- 6370 - 0x18e2  :  251 - 0xfb
    "11111001", -- 6371 - 0x18e3  :  249 - 0xf9
    "11111000", -- 6372 - 0x18e4  :  248 - 0xf8
    "11111000", -- 6373 - 0x18e5  :  248 - 0xf8
    "11111000", -- 6374 - 0x18e6  :  248 - 0xf8
    "11111000", -- 6375 - 0x18e7  :  248 - 0xf8
    "00000000", -- 6376 - 0x18e8  :    0 - 0x0
    "00000000", -- 6377 - 0x18e9  :    0 - 0x0
    "00000000", -- 6378 - 0x18ea  :    0 - 0x0
    "00000000", -- 6379 - 0x18eb  :    0 - 0x0
    "00000010", -- 6380 - 0x18ec  :    2 - 0x2
    "00000010", -- 6381 - 0x18ed  :    2 - 0x2
    "00000010", -- 6382 - 0x18ee  :    2 - 0x2
    "00000010", -- 6383 - 0x18ef  :    2 - 0x2
    "11111111", -- 6384 - 0x18f0  :  255 - 0xff -- Background 0x8f
    "11111111", -- 6385 - 0x18f1  :  255 - 0xff
    "01111000", -- 6386 - 0x18f2  :  120 - 0x78
    "00111000", -- 6387 - 0x18f3  :   56 - 0x38
    "00011000", -- 6388 - 0x18f4  :   24 - 0x18
    "00001000", -- 6389 - 0x18f5  :    8 - 0x8
    "10000000", -- 6390 - 0x18f6  :  128 - 0x80
    "11000000", -- 6391 - 0x18f7  :  192 - 0xc0
    "00000000", -- 6392 - 0x18f8  :    0 - 0x0
    "00000000", -- 6393 - 0x18f9  :    0 - 0x0
    "00000000", -- 6394 - 0x18fa  :    0 - 0x0
    "00000011", -- 6395 - 0x18fb  :    3 - 0x3
    "01000011", -- 6396 - 0x18fc  :   67 - 0x43
    "01100010", -- 6397 - 0x18fd  :   98 - 0x62
    "10110010", -- 6398 - 0x18fe  :  178 - 0xb2
    "11011010", -- 6399 - 0x18ff  :  218 - 0xda
    "11111111", -- 6400 - 0x1900  :  255 - 0xff -- Background 0x90
    "11111111", -- 6401 - 0x1901  :  255 - 0xff
    "00000001", -- 6402 - 0x1902  :    1 - 0x1
    "00000001", -- 6403 - 0x1903  :    1 - 0x1
    "00000001", -- 6404 - 0x1904  :    1 - 0x1
    "00000000", -- 6405 - 0x1905  :    0 - 0x0
    "11111111", -- 6406 - 0x1906  :  255 - 0xff
    "11111111", -- 6407 - 0x1907  :  255 - 0xff
    "00000000", -- 6408 - 0x1908  :    0 - 0x0
    "00000000", -- 6409 - 0x1909  :    0 - 0x0
    "00000000", -- 6410 - 0x190a  :    0 - 0x0
    "11111100", -- 6411 - 0x190b  :  252 - 0xfc
    "11111100", -- 6412 - 0x190c  :  252 - 0xfc
    "00000000", -- 6413 - 0x190d  :    0 - 0x0
    "11111111", -- 6414 - 0x190e  :  255 - 0xff
    "11111111", -- 6415 - 0x190f  :  255 - 0xff
    "11111111", -- 6416 - 0x1910  :  255 - 0xff -- Background 0x91
    "11111111", -- 6417 - 0x1911  :  255 - 0xff
    "11111111", -- 6418 - 0x1912  :  255 - 0xff
    "11111111", -- 6419 - 0x1913  :  255 - 0xff
    "11111111", -- 6420 - 0x1914  :  255 - 0xff
    "11111111", -- 6421 - 0x1915  :  255 - 0xff
    "01111111", -- 6422 - 0x1916  :  127 - 0x7f
    "00111111", -- 6423 - 0x1917  :   63 - 0x3f
    "00000000", -- 6424 - 0x1918  :    0 - 0x0
    "00000000", -- 6425 - 0x1919  :    0 - 0x0
    "00000000", -- 6426 - 0x191a  :    0 - 0x0
    "00000000", -- 6427 - 0x191b  :    0 - 0x0
    "00000000", -- 6428 - 0x191c  :    0 - 0x0
    "00000000", -- 6429 - 0x191d  :    0 - 0x0
    "00000000", -- 6430 - 0x191e  :    0 - 0x0
    "00000000", -- 6431 - 0x191f  :    0 - 0x0
    "11000111", -- 6432 - 0x1920  :  199 - 0xc7 -- Background 0x92
    "11000111", -- 6433 - 0x1921  :  199 - 0xc7
    "11000111", -- 6434 - 0x1922  :  199 - 0xc7
    "11000111", -- 6435 - 0x1923  :  199 - 0xc7
    "11000111", -- 6436 - 0x1924  :  199 - 0xc7
    "11000111", -- 6437 - 0x1925  :  199 - 0xc7
    "11000111", -- 6438 - 0x1926  :  199 - 0xc7
    "11000111", -- 6439 - 0x1927  :  199 - 0xc7
    "00010111", -- 6440 - 0x1928  :   23 - 0x17
    "00010111", -- 6441 - 0x1929  :   23 - 0x17
    "00010111", -- 6442 - 0x192a  :   23 - 0x17
    "00010111", -- 6443 - 0x192b  :   23 - 0x17
    "00010111", -- 6444 - 0x192c  :   23 - 0x17
    "00010111", -- 6445 - 0x192d  :   23 - 0x17
    "00010111", -- 6446 - 0x192e  :   23 - 0x17
    "00010111", -- 6447 - 0x192f  :   23 - 0x17
    "11111111", -- 6448 - 0x1930  :  255 - 0xff -- Background 0x93
    "11111111", -- 6449 - 0x1931  :  255 - 0xff
    "11111111", -- 6450 - 0x1932  :  255 - 0xff
    "11111111", -- 6451 - 0x1933  :  255 - 0xff
    "11111001", -- 6452 - 0x1934  :  249 - 0xf9
    "11111001", -- 6453 - 0x1935  :  249 - 0xf9
    "11111111", -- 6454 - 0x1936  :  255 - 0xff
    "11111111", -- 6455 - 0x1937  :  255 - 0xff
    "11111111", -- 6456 - 0x1938  :  255 - 0xff
    "11111111", -- 6457 - 0x1939  :  255 - 0xff
    "11111111", -- 6458 - 0x193a  :  255 - 0xff
    "11111111", -- 6459 - 0x193b  :  255 - 0xff
    "11111001", -- 6460 - 0x193c  :  249 - 0xf9
    "11111001", -- 6461 - 0x193d  :  249 - 0xf9
    "11111111", -- 6462 - 0x193e  :  255 - 0xff
    "11111111", -- 6463 - 0x193f  :  255 - 0xff
    "11110111", -- 6464 - 0x1940  :  247 - 0xf7 -- Background 0x94
    "11111011", -- 6465 - 0x1941  :  251 - 0xfb
    "11111011", -- 6466 - 0x1942  :  251 - 0xfb
    "11111101", -- 6467 - 0x1943  :  253 - 0xfd
    "11111100", -- 6468 - 0x1944  :  252 - 0xfc
    "11111100", -- 6469 - 0x1945  :  252 - 0xfc
    "01111100", -- 6470 - 0x1946  :  124 - 0x7c
    "01111100", -- 6471 - 0x1947  :  124 - 0x7c
    "11110000", -- 6472 - 0x1948  :  240 - 0xf0
    "11111000", -- 6473 - 0x1949  :  248 - 0xf8
    "11111000", -- 6474 - 0x194a  :  248 - 0xf8
    "11111100", -- 6475 - 0x194b  :  252 - 0xfc
    "11111100", -- 6476 - 0x194c  :  252 - 0xfc
    "11111100", -- 6477 - 0x194d  :  252 - 0xfc
    "01111100", -- 6478 - 0x194e  :  124 - 0x7c
    "01111100", -- 6479 - 0x194f  :  124 - 0x7c
    "11000111", -- 6480 - 0x1950  :  199 - 0xc7 -- Background 0x95
    "10001111", -- 6481 - 0x1951  :  143 - 0x8f
    "10001111", -- 6482 - 0x1952  :  143 - 0x8f
    "00011111", -- 6483 - 0x1953  :   31 - 0x1f
    "00011111", -- 6484 - 0x1954  :   31 - 0x1f
    "00111111", -- 6485 - 0x1955  :   63 - 0x3f
    "00111111", -- 6486 - 0x1956  :   63 - 0x3f
    "01111111", -- 6487 - 0x1957  :  127 - 0x7f
    "00010111", -- 6488 - 0x1958  :   23 - 0x17
    "00101111", -- 6489 - 0x1959  :   47 - 0x2f
    "00101111", -- 6490 - 0x195a  :   47 - 0x2f
    "01011111", -- 6491 - 0x195b  :   95 - 0x5f
    "01011111", -- 6492 - 0x195c  :   95 - 0x5f
    "10111111", -- 6493 - 0x195d  :  191 - 0xbf
    "10111111", -- 6494 - 0x195e  :  191 - 0xbf
    "01111111", -- 6495 - 0x195f  :  127 - 0x7f
    "00001111", -- 6496 - 0x1960  :   15 - 0xf -- Background 0x96
    "00001111", -- 6497 - 0x1961  :   15 - 0xf
    "10000111", -- 6498 - 0x1962  :  135 - 0x87
    "10000111", -- 6499 - 0x1963  :  135 - 0x87
    "11000010", -- 6500 - 0x1964  :  194 - 0xc2
    "11000010", -- 6501 - 0x1965  :  194 - 0xc2
    "11100000", -- 6502 - 0x1966  :  224 - 0xe0
    "11100000", -- 6503 - 0x1967  :  224 - 0xe0
    "01100000", -- 6504 - 0x1968  :   96 - 0x60
    "01100000", -- 6505 - 0x1969  :   96 - 0x60
    "10110000", -- 6506 - 0x196a  :  176 - 0xb0
    "10110000", -- 6507 - 0x196b  :  176 - 0xb0
    "11011000", -- 6508 - 0x196c  :  216 - 0xd8
    "11011000", -- 6509 - 0x196d  :  216 - 0xd8
    "11101100", -- 6510 - 0x196e  :  236 - 0xec
    "11101100", -- 6511 - 0x196f  :  236 - 0xec
    "10000011", -- 6512 - 0x1970  :  131 - 0x83 -- Background 0x97
    "10001111", -- 6513 - 0x1971  :  143 - 0x8f
    "00001111", -- 6514 - 0x1972  :   15 - 0xf
    "00011111", -- 6515 - 0x1973  :   31 - 0x1f
    "00011111", -- 6516 - 0x1974  :   31 - 0x1f
    "00111111", -- 6517 - 0x1975  :   63 - 0x3f
    "00111111", -- 6518 - 0x1976  :   63 - 0x3f
    "00111111", -- 6519 - 0x1977  :   63 - 0x3f
    "00110011", -- 6520 - 0x1978  :   51 - 0x33
    "00101111", -- 6521 - 0x1979  :   47 - 0x2f
    "01101111", -- 6522 - 0x197a  :  111 - 0x6f
    "01011111", -- 6523 - 0x197b  :   95 - 0x5f
    "11011111", -- 6524 - 0x197c  :  223 - 0xdf
    "10111111", -- 6525 - 0x197d  :  191 - 0xbf
    "10111111", -- 6526 - 0x197e  :  191 - 0xbf
    "10111111", -- 6527 - 0x197f  :  191 - 0xbf
    "11111111", -- 6528 - 0x1980  :  255 - 0xff -- Background 0x98
    "11111111", -- 6529 - 0x1981  :  255 - 0xff
    "11111111", -- 6530 - 0x1982  :  255 - 0xff
    "11111110", -- 6531 - 0x1983  :  254 - 0xfe
    "11111001", -- 6532 - 0x1984  :  249 - 0xf9
    "11100111", -- 6533 - 0x1985  :  231 - 0xe7
    "11111100", -- 6534 - 0x1986  :  252 - 0xfc
    "11110000", -- 6535 - 0x1987  :  240 - 0xf0
    "11111111", -- 6536 - 0x1988  :  255 - 0xff
    "11111111", -- 6537 - 0x1989  :  255 - 0xff
    "11111111", -- 6538 - 0x198a  :  255 - 0xff
    "11111110", -- 6539 - 0x198b  :  254 - 0xfe
    "11111001", -- 6540 - 0x198c  :  249 - 0xf9
    "11100111", -- 6541 - 0x198d  :  231 - 0xe7
    "11111100", -- 6542 - 0x198e  :  252 - 0xfc
    "11110011", -- 6543 - 0x198f  :  243 - 0xf3
    "11110111", -- 6544 - 0x1990  :  247 - 0xf7 -- Background 0x99
    "11111011", -- 6545 - 0x1991  :  251 - 0xfb
    "11111011", -- 6546 - 0x1992  :  251 - 0xfb
    "01110011", -- 6547 - 0x1993  :  115 - 0x73
    "11000001", -- 6548 - 0x1994  :  193 - 0xc1
    "00000011", -- 6549 - 0x1995  :    3 - 0x3
    "00001111", -- 6550 - 0x1996  :   15 - 0xf
    "00111111", -- 6551 - 0x1997  :   63 - 0x3f
    "11110000", -- 6552 - 0x1998  :  240 - 0xf0
    "11111000", -- 6553 - 0x1999  :  248 - 0xf8
    "11111000", -- 6554 - 0x199a  :  248 - 0xf8
    "01110000", -- 6555 - 0x199b  :  112 - 0x70
    "11001100", -- 6556 - 0x199c  :  204 - 0xcc
    "00110000", -- 6557 - 0x199d  :   48 - 0x30
    "11000000", -- 6558 - 0x199e  :  192 - 0xc0
    "00000000", -- 6559 - 0x199f  :    0 - 0x0
    "11111111", -- 6560 - 0x19a0  :  255 - 0xff -- Background 0x9a
    "11111111", -- 6561 - 0x19a1  :  255 - 0xff
    "11111111", -- 6562 - 0x19a2  :  255 - 0xff
    "10000000", -- 6563 - 0x19a3  :  128 - 0x80
    "10000000", -- 6564 - 0x19a4  :  128 - 0x80
    "10000000", -- 6565 - 0x19a5  :  128 - 0x80
    "10001111", -- 6566 - 0x19a6  :  143 - 0x8f
    "10001111", -- 6567 - 0x19a7  :  143 - 0x8f
    "00000000", -- 6568 - 0x19a8  :    0 - 0x0
    "00000000", -- 6569 - 0x19a9  :    0 - 0x0
    "00000000", -- 6570 - 0x19aa  :    0 - 0x0
    "00000000", -- 6571 - 0x19ab  :    0 - 0x0
    "00111111", -- 6572 - 0x19ac  :   63 - 0x3f
    "00100000", -- 6573 - 0x19ad  :   32 - 0x20
    "00101111", -- 6574 - 0x19ae  :   47 - 0x2f
    "00101111", -- 6575 - 0x19af  :   47 - 0x2f
    "11111111", -- 6576 - 0x19b0  :  255 - 0xff -- Background 0x9b
    "11111111", -- 6577 - 0x19b1  :  255 - 0xff
    "11111111", -- 6578 - 0x19b2  :  255 - 0xff
    "00001111", -- 6579 - 0x19b3  :   15 - 0xf
    "00001111", -- 6580 - 0x19b4  :   15 - 0xf
    "00000111", -- 6581 - 0x19b5  :    7 - 0x7
    "11110111", -- 6582 - 0x19b6  :  247 - 0xf7
    "11110001", -- 6583 - 0x19b7  :  241 - 0xf1
    "00000000", -- 6584 - 0x19b8  :    0 - 0x0
    "00000000", -- 6585 - 0x19b9  :    0 - 0x0
    "00000000", -- 6586 - 0x19ba  :    0 - 0x0
    "00000000", -- 6587 - 0x19bb  :    0 - 0x0
    "11100000", -- 6588 - 0x19bc  :  224 - 0xe0
    "00000000", -- 6589 - 0x19bd  :    0 - 0x0
    "11110000", -- 6590 - 0x19be  :  240 - 0xf0
    "11110000", -- 6591 - 0x19bf  :  240 - 0xf0
    "00011100", -- 6592 - 0x19c0  :   28 - 0x1c -- Background 0x9c
    "00011110", -- 6593 - 0x19c1  :   30 - 0x1e
    "00011111", -- 6594 - 0x19c2  :   31 - 0x1f
    "00011111", -- 6595 - 0x19c3  :   31 - 0x1f
    "00011111", -- 6596 - 0x19c4  :   31 - 0x1f
    "00011111", -- 6597 - 0x19c5  :   31 - 0x1f
    "00011111", -- 6598 - 0x19c6  :   31 - 0x1f
    "00011111", -- 6599 - 0x19c7  :   31 - 0x1f
    "01011101", -- 6600 - 0x19c8  :   93 - 0x5d
    "01011110", -- 6601 - 0x19c9  :   94 - 0x5e
    "01011111", -- 6602 - 0x19ca  :   95 - 0x5f
    "01011111", -- 6603 - 0x19cb  :   95 - 0x5f
    "01011111", -- 6604 - 0x19cc  :   95 - 0x5f
    "01011111", -- 6605 - 0x19cd  :   95 - 0x5f
    "01011111", -- 6606 - 0x19ce  :   95 - 0x5f
    "01011111", -- 6607 - 0x19cf  :   95 - 0x5f
    "00111110", -- 6608 - 0x19d0  :   62 - 0x3e -- Background 0x9d
    "00011100", -- 6609 - 0x19d1  :   28 - 0x1c
    "00001000", -- 6610 - 0x19d2  :    8 - 0x8
    "10000000", -- 6611 - 0x19d3  :  128 - 0x80
    "11000001", -- 6612 - 0x19d4  :  193 - 0xc1
    "11100011", -- 6613 - 0x19d5  :  227 - 0xe3
    "11110111", -- 6614 - 0x19d6  :  247 - 0xf7
    "11111111", -- 6615 - 0x19d7  :  255 - 0xff
    "10000000", -- 6616 - 0x19d8  :  128 - 0x80
    "11000001", -- 6617 - 0x19d9  :  193 - 0xc1
    "01100011", -- 6618 - 0x19da  :   99 - 0x63
    "10110110", -- 6619 - 0x19db  :  182 - 0xb6
    "11011001", -- 6620 - 0x19dc  :  217 - 0xd9
    "11101011", -- 6621 - 0x19dd  :  235 - 0xeb
    "11110111", -- 6622 - 0x19de  :  247 - 0xf7
    "11111111", -- 6623 - 0x19df  :  255 - 0xff
    "00011100", -- 6624 - 0x19e0  :   28 - 0x1c -- Background 0x9e
    "00111100", -- 6625 - 0x19e1  :   60 - 0x3c
    "01111100", -- 6626 - 0x19e2  :  124 - 0x7c
    "11111100", -- 6627 - 0x19e3  :  252 - 0xfc
    "11111100", -- 6628 - 0x19e4  :  252 - 0xfc
    "11111100", -- 6629 - 0x19e5  :  252 - 0xfc
    "11111100", -- 6630 - 0x19e6  :  252 - 0xfc
    "11111100", -- 6631 - 0x19e7  :  252 - 0xfc
    "11011101", -- 6632 - 0x19e8  :  221 - 0xdd
    "10111101", -- 6633 - 0x19e9  :  189 - 0xbd
    "01111101", -- 6634 - 0x19ea  :  125 - 0x7d
    "11111101", -- 6635 - 0x19eb  :  253 - 0xfd
    "11111101", -- 6636 - 0x19ec  :  253 - 0xfd
    "11111101", -- 6637 - 0x19ed  :  253 - 0xfd
    "11111101", -- 6638 - 0x19ee  :  253 - 0xfd
    "11111101", -- 6639 - 0x19ef  :  253 - 0xfd
    "01111100", -- 6640 - 0x19f0  :  124 - 0x7c -- Background 0x9f
    "01111100", -- 6641 - 0x19f1  :  124 - 0x7c
    "01111000", -- 6642 - 0x19f2  :  120 - 0x78
    "01111000", -- 6643 - 0x19f3  :  120 - 0x78
    "01110001", -- 6644 - 0x19f4  :  113 - 0x71
    "01110001", -- 6645 - 0x19f5  :  113 - 0x71
    "01100011", -- 6646 - 0x19f6  :   99 - 0x63
    "01100011", -- 6647 - 0x19f7  :   99 - 0x63
    "00000001", -- 6648 - 0x19f8  :    1 - 0x1
    "00000001", -- 6649 - 0x19f9  :    1 - 0x1
    "00000010", -- 6650 - 0x19fa  :    2 - 0x2
    "00000010", -- 6651 - 0x19fb  :    2 - 0x2
    "00000101", -- 6652 - 0x19fc  :    5 - 0x5
    "00000101", -- 6653 - 0x19fd  :    5 - 0x5
    "00001011", -- 6654 - 0x19fe  :   11 - 0xb
    "00001011", -- 6655 - 0x19ff  :   11 - 0xb
    "01110001", -- 6656 - 0x1a00  :  113 - 0x71 -- Background 0xa0
    "01110000", -- 6657 - 0x1a01  :  112 - 0x70
    "11111000", -- 6658 - 0x1a02  :  248 - 0xf8
    "11111000", -- 6659 - 0x1a03  :  248 - 0xf8
    "11111100", -- 6660 - 0x1a04  :  252 - 0xfc
    "11111100", -- 6661 - 0x1a05  :  252 - 0xfc
    "11111110", -- 6662 - 0x1a06  :  254 - 0xfe
    "11111110", -- 6663 - 0x1a07  :  254 - 0xfe
    "01110100", -- 6664 - 0x1a08  :  116 - 0x74
    "01110110", -- 6665 - 0x1a09  :  118 - 0x76
    "11111010", -- 6666 - 0x1a0a  :  250 - 0xfa
    "11111011", -- 6667 - 0x1a0b  :  251 - 0xfb
    "11111101", -- 6668 - 0x1a0c  :  253 - 0xfd
    "11111101", -- 6669 - 0x1a0d  :  253 - 0xfd
    "11111110", -- 6670 - 0x1a0e  :  254 - 0xfe
    "11111110", -- 6671 - 0x1a0f  :  254 - 0xfe
    "11111000", -- 6672 - 0x1a10  :  248 - 0xf8 -- Background 0xa1
    "11111000", -- 6673 - 0x1a11  :  248 - 0xf8
    "11111000", -- 6674 - 0x1a12  :  248 - 0xf8
    "01111000", -- 6675 - 0x1a13  :  120 - 0x78
    "01111000", -- 6676 - 0x1a14  :  120 - 0x78
    "00111000", -- 6677 - 0x1a15  :   56 - 0x38
    "00111000", -- 6678 - 0x1a16  :   56 - 0x38
    "00011000", -- 6679 - 0x1a17  :   24 - 0x18
    "00000010", -- 6680 - 0x1a18  :    2 - 0x2
    "00000010", -- 6681 - 0x1a19  :    2 - 0x2
    "00000010", -- 6682 - 0x1a1a  :    2 - 0x2
    "00000010", -- 6683 - 0x1a1b  :    2 - 0x2
    "00000010", -- 6684 - 0x1a1c  :    2 - 0x2
    "10000010", -- 6685 - 0x1a1d  :  130 - 0x82
    "10000010", -- 6686 - 0x1a1e  :  130 - 0x82
    "11000010", -- 6687 - 0x1a1f  :  194 - 0xc2
    "11100000", -- 6688 - 0x1a20  :  224 - 0xe0 -- Background 0xa2
    "11110000", -- 6689 - 0x1a21  :  240 - 0xf0
    "11111000", -- 6690 - 0x1a22  :  248 - 0xf8
    "11111000", -- 6691 - 0x1a23  :  248 - 0xf8
    "11111100", -- 6692 - 0x1a24  :  252 - 0xfc
    "11111100", -- 6693 - 0x1a25  :  252 - 0xfc
    "11111110", -- 6694 - 0x1a26  :  254 - 0xfe
    "11111111", -- 6695 - 0x1a27  :  255 - 0xff
    "11101010", -- 6696 - 0x1a28  :  234 - 0xea
    "11110110", -- 6697 - 0x1a29  :  246 - 0xf6
    "11111010", -- 6698 - 0x1a2a  :  250 - 0xfa
    "11111010", -- 6699 - 0x1a2b  :  250 - 0xfa
    "11111100", -- 6700 - 0x1a2c  :  252 - 0xfc
    "11111100", -- 6701 - 0x1a2d  :  252 - 0xfc
    "11111110", -- 6702 - 0x1a2e  :  254 - 0xfe
    "11111111", -- 6703 - 0x1a2f  :  255 - 0xff
    "11111111", -- 6704 - 0x1a30  :  255 - 0xff -- Background 0xa3
    "11111111", -- 6705 - 0x1a31  :  255 - 0xff
    "11111111", -- 6706 - 0x1a32  :  255 - 0xff
    "11111111", -- 6707 - 0x1a33  :  255 - 0xff
    "11111111", -- 6708 - 0x1a34  :  255 - 0xff
    "11111111", -- 6709 - 0x1a35  :  255 - 0xff
    "11111111", -- 6710 - 0x1a36  :  255 - 0xff
    "11111111", -- 6711 - 0x1a37  :  255 - 0xff
    "11111111", -- 6712 - 0x1a38  :  255 - 0xff
    "11111111", -- 6713 - 0x1a39  :  255 - 0xff
    "11111111", -- 6714 - 0x1a3a  :  255 - 0xff
    "11111111", -- 6715 - 0x1a3b  :  255 - 0xff
    "11111111", -- 6716 - 0x1a3c  :  255 - 0xff
    "11111111", -- 6717 - 0x1a3d  :  255 - 0xff
    "11111111", -- 6718 - 0x1a3e  :  255 - 0xff
    "11111111", -- 6719 - 0x1a3f  :  255 - 0xff
    "00011111", -- 6720 - 0x1a40  :   31 - 0x1f -- Background 0xa4
    "00011111", -- 6721 - 0x1a41  :   31 - 0x1f
    "00011111", -- 6722 - 0x1a42  :   31 - 0x1f
    "00011111", -- 6723 - 0x1a43  :   31 - 0x1f
    "00011111", -- 6724 - 0x1a44  :   31 - 0x1f
    "00011111", -- 6725 - 0x1a45  :   31 - 0x1f
    "00011111", -- 6726 - 0x1a46  :   31 - 0x1f
    "00011111", -- 6727 - 0x1a47  :   31 - 0x1f
    "01000000", -- 6728 - 0x1a48  :   64 - 0x40
    "01000000", -- 6729 - 0x1a49  :   64 - 0x40
    "01000000", -- 6730 - 0x1a4a  :   64 - 0x40
    "01000000", -- 6731 - 0x1a4b  :   64 - 0x40
    "01000000", -- 6732 - 0x1a4c  :   64 - 0x40
    "01000000", -- 6733 - 0x1a4d  :   64 - 0x40
    "01000000", -- 6734 - 0x1a4e  :   64 - 0x40
    "01000000", -- 6735 - 0x1a4f  :   64 - 0x40
    "11111000", -- 6736 - 0x1a50  :  248 - 0xf8 -- Background 0xa5
    "11111111", -- 6737 - 0x1a51  :  255 - 0xff
    "11111111", -- 6738 - 0x1a52  :  255 - 0xff
    "11111000", -- 6739 - 0x1a53  :  248 - 0xf8
    "11111000", -- 6740 - 0x1a54  :  248 - 0xf8
    "11111000", -- 6741 - 0x1a55  :  248 - 0xf8
    "11111000", -- 6742 - 0x1a56  :  248 - 0xf8
    "11111000", -- 6743 - 0x1a57  :  248 - 0xf8
    "11111000", -- 6744 - 0x1a58  :  248 - 0xf8
    "11111111", -- 6745 - 0x1a59  :  255 - 0xff
    "11111111", -- 6746 - 0x1a5a  :  255 - 0xff
    "11111000", -- 6747 - 0x1a5b  :  248 - 0xf8
    "11111011", -- 6748 - 0x1a5c  :  251 - 0xfb
    "11111010", -- 6749 - 0x1a5d  :  250 - 0xfa
    "11111010", -- 6750 - 0x1a5e  :  250 - 0xfa
    "11111010", -- 6751 - 0x1a5f  :  250 - 0xfa
    "11111100", -- 6752 - 0x1a60  :  252 - 0xfc -- Background 0xa6
    "11111000", -- 6753 - 0x1a61  :  248 - 0xf8
    "11110000", -- 6754 - 0x1a62  :  240 - 0xf0
    "00000001", -- 6755 - 0x1a63  :    1 - 0x1
    "00000001", -- 6756 - 0x1a64  :    1 - 0x1
    "00000011", -- 6757 - 0x1a65  :    3 - 0x3
    "11000011", -- 6758 - 0x1a66  :  195 - 0xc3
    "10000111", -- 6759 - 0x1a67  :  135 - 0x87
    "11111100", -- 6760 - 0x1a68  :  252 - 0xfc
    "11111010", -- 6761 - 0x1a69  :  250 - 0xfa
    "11110110", -- 6762 - 0x1a6a  :  246 - 0xf6
    "00001101", -- 6763 - 0x1a6b  :   13 - 0xd
    "11111001", -- 6764 - 0x1a6c  :  249 - 0xf9
    "00000011", -- 6765 - 0x1a6d  :    3 - 0x3
    "00010011", -- 6766 - 0x1a6e  :   19 - 0x13
    "00110111", -- 6767 - 0x1a6f  :   55 - 0x37
    "01111111", -- 6768 - 0x1a70  :  127 - 0x7f -- Background 0xa7
    "11111001", -- 6769 - 0x1a71  :  249 - 0xf9
    "11111001", -- 6770 - 0x1a72  :  249 - 0xf9
    "11111111", -- 6771 - 0x1a73  :  255 - 0xff
    "11111110", -- 6772 - 0x1a74  :  254 - 0xfe
    "11111100", -- 6773 - 0x1a75  :  252 - 0xfc
    "11111111", -- 6774 - 0x1a76  :  255 - 0xff
    "11111111", -- 6775 - 0x1a77  :  255 - 0xff
    "01111111", -- 6776 - 0x1a78  :  127 - 0x7f
    "11111001", -- 6777 - 0x1a79  :  249 - 0xf9
    "11111001", -- 6778 - 0x1a7a  :  249 - 0xf9
    "11111111", -- 6779 - 0x1a7b  :  255 - 0xff
    "11111110", -- 6780 - 0x1a7c  :  254 - 0xfe
    "11111100", -- 6781 - 0x1a7d  :  252 - 0xfc
    "11111111", -- 6782 - 0x1a7e  :  255 - 0xff
    "11111111", -- 6783 - 0x1a7f  :  255 - 0xff
    "11110000", -- 6784 - 0x1a80  :  240 - 0xf0 -- Background 0xa8
    "11110000", -- 6785 - 0x1a81  :  240 - 0xf0
    "11111000", -- 6786 - 0x1a82  :  248 - 0xf8
    "01111000", -- 6787 - 0x1a83  :  120 - 0x78
    "11111100", -- 6788 - 0x1a84  :  252 - 0xfc
    "11110100", -- 6789 - 0x1a85  :  244 - 0xf4
    "11110110", -- 6790 - 0x1a86  :  246 - 0xf6
    "11111010", -- 6791 - 0x1a87  :  250 - 0xfa
    "11110110", -- 6792 - 0x1a88  :  246 - 0xf6
    "11110110", -- 6793 - 0x1a89  :  246 - 0xf6
    "11111011", -- 6794 - 0x1a8a  :  251 - 0xfb
    "01111011", -- 6795 - 0x1a8b  :  123 - 0x7b
    "11111101", -- 6796 - 0x1a8c  :  253 - 0xfd
    "11110101", -- 6797 - 0x1a8d  :  245 - 0xf5
    "11110110", -- 6798 - 0x1a8e  :  246 - 0xf6
    "11111010", -- 6799 - 0x1a8f  :  250 - 0xfa
    "00111111", -- 6800 - 0x1a90  :   63 - 0x3f -- Background 0xa9
    "00111111", -- 6801 - 0x1a91  :   63 - 0x3f
    "00111111", -- 6802 - 0x1a92  :   63 - 0x3f
    "00111111", -- 6803 - 0x1a93  :   63 - 0x3f
    "00111111", -- 6804 - 0x1a94  :   63 - 0x3f
    "00011111", -- 6805 - 0x1a95  :   31 - 0x1f
    "00001111", -- 6806 - 0x1a96  :   15 - 0xf
    "00000111", -- 6807 - 0x1a97  :    7 - 0x7
    "10111111", -- 6808 - 0x1a98  :  191 - 0xbf
    "10111111", -- 6809 - 0x1a99  :  191 - 0xbf
    "00111111", -- 6810 - 0x1a9a  :   63 - 0x3f
    "00111111", -- 6811 - 0x1a9b  :   63 - 0x3f
    "10111111", -- 6812 - 0x1a9c  :  191 - 0xbf
    "10011111", -- 6813 - 0x1a9d  :  159 - 0x9f
    "11001111", -- 6814 - 0x1a9e  :  207 - 0xcf
    "11010111", -- 6815 - 0x1a9f  :  215 - 0xd7
    "11100000", -- 6816 - 0x1aa0  :  224 - 0xe0 -- Background 0xaa
    "11111000", -- 6817 - 0x1aa1  :  248 - 0xf8
    "11111111", -- 6818 - 0x1aa2  :  255 - 0xff
    "11110011", -- 6819 - 0x1aa3  :  243 - 0xf3
    "11111100", -- 6820 - 0x1aa4  :  252 - 0xfc
    "11111111", -- 6821 - 0x1aa5  :  255 - 0xff
    "11111111", -- 6822 - 0x1aa6  :  255 - 0xff
    "11111111", -- 6823 - 0x1aa7  :  255 - 0xff
    "11100100", -- 6824 - 0x1aa8  :  228 - 0xe4
    "11111000", -- 6825 - 0x1aa9  :  248 - 0xf8
    "11111111", -- 6826 - 0x1aaa  :  255 - 0xff
    "11110011", -- 6827 - 0x1aab  :  243 - 0xf3
    "11111100", -- 6828 - 0x1aac  :  252 - 0xfc
    "11111111", -- 6829 - 0x1aad  :  255 - 0xff
    "11111111", -- 6830 - 0x1aae  :  255 - 0xff
    "11111111", -- 6831 - 0x1aaf  :  255 - 0xff
    "11111111", -- 6832 - 0x1ab0  :  255 - 0xff -- Background 0xab
    "11111111", -- 6833 - 0x1ab1  :  255 - 0xff
    "00111111", -- 6834 - 0x1ab2  :   63 - 0x3f
    "11001111", -- 6835 - 0x1ab3  :  207 - 0xcf
    "11110011", -- 6836 - 0x1ab4  :  243 - 0xf3
    "00111101", -- 6837 - 0x1ab5  :   61 - 0x3d
    "11011000", -- 6838 - 0x1ab6  :  216 - 0xd8
    "10110000", -- 6839 - 0x1ab7  :  176 - 0xb0
    "00000000", -- 6840 - 0x1ab8  :    0 - 0x0
    "00000000", -- 6841 - 0x1ab9  :    0 - 0x0
    "00000000", -- 6842 - 0x1aba  :    0 - 0x0
    "11000000", -- 6843 - 0x1abb  :  192 - 0xc0
    "11110000", -- 6844 - 0x1abc  :  240 - 0xf0
    "00111100", -- 6845 - 0x1abd  :   60 - 0x3c
    "11011000", -- 6846 - 0x1abe  :  216 - 0xd8
    "10110110", -- 6847 - 0x1abf  :  182 - 0xb6
    "10001111", -- 6848 - 0x1ac0  :  143 - 0x8f -- Background 0xac
    "11101111", -- 6849 - 0x1ac1  :  239 - 0xef
    "11100000", -- 6850 - 0x1ac2  :  224 - 0xe0
    "11111000", -- 6851 - 0x1ac3  :  248 - 0xf8
    "11111000", -- 6852 - 0x1ac4  :  248 - 0xf8
    "11111111", -- 6853 - 0x1ac5  :  255 - 0xff
    "11111111", -- 6854 - 0x1ac6  :  255 - 0xff
    "11111111", -- 6855 - 0x1ac7  :  255 - 0xff
    "00001111", -- 6856 - 0x1ac8  :   15 - 0xf
    "00001111", -- 6857 - 0x1ac9  :   15 - 0xf
    "00000000", -- 6858 - 0x1aca  :    0 - 0x0
    "00000011", -- 6859 - 0x1acb  :    3 - 0x3
    "00000000", -- 6860 - 0x1acc  :    0 - 0x0
    "00000000", -- 6861 - 0x1acd  :    0 - 0x0
    "00000000", -- 6862 - 0x1ace  :    0 - 0x0
    "00000000", -- 6863 - 0x1acf  :    0 - 0x0
    "11110001", -- 6864 - 0x1ad0  :  241 - 0xf1 -- Background 0xad
    "11110001", -- 6865 - 0x1ad1  :  241 - 0xf1
    "00000001", -- 6866 - 0x1ad2  :    1 - 0x1
    "00000001", -- 6867 - 0x1ad3  :    1 - 0x1
    "00000001", -- 6868 - 0x1ad4  :    1 - 0x1
    "11111111", -- 6869 - 0x1ad5  :  255 - 0xff
    "11111111", -- 6870 - 0x1ad6  :  255 - 0xff
    "11111111", -- 6871 - 0x1ad7  :  255 - 0xff
    "11110100", -- 6872 - 0x1ad8  :  244 - 0xf4
    "11110100", -- 6873 - 0x1ad9  :  244 - 0xf4
    "00000100", -- 6874 - 0x1ada  :    4 - 0x4
    "11111100", -- 6875 - 0x1adb  :  252 - 0xfc
    "00000000", -- 6876 - 0x1adc  :    0 - 0x0
    "00000000", -- 6877 - 0x1add  :    0 - 0x0
    "00000000", -- 6878 - 0x1ade  :    0 - 0x0
    "00000000", -- 6879 - 0x1adf  :    0 - 0x0
    "00011111", -- 6880 - 0x1ae0  :   31 - 0x1f -- Background 0xae
    "00011111", -- 6881 - 0x1ae1  :   31 - 0x1f
    "00011111", -- 6882 - 0x1ae2  :   31 - 0x1f
    "00011111", -- 6883 - 0x1ae3  :   31 - 0x1f
    "00011111", -- 6884 - 0x1ae4  :   31 - 0x1f
    "00011111", -- 6885 - 0x1ae5  :   31 - 0x1f
    "00011111", -- 6886 - 0x1ae6  :   31 - 0x1f
    "00011111", -- 6887 - 0x1ae7  :   31 - 0x1f
    "01011111", -- 6888 - 0x1ae8  :   95 - 0x5f
    "01011111", -- 6889 - 0x1ae9  :   95 - 0x5f
    "01011111", -- 6890 - 0x1aea  :   95 - 0x5f
    "01011111", -- 6891 - 0x1aeb  :   95 - 0x5f
    "01011111", -- 6892 - 0x1aec  :   95 - 0x5f
    "01011111", -- 6893 - 0x1aed  :   95 - 0x5f
    "01011111", -- 6894 - 0x1aee  :   95 - 0x5f
    "01011111", -- 6895 - 0x1aef  :   95 - 0x5f
    "11111100", -- 6896 - 0x1af0  :  252 - 0xfc -- Background 0xaf
    "11111100", -- 6897 - 0x1af1  :  252 - 0xfc
    "11111100", -- 6898 - 0x1af2  :  252 - 0xfc
    "11111100", -- 6899 - 0x1af3  :  252 - 0xfc
    "11110100", -- 6900 - 0x1af4  :  244 - 0xf4
    "11110100", -- 6901 - 0x1af5  :  244 - 0xf4
    "11110100", -- 6902 - 0x1af6  :  244 - 0xf4
    "11110100", -- 6903 - 0x1af7  :  244 - 0xf4
    "11111101", -- 6904 - 0x1af8  :  253 - 0xfd
    "11111101", -- 6905 - 0x1af9  :  253 - 0xfd
    "11111101", -- 6906 - 0x1afa  :  253 - 0xfd
    "11111101", -- 6907 - 0x1afb  :  253 - 0xfd
    "11110101", -- 6908 - 0x1afc  :  245 - 0xf5
    "11110101", -- 6909 - 0x1afd  :  245 - 0xf5
    "11110101", -- 6910 - 0x1afe  :  245 - 0xf5
    "11110101", -- 6911 - 0x1aff  :  245 - 0xf5
    "00001100", -- 6912 - 0x1b00  :   12 - 0xc -- Background 0xb0
    "00011100", -- 6913 - 0x1b01  :   28 - 0x1c
    "00001100", -- 6914 - 0x1b02  :   12 - 0xc
    "00001100", -- 6915 - 0x1b03  :   12 - 0xc
    "00001100", -- 6916 - 0x1b04  :   12 - 0xc
    "00001100", -- 6917 - 0x1b05  :   12 - 0xc
    "00111111", -- 6918 - 0x1b06  :   63 - 0x3f
    "00000000", -- 6919 - 0x1b07  :    0 - 0x0
    "00001100", -- 6920 - 0x1b08  :   12 - 0xc
    "00011100", -- 6921 - 0x1b09  :   28 - 0x1c
    "00001100", -- 6922 - 0x1b0a  :   12 - 0xc
    "00001100", -- 6923 - 0x1b0b  :   12 - 0xc
    "00001100", -- 6924 - 0x1b0c  :   12 - 0xc
    "00001100", -- 6925 - 0x1b0d  :   12 - 0xc
    "00111111", -- 6926 - 0x1b0e  :   63 - 0x3f
    "00000000", -- 6927 - 0x1b0f  :    0 - 0x0
    "00111110", -- 6928 - 0x1b10  :   62 - 0x3e -- Background 0xb1
    "01100011", -- 6929 - 0x1b11  :   99 - 0x63
    "00000111", -- 6930 - 0x1b12  :    7 - 0x7
    "00011110", -- 6931 - 0x1b13  :   30 - 0x1e
    "00111100", -- 6932 - 0x1b14  :   60 - 0x3c
    "01110000", -- 6933 - 0x1b15  :  112 - 0x70
    "01111111", -- 6934 - 0x1b16  :  127 - 0x7f
    "00000000", -- 6935 - 0x1b17  :    0 - 0x0
    "00111110", -- 6936 - 0x1b18  :   62 - 0x3e
    "01100011", -- 6937 - 0x1b19  :   99 - 0x63
    "00000111", -- 6938 - 0x1b1a  :    7 - 0x7
    "00011110", -- 6939 - 0x1b1b  :   30 - 0x1e
    "00111100", -- 6940 - 0x1b1c  :   60 - 0x3c
    "01110000", -- 6941 - 0x1b1d  :  112 - 0x70
    "01111111", -- 6942 - 0x1b1e  :  127 - 0x7f
    "00000000", -- 6943 - 0x1b1f  :    0 - 0x0
    "01111110", -- 6944 - 0x1b20  :  126 - 0x7e -- Background 0xb2
    "01100011", -- 6945 - 0x1b21  :   99 - 0x63
    "01100011", -- 6946 - 0x1b22  :   99 - 0x63
    "01100011", -- 6947 - 0x1b23  :   99 - 0x63
    "01111110", -- 6948 - 0x1b24  :  126 - 0x7e
    "01100000", -- 6949 - 0x1b25  :   96 - 0x60
    "01100000", -- 6950 - 0x1b26  :   96 - 0x60
    "00000000", -- 6951 - 0x1b27  :    0 - 0x0
    "01111110", -- 6952 - 0x1b28  :  126 - 0x7e
    "01100011", -- 6953 - 0x1b29  :   99 - 0x63
    "01100011", -- 6954 - 0x1b2a  :   99 - 0x63
    "01100011", -- 6955 - 0x1b2b  :   99 - 0x63
    "01111110", -- 6956 - 0x1b2c  :  126 - 0x7e
    "01100000", -- 6957 - 0x1b2d  :   96 - 0x60
    "01100000", -- 6958 - 0x1b2e  :   96 - 0x60
    "00000000", -- 6959 - 0x1b2f  :    0 - 0x0
    "01100011", -- 6960 - 0x1b30  :   99 - 0x63 -- Background 0xb3
    "01100011", -- 6961 - 0x1b31  :   99 - 0x63
    "01100011", -- 6962 - 0x1b32  :   99 - 0x63
    "01100011", -- 6963 - 0x1b33  :   99 - 0x63
    "01100011", -- 6964 - 0x1b34  :   99 - 0x63
    "01100011", -- 6965 - 0x1b35  :   99 - 0x63
    "00111110", -- 6966 - 0x1b36  :   62 - 0x3e
    "00000000", -- 6967 - 0x1b37  :    0 - 0x0
    "01100011", -- 6968 - 0x1b38  :   99 - 0x63
    "01100011", -- 6969 - 0x1b39  :   99 - 0x63
    "01100011", -- 6970 - 0x1b3a  :   99 - 0x63
    "01100011", -- 6971 - 0x1b3b  :   99 - 0x63
    "01100011", -- 6972 - 0x1b3c  :   99 - 0x63
    "01100011", -- 6973 - 0x1b3d  :   99 - 0x63
    "00111110", -- 6974 - 0x1b3e  :   62 - 0x3e
    "00000000", -- 6975 - 0x1b3f  :    0 - 0x0
    "01100011", -- 6976 - 0x1b40  :   99 - 0x63 -- Background 0xb4
    "01100011", -- 6977 - 0x1b41  :   99 - 0x63
    "01100011", -- 6978 - 0x1b42  :   99 - 0x63
    "01111111", -- 6979 - 0x1b43  :  127 - 0x7f
    "01100011", -- 6980 - 0x1b44  :   99 - 0x63
    "01100011", -- 6981 - 0x1b45  :   99 - 0x63
    "01100011", -- 6982 - 0x1b46  :   99 - 0x63
    "00000000", -- 6983 - 0x1b47  :    0 - 0x0
    "01100011", -- 6984 - 0x1b48  :   99 - 0x63
    "01100011", -- 6985 - 0x1b49  :   99 - 0x63
    "01100011", -- 6986 - 0x1b4a  :   99 - 0x63
    "01111111", -- 6987 - 0x1b4b  :  127 - 0x7f
    "01100011", -- 6988 - 0x1b4c  :   99 - 0x63
    "01100011", -- 6989 - 0x1b4d  :   99 - 0x63
    "01100011", -- 6990 - 0x1b4e  :   99 - 0x63
    "00000000", -- 6991 - 0x1b4f  :    0 - 0x0
    "00111111", -- 6992 - 0x1b50  :   63 - 0x3f -- Background 0xb5
    "00001100", -- 6993 - 0x1b51  :   12 - 0xc
    "00001100", -- 6994 - 0x1b52  :   12 - 0xc
    "00001100", -- 6995 - 0x1b53  :   12 - 0xc
    "00001100", -- 6996 - 0x1b54  :   12 - 0xc
    "00001100", -- 6997 - 0x1b55  :   12 - 0xc
    "00111111", -- 6998 - 0x1b56  :   63 - 0x3f
    "00000000", -- 6999 - 0x1b57  :    0 - 0x0
    "00111111", -- 7000 - 0x1b58  :   63 - 0x3f
    "00001100", -- 7001 - 0x1b59  :   12 - 0xc
    "00001100", -- 7002 - 0x1b5a  :   12 - 0xc
    "00001100", -- 7003 - 0x1b5b  :   12 - 0xc
    "00001100", -- 7004 - 0x1b5c  :   12 - 0xc
    "00001100", -- 7005 - 0x1b5d  :   12 - 0xc
    "00111111", -- 7006 - 0x1b5e  :   63 - 0x3f
    "00000000", -- 7007 - 0x1b5f  :    0 - 0x0
    "00000000", -- 7008 - 0x1b60  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 7009 - 0x1b61  :    0 - 0x0
    "00000000", -- 7010 - 0x1b62  :    0 - 0x0
    "01111110", -- 7011 - 0x1b63  :  126 - 0x7e
    "00000000", -- 7012 - 0x1b64  :    0 - 0x0
    "00000000", -- 7013 - 0x1b65  :    0 - 0x0
    "00000000", -- 7014 - 0x1b66  :    0 - 0x0
    "00000000", -- 7015 - 0x1b67  :    0 - 0x0
    "00000000", -- 7016 - 0x1b68  :    0 - 0x0
    "00000000", -- 7017 - 0x1b69  :    0 - 0x0
    "00000000", -- 7018 - 0x1b6a  :    0 - 0x0
    "01111110", -- 7019 - 0x1b6b  :  126 - 0x7e
    "00000000", -- 7020 - 0x1b6c  :    0 - 0x0
    "00000000", -- 7021 - 0x1b6d  :    0 - 0x0
    "00000000", -- 7022 - 0x1b6e  :    0 - 0x0
    "00000000", -- 7023 - 0x1b6f  :    0 - 0x0
    "00111100", -- 7024 - 0x1b70  :   60 - 0x3c -- Background 0xb7
    "01100110", -- 7025 - 0x1b71  :  102 - 0x66
    "01100000", -- 7026 - 0x1b72  :   96 - 0x60
    "00111110", -- 7027 - 0x1b73  :   62 - 0x3e
    "00000011", -- 7028 - 0x1b74  :    3 - 0x3
    "01100011", -- 7029 - 0x1b75  :   99 - 0x63
    "00111110", -- 7030 - 0x1b76  :   62 - 0x3e
    "00000000", -- 7031 - 0x1b77  :    0 - 0x0
    "00111100", -- 7032 - 0x1b78  :   60 - 0x3c
    "01100110", -- 7033 - 0x1b79  :  102 - 0x66
    "01100000", -- 7034 - 0x1b7a  :   96 - 0x60
    "00111110", -- 7035 - 0x1b7b  :   62 - 0x3e
    "00000011", -- 7036 - 0x1b7c  :    3 - 0x3
    "01100011", -- 7037 - 0x1b7d  :   99 - 0x63
    "00111110", -- 7038 - 0x1b7e  :   62 - 0x3e
    "00000000", -- 7039 - 0x1b7f  :    0 - 0x0
    "00011110", -- 7040 - 0x1b80  :   30 - 0x1e -- Background 0xb8
    "00110011", -- 7041 - 0x1b81  :   51 - 0x33
    "01100000", -- 7042 - 0x1b82  :   96 - 0x60
    "01100000", -- 7043 - 0x1b83  :   96 - 0x60
    "01100000", -- 7044 - 0x1b84  :   96 - 0x60
    "00110011", -- 7045 - 0x1b85  :   51 - 0x33
    "00011110", -- 7046 - 0x1b86  :   30 - 0x1e
    "00000000", -- 7047 - 0x1b87  :    0 - 0x0
    "00011110", -- 7048 - 0x1b88  :   30 - 0x1e
    "00110011", -- 7049 - 0x1b89  :   51 - 0x33
    "01100000", -- 7050 - 0x1b8a  :   96 - 0x60
    "01100000", -- 7051 - 0x1b8b  :   96 - 0x60
    "01100000", -- 7052 - 0x1b8c  :   96 - 0x60
    "00110011", -- 7053 - 0x1b8d  :   51 - 0x33
    "00011110", -- 7054 - 0x1b8e  :   30 - 0x1e
    "00000000", -- 7055 - 0x1b8f  :    0 - 0x0
    "00111110", -- 7056 - 0x1b90  :   62 - 0x3e -- Background 0xb9
    "01100011", -- 7057 - 0x1b91  :   99 - 0x63
    "01100011", -- 7058 - 0x1b92  :   99 - 0x63
    "01100011", -- 7059 - 0x1b93  :   99 - 0x63
    "01100011", -- 7060 - 0x1b94  :   99 - 0x63
    "01100011", -- 7061 - 0x1b95  :   99 - 0x63
    "00111110", -- 7062 - 0x1b96  :   62 - 0x3e
    "00000000", -- 7063 - 0x1b97  :    0 - 0x0
    "00111110", -- 7064 - 0x1b98  :   62 - 0x3e
    "01100011", -- 7065 - 0x1b99  :   99 - 0x63
    "01100011", -- 7066 - 0x1b9a  :   99 - 0x63
    "01100011", -- 7067 - 0x1b9b  :   99 - 0x63
    "01100011", -- 7068 - 0x1b9c  :   99 - 0x63
    "01100011", -- 7069 - 0x1b9d  :   99 - 0x63
    "00111110", -- 7070 - 0x1b9e  :   62 - 0x3e
    "00000000", -- 7071 - 0x1b9f  :    0 - 0x0
    "01111110", -- 7072 - 0x1ba0  :  126 - 0x7e -- Background 0xba
    "01100011", -- 7073 - 0x1ba1  :   99 - 0x63
    "01100011", -- 7074 - 0x1ba2  :   99 - 0x63
    "01100111", -- 7075 - 0x1ba3  :  103 - 0x67
    "01111100", -- 7076 - 0x1ba4  :  124 - 0x7c
    "01101110", -- 7077 - 0x1ba5  :  110 - 0x6e
    "01100111", -- 7078 - 0x1ba6  :  103 - 0x67
    "00000000", -- 7079 - 0x1ba7  :    0 - 0x0
    "01111110", -- 7080 - 0x1ba8  :  126 - 0x7e
    "01100011", -- 7081 - 0x1ba9  :   99 - 0x63
    "01100011", -- 7082 - 0x1baa  :   99 - 0x63
    "01100111", -- 7083 - 0x1bab  :  103 - 0x67
    "01111100", -- 7084 - 0x1bac  :  124 - 0x7c
    "01101110", -- 7085 - 0x1bad  :  110 - 0x6e
    "01100111", -- 7086 - 0x1bae  :  103 - 0x67
    "00000000", -- 7087 - 0x1baf  :    0 - 0x0
    "01111111", -- 7088 - 0x1bb0  :  127 - 0x7f -- Background 0xbb
    "01100000", -- 7089 - 0x1bb1  :   96 - 0x60
    "01100000", -- 7090 - 0x1bb2  :   96 - 0x60
    "01111110", -- 7091 - 0x1bb3  :  126 - 0x7e
    "01100000", -- 7092 - 0x1bb4  :   96 - 0x60
    "01100000", -- 7093 - 0x1bb5  :   96 - 0x60
    "01111111", -- 7094 - 0x1bb6  :  127 - 0x7f
    "00000000", -- 7095 - 0x1bb7  :    0 - 0x0
    "01111111", -- 7096 - 0x1bb8  :  127 - 0x7f
    "01100000", -- 7097 - 0x1bb9  :   96 - 0x60
    "01100000", -- 7098 - 0x1bba  :   96 - 0x60
    "01111110", -- 7099 - 0x1bbb  :  126 - 0x7e
    "01100000", -- 7100 - 0x1bbc  :   96 - 0x60
    "01100000", -- 7101 - 0x1bbd  :   96 - 0x60
    "01111111", -- 7102 - 0x1bbe  :  127 - 0x7f
    "00000000", -- 7103 - 0x1bbf  :    0 - 0x0
    "00000000", -- 7104 - 0x1bc0  :    0 - 0x0 -- Background 0xbc
    "00100010", -- 7105 - 0x1bc1  :   34 - 0x22
    "01100101", -- 7106 - 0x1bc2  :  101 - 0x65
    "00100101", -- 7107 - 0x1bc3  :   37 - 0x25
    "00100101", -- 7108 - 0x1bc4  :   37 - 0x25
    "01110010", -- 7109 - 0x1bc5  :  114 - 0x72
    "00000000", -- 7110 - 0x1bc6  :    0 - 0x0
    "00000000", -- 7111 - 0x1bc7  :    0 - 0x0
    "00000000", -- 7112 - 0x1bc8  :    0 - 0x0
    "00000000", -- 7113 - 0x1bc9  :    0 - 0x0
    "00000000", -- 7114 - 0x1bca  :    0 - 0x0
    "00000000", -- 7115 - 0x1bcb  :    0 - 0x0
    "00000000", -- 7116 - 0x1bcc  :    0 - 0x0
    "00000000", -- 7117 - 0x1bcd  :    0 - 0x0
    "00000000", -- 7118 - 0x1bce  :    0 - 0x0
    "00000000", -- 7119 - 0x1bcf  :    0 - 0x0
    "00000000", -- 7120 - 0x1bd0  :    0 - 0x0 -- Background 0xbd
    "01110010", -- 7121 - 0x1bd1  :  114 - 0x72
    "01000101", -- 7122 - 0x1bd2  :   69 - 0x45
    "01100101", -- 7123 - 0x1bd3  :  101 - 0x65
    "00010101", -- 7124 - 0x1bd4  :   21 - 0x15
    "01100010", -- 7125 - 0x1bd5  :   98 - 0x62
    "00000000", -- 7126 - 0x1bd6  :    0 - 0x0
    "00000000", -- 7127 - 0x1bd7  :    0 - 0x0
    "00000000", -- 7128 - 0x1bd8  :    0 - 0x0
    "00000000", -- 7129 - 0x1bd9  :    0 - 0x0
    "00000000", -- 7130 - 0x1bda  :    0 - 0x0
    "00000000", -- 7131 - 0x1bdb  :    0 - 0x0
    "00000000", -- 7132 - 0x1bdc  :    0 - 0x0
    "00000000", -- 7133 - 0x1bdd  :    0 - 0x0
    "00000000", -- 7134 - 0x1bde  :    0 - 0x0
    "00000000", -- 7135 - 0x1bdf  :    0 - 0x0
    "00000000", -- 7136 - 0x1be0  :    0 - 0x0 -- Background 0xbe
    "01100111", -- 7137 - 0x1be1  :  103 - 0x67
    "01010010", -- 7138 - 0x1be2  :   82 - 0x52
    "01100010", -- 7139 - 0x1be3  :   98 - 0x62
    "01000010", -- 7140 - 0x1be4  :   66 - 0x42
    "01000010", -- 7141 - 0x1be5  :   66 - 0x42
    "00000000", -- 7142 - 0x1be6  :    0 - 0x0
    "00000000", -- 7143 - 0x1be7  :    0 - 0x0
    "00000000", -- 7144 - 0x1be8  :    0 - 0x0
    "00000000", -- 7145 - 0x1be9  :    0 - 0x0
    "00000000", -- 7146 - 0x1bea  :    0 - 0x0
    "00000000", -- 7147 - 0x1beb  :    0 - 0x0
    "00000000", -- 7148 - 0x1bec  :    0 - 0x0
    "00000000", -- 7149 - 0x1bed  :    0 - 0x0
    "00000000", -- 7150 - 0x1bee  :    0 - 0x0
    "00000000", -- 7151 - 0x1bef  :    0 - 0x0
    "00000000", -- 7152 - 0x1bf0  :    0 - 0x0 -- Background 0xbf
    "01100000", -- 7153 - 0x1bf1  :   96 - 0x60
    "10000000", -- 7154 - 0x1bf2  :  128 - 0x80
    "01000000", -- 7155 - 0x1bf3  :   64 - 0x40
    "00100000", -- 7156 - 0x1bf4  :   32 - 0x20
    "11000110", -- 7157 - 0x1bf5  :  198 - 0xc6
    "00000000", -- 7158 - 0x1bf6  :    0 - 0x0
    "00000000", -- 7159 - 0x1bf7  :    0 - 0x0
    "00000000", -- 7160 - 0x1bf8  :    0 - 0x0
    "00000000", -- 7161 - 0x1bf9  :    0 - 0x0
    "00000000", -- 7162 - 0x1bfa  :    0 - 0x0
    "00000000", -- 7163 - 0x1bfb  :    0 - 0x0
    "00000000", -- 7164 - 0x1bfc  :    0 - 0x0
    "00000000", -- 7165 - 0x1bfd  :    0 - 0x0
    "00000000", -- 7166 - 0x1bfe  :    0 - 0x0
    "00000000", -- 7167 - 0x1bff  :    0 - 0x0
    "01100011", -- 7168 - 0x1c00  :   99 - 0x63 -- Background 0xc0
    "01100110", -- 7169 - 0x1c01  :  102 - 0x66
    "01101100", -- 7170 - 0x1c02  :  108 - 0x6c
    "01111000", -- 7171 - 0x1c03  :  120 - 0x78
    "01111100", -- 7172 - 0x1c04  :  124 - 0x7c
    "01100110", -- 7173 - 0x1c05  :  102 - 0x66
    "01100011", -- 7174 - 0x1c06  :   99 - 0x63
    "00000000", -- 7175 - 0x1c07  :    0 - 0x0
    "01100011", -- 7176 - 0x1c08  :   99 - 0x63
    "01100110", -- 7177 - 0x1c09  :  102 - 0x66
    "01101100", -- 7178 - 0x1c0a  :  108 - 0x6c
    "01111000", -- 7179 - 0x1c0b  :  120 - 0x78
    "01111100", -- 7180 - 0x1c0c  :  124 - 0x7c
    "01100110", -- 7181 - 0x1c0d  :  102 - 0x66
    "01100011", -- 7182 - 0x1c0e  :   99 - 0x63
    "00000000", -- 7183 - 0x1c0f  :    0 - 0x0
    "00111111", -- 7184 - 0x1c10  :   63 - 0x3f -- Background 0xc1
    "00001100", -- 7185 - 0x1c11  :   12 - 0xc
    "00001100", -- 7186 - 0x1c12  :   12 - 0xc
    "00001100", -- 7187 - 0x1c13  :   12 - 0xc
    "00001100", -- 7188 - 0x1c14  :   12 - 0xc
    "00001100", -- 7189 - 0x1c15  :   12 - 0xc
    "00111111", -- 7190 - 0x1c16  :   63 - 0x3f
    "00000000", -- 7191 - 0x1c17  :    0 - 0x0
    "00111111", -- 7192 - 0x1c18  :   63 - 0x3f
    "00001100", -- 7193 - 0x1c19  :   12 - 0xc
    "00001100", -- 7194 - 0x1c1a  :   12 - 0xc
    "00001100", -- 7195 - 0x1c1b  :   12 - 0xc
    "00001100", -- 7196 - 0x1c1c  :   12 - 0xc
    "00001100", -- 7197 - 0x1c1d  :   12 - 0xc
    "00111111", -- 7198 - 0x1c1e  :   63 - 0x3f
    "00000000", -- 7199 - 0x1c1f  :    0 - 0x0
    "01100011", -- 7200 - 0x1c20  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 7201 - 0x1c21  :  119 - 0x77
    "01111111", -- 7202 - 0x1c22  :  127 - 0x7f
    "01111111", -- 7203 - 0x1c23  :  127 - 0x7f
    "01101011", -- 7204 - 0x1c24  :  107 - 0x6b
    "01100011", -- 7205 - 0x1c25  :   99 - 0x63
    "01100011", -- 7206 - 0x1c26  :   99 - 0x63
    "00000000", -- 7207 - 0x1c27  :    0 - 0x0
    "01100011", -- 7208 - 0x1c28  :   99 - 0x63
    "01110111", -- 7209 - 0x1c29  :  119 - 0x77
    "01111111", -- 7210 - 0x1c2a  :  127 - 0x7f
    "01111111", -- 7211 - 0x1c2b  :  127 - 0x7f
    "01101011", -- 7212 - 0x1c2c  :  107 - 0x6b
    "01100011", -- 7213 - 0x1c2d  :   99 - 0x63
    "01100011", -- 7214 - 0x1c2e  :   99 - 0x63
    "00000000", -- 7215 - 0x1c2f  :    0 - 0x0
    "00011100", -- 7216 - 0x1c30  :   28 - 0x1c -- Background 0xc3
    "00110110", -- 7217 - 0x1c31  :   54 - 0x36
    "01100011", -- 7218 - 0x1c32  :   99 - 0x63
    "01100011", -- 7219 - 0x1c33  :   99 - 0x63
    "01111111", -- 7220 - 0x1c34  :  127 - 0x7f
    "01100011", -- 7221 - 0x1c35  :   99 - 0x63
    "01100011", -- 7222 - 0x1c36  :   99 - 0x63
    "00000000", -- 7223 - 0x1c37  :    0 - 0x0
    "00011100", -- 7224 - 0x1c38  :   28 - 0x1c
    "00110110", -- 7225 - 0x1c39  :   54 - 0x36
    "01100011", -- 7226 - 0x1c3a  :   99 - 0x63
    "01100011", -- 7227 - 0x1c3b  :   99 - 0x63
    "01111111", -- 7228 - 0x1c3c  :  127 - 0x7f
    "01100011", -- 7229 - 0x1c3d  :   99 - 0x63
    "01100011", -- 7230 - 0x1c3e  :   99 - 0x63
    "00000000", -- 7231 - 0x1c3f  :    0 - 0x0
    "00011111", -- 7232 - 0x1c40  :   31 - 0x1f -- Background 0xc4
    "00110000", -- 7233 - 0x1c41  :   48 - 0x30
    "01100000", -- 7234 - 0x1c42  :   96 - 0x60
    "01100111", -- 7235 - 0x1c43  :  103 - 0x67
    "01100011", -- 7236 - 0x1c44  :   99 - 0x63
    "00110011", -- 7237 - 0x1c45  :   51 - 0x33
    "00011111", -- 7238 - 0x1c46  :   31 - 0x1f
    "00000000", -- 7239 - 0x1c47  :    0 - 0x0
    "00011111", -- 7240 - 0x1c48  :   31 - 0x1f
    "00110000", -- 7241 - 0x1c49  :   48 - 0x30
    "01100000", -- 7242 - 0x1c4a  :   96 - 0x60
    "01100111", -- 7243 - 0x1c4b  :  103 - 0x67
    "01100011", -- 7244 - 0x1c4c  :   99 - 0x63
    "00110011", -- 7245 - 0x1c4d  :   51 - 0x33
    "00011111", -- 7246 - 0x1c4e  :   31 - 0x1f
    "00000000", -- 7247 - 0x1c4f  :    0 - 0x0
    "01100011", -- 7248 - 0x1c50  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 7249 - 0x1c51  :   99 - 0x63
    "01100011", -- 7250 - 0x1c52  :   99 - 0x63
    "01100011", -- 7251 - 0x1c53  :   99 - 0x63
    "01100011", -- 7252 - 0x1c54  :   99 - 0x63
    "01100011", -- 7253 - 0x1c55  :   99 - 0x63
    "00111110", -- 7254 - 0x1c56  :   62 - 0x3e
    "00000000", -- 7255 - 0x1c57  :    0 - 0x0
    "01100011", -- 7256 - 0x1c58  :   99 - 0x63
    "01100011", -- 7257 - 0x1c59  :   99 - 0x63
    "01100011", -- 7258 - 0x1c5a  :   99 - 0x63
    "01100011", -- 7259 - 0x1c5b  :   99 - 0x63
    "01100011", -- 7260 - 0x1c5c  :   99 - 0x63
    "01100011", -- 7261 - 0x1c5d  :   99 - 0x63
    "00111110", -- 7262 - 0x1c5e  :   62 - 0x3e
    "00000000", -- 7263 - 0x1c5f  :    0 - 0x0
    "01111110", -- 7264 - 0x1c60  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 7265 - 0x1c61  :   99 - 0x63
    "01100011", -- 7266 - 0x1c62  :   99 - 0x63
    "01100111", -- 7267 - 0x1c63  :  103 - 0x67
    "01111100", -- 7268 - 0x1c64  :  124 - 0x7c
    "01101110", -- 7269 - 0x1c65  :  110 - 0x6e
    "01100111", -- 7270 - 0x1c66  :  103 - 0x67
    "00000000", -- 7271 - 0x1c67  :    0 - 0x0
    "01111110", -- 7272 - 0x1c68  :  126 - 0x7e
    "01100011", -- 7273 - 0x1c69  :   99 - 0x63
    "01100011", -- 7274 - 0x1c6a  :   99 - 0x63
    "01100111", -- 7275 - 0x1c6b  :  103 - 0x67
    "01111100", -- 7276 - 0x1c6c  :  124 - 0x7c
    "01101110", -- 7277 - 0x1c6d  :  110 - 0x6e
    "01100111", -- 7278 - 0x1c6e  :  103 - 0x67
    "00000000", -- 7279 - 0x1c6f  :    0 - 0x0
    "01111111", -- 7280 - 0x1c70  :  127 - 0x7f -- Background 0xc7
    "01100000", -- 7281 - 0x1c71  :   96 - 0x60
    "01100000", -- 7282 - 0x1c72  :   96 - 0x60
    "01111110", -- 7283 - 0x1c73  :  126 - 0x7e
    "01100000", -- 7284 - 0x1c74  :   96 - 0x60
    "01100000", -- 7285 - 0x1c75  :   96 - 0x60
    "01111111", -- 7286 - 0x1c76  :  127 - 0x7f
    "00000000", -- 7287 - 0x1c77  :    0 - 0x0
    "01111111", -- 7288 - 0x1c78  :  127 - 0x7f
    "01100000", -- 7289 - 0x1c79  :   96 - 0x60
    "01100000", -- 7290 - 0x1c7a  :   96 - 0x60
    "01111110", -- 7291 - 0x1c7b  :  126 - 0x7e
    "01100000", -- 7292 - 0x1c7c  :   96 - 0x60
    "01100000", -- 7293 - 0x1c7d  :   96 - 0x60
    "01111111", -- 7294 - 0x1c7e  :  127 - 0x7f
    "00000000", -- 7295 - 0x1c7f  :    0 - 0x0
    "00110110", -- 7296 - 0x1c80  :   54 - 0x36 -- Background 0xc8
    "00110110", -- 7297 - 0x1c81  :   54 - 0x36
    "00010010", -- 7298 - 0x1c82  :   18 - 0x12
    "00000000", -- 7299 - 0x1c83  :    0 - 0x0
    "00000000", -- 7300 - 0x1c84  :    0 - 0x0
    "00000000", -- 7301 - 0x1c85  :    0 - 0x0
    "00000000", -- 7302 - 0x1c86  :    0 - 0x0
    "00000000", -- 7303 - 0x1c87  :    0 - 0x0
    "00110110", -- 7304 - 0x1c88  :   54 - 0x36
    "00110110", -- 7305 - 0x1c89  :   54 - 0x36
    "00010010", -- 7306 - 0x1c8a  :   18 - 0x12
    "00000000", -- 7307 - 0x1c8b  :    0 - 0x0
    "00000000", -- 7308 - 0x1c8c  :    0 - 0x0
    "00000000", -- 7309 - 0x1c8d  :    0 - 0x0
    "00000000", -- 7310 - 0x1c8e  :    0 - 0x0
    "00000000", -- 7311 - 0x1c8f  :    0 - 0x0
    "00111110", -- 7312 - 0x1c90  :   62 - 0x3e -- Background 0xc9
    "01100011", -- 7313 - 0x1c91  :   99 - 0x63
    "01100011", -- 7314 - 0x1c92  :   99 - 0x63
    "01100011", -- 7315 - 0x1c93  :   99 - 0x63
    "01100011", -- 7316 - 0x1c94  :   99 - 0x63
    "01100011", -- 7317 - 0x1c95  :   99 - 0x63
    "00111110", -- 7318 - 0x1c96  :   62 - 0x3e
    "00000000", -- 7319 - 0x1c97  :    0 - 0x0
    "00111110", -- 7320 - 0x1c98  :   62 - 0x3e
    "01100011", -- 7321 - 0x1c99  :   99 - 0x63
    "01100011", -- 7322 - 0x1c9a  :   99 - 0x63
    "01100011", -- 7323 - 0x1c9b  :   99 - 0x63
    "01100011", -- 7324 - 0x1c9c  :   99 - 0x63
    "01100011", -- 7325 - 0x1c9d  :   99 - 0x63
    "00111110", -- 7326 - 0x1c9e  :   62 - 0x3e
    "00000000", -- 7327 - 0x1c9f  :    0 - 0x0
    "00111100", -- 7328 - 0x1ca0  :   60 - 0x3c -- Background 0xca
    "01100110", -- 7329 - 0x1ca1  :  102 - 0x66
    "01100000", -- 7330 - 0x1ca2  :   96 - 0x60
    "00111110", -- 7331 - 0x1ca3  :   62 - 0x3e
    "00000011", -- 7332 - 0x1ca4  :    3 - 0x3
    "01100011", -- 7333 - 0x1ca5  :   99 - 0x63
    "00111110", -- 7334 - 0x1ca6  :   62 - 0x3e
    "00000000", -- 7335 - 0x1ca7  :    0 - 0x0
    "00111100", -- 7336 - 0x1ca8  :   60 - 0x3c
    "01100110", -- 7337 - 0x1ca9  :  102 - 0x66
    "01100000", -- 7338 - 0x1caa  :   96 - 0x60
    "00111110", -- 7339 - 0x1cab  :   62 - 0x3e
    "00000011", -- 7340 - 0x1cac  :    3 - 0x3
    "01100011", -- 7341 - 0x1cad  :   99 - 0x63
    "00111110", -- 7342 - 0x1cae  :   62 - 0x3e
    "00000000", -- 7343 - 0x1caf  :    0 - 0x0
    "00000000", -- 7344 - 0x1cb0  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 7345 - 0x1cb1  :    0 - 0x0
    "00000000", -- 7346 - 0x1cb2  :    0 - 0x0
    "00000000", -- 7347 - 0x1cb3  :    0 - 0x0
    "00000000", -- 7348 - 0x1cb4  :    0 - 0x0
    "00000000", -- 7349 - 0x1cb5  :    0 - 0x0
    "00000000", -- 7350 - 0x1cb6  :    0 - 0x0
    "00000000", -- 7351 - 0x1cb7  :    0 - 0x0
    "00000000", -- 7352 - 0x1cb8  :    0 - 0x0
    "00111000", -- 7353 - 0x1cb9  :   56 - 0x38
    "01111100", -- 7354 - 0x1cba  :  124 - 0x7c
    "11111110", -- 7355 - 0x1cbb  :  254 - 0xfe
    "11111110", -- 7356 - 0x1cbc  :  254 - 0xfe
    "11111110", -- 7357 - 0x1cbd  :  254 - 0xfe
    "01111100", -- 7358 - 0x1cbe  :  124 - 0x7c
    "00111000", -- 7359 - 0x1cbf  :   56 - 0x38
    "00000000", -- 7360 - 0x1cc0  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 7361 - 0x1cc1  :    0 - 0x0
    "00000000", -- 7362 - 0x1cc2  :    0 - 0x0
    "00000000", -- 7363 - 0x1cc3  :    0 - 0x0
    "00000000", -- 7364 - 0x1cc4  :    0 - 0x0
    "00000000", -- 7365 - 0x1cc5  :    0 - 0x0
    "00000000", -- 7366 - 0x1cc6  :    0 - 0x0
    "00000000", -- 7367 - 0x1cc7  :    0 - 0x0
    "00000000", -- 7368 - 0x1cc8  :    0 - 0x0
    "00000000", -- 7369 - 0x1cc9  :    0 - 0x0
    "00000000", -- 7370 - 0x1cca  :    0 - 0x0
    "00000000", -- 7371 - 0x1ccb  :    0 - 0x0
    "00000000", -- 7372 - 0x1ccc  :    0 - 0x0
    "00000000", -- 7373 - 0x1ccd  :    0 - 0x0
    "00000000", -- 7374 - 0x1cce  :    0 - 0x0
    "00000000", -- 7375 - 0x1ccf  :    0 - 0x0
    "00000000", -- 7376 - 0x1cd0  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 7377 - 0x1cd1  :    0 - 0x0
    "00000000", -- 7378 - 0x1cd2  :    0 - 0x0
    "00000000", -- 7379 - 0x1cd3  :    0 - 0x0
    "00000000", -- 7380 - 0x1cd4  :    0 - 0x0
    "00000000", -- 7381 - 0x1cd5  :    0 - 0x0
    "00000000", -- 7382 - 0x1cd6  :    0 - 0x0
    "00000000", -- 7383 - 0x1cd7  :    0 - 0x0
    "00000000", -- 7384 - 0x1cd8  :    0 - 0x0
    "00000000", -- 7385 - 0x1cd9  :    0 - 0x0
    "00000000", -- 7386 - 0x1cda  :    0 - 0x0
    "00000000", -- 7387 - 0x1cdb  :    0 - 0x0
    "00000000", -- 7388 - 0x1cdc  :    0 - 0x0
    "00000000", -- 7389 - 0x1cdd  :    0 - 0x0
    "00000000", -- 7390 - 0x1cde  :    0 - 0x0
    "00000000", -- 7391 - 0x1cdf  :    0 - 0x0
    "00000000", -- 7392 - 0x1ce0  :    0 - 0x0 -- Background 0xce
    "00000000", -- 7393 - 0x1ce1  :    0 - 0x0
    "00000000", -- 7394 - 0x1ce2  :    0 - 0x0
    "00000000", -- 7395 - 0x1ce3  :    0 - 0x0
    "00000000", -- 7396 - 0x1ce4  :    0 - 0x0
    "00000000", -- 7397 - 0x1ce5  :    0 - 0x0
    "00000000", -- 7398 - 0x1ce6  :    0 - 0x0
    "00000000", -- 7399 - 0x1ce7  :    0 - 0x0
    "00000000", -- 7400 - 0x1ce8  :    0 - 0x0
    "00000000", -- 7401 - 0x1ce9  :    0 - 0x0
    "00000000", -- 7402 - 0x1cea  :    0 - 0x0
    "00000000", -- 7403 - 0x1ceb  :    0 - 0x0
    "00000000", -- 7404 - 0x1cec  :    0 - 0x0
    "00000000", -- 7405 - 0x1ced  :    0 - 0x0
    "00000000", -- 7406 - 0x1cee  :    0 - 0x0
    "00000000", -- 7407 - 0x1cef  :    0 - 0x0
    "00000000", -- 7408 - 0x1cf0  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 7409 - 0x1cf1  :    0 - 0x0
    "00000000", -- 7410 - 0x1cf2  :    0 - 0x0
    "00000000", -- 7411 - 0x1cf3  :    0 - 0x0
    "00000000", -- 7412 - 0x1cf4  :    0 - 0x0
    "00000000", -- 7413 - 0x1cf5  :    0 - 0x0
    "00000000", -- 7414 - 0x1cf6  :    0 - 0x0
    "00000000", -- 7415 - 0x1cf7  :    0 - 0x0
    "00000000", -- 7416 - 0x1cf8  :    0 - 0x0
    "00000000", -- 7417 - 0x1cf9  :    0 - 0x0
    "00000000", -- 7418 - 0x1cfa  :    0 - 0x0
    "00000000", -- 7419 - 0x1cfb  :    0 - 0x0
    "00000000", -- 7420 - 0x1cfc  :    0 - 0x0
    "00000000", -- 7421 - 0x1cfd  :    0 - 0x0
    "00000000", -- 7422 - 0x1cfe  :    0 - 0x0
    "00000000", -- 7423 - 0x1cff  :    0 - 0x0
    "01000111", -- 7424 - 0x1d00  :   71 - 0x47 -- Background 0xd0
    "01000111", -- 7425 - 0x1d01  :   71 - 0x47
    "00001111", -- 7426 - 0x1d02  :   15 - 0xf
    "00001111", -- 7427 - 0x1d03  :   15 - 0xf
    "00011111", -- 7428 - 0x1d04  :   31 - 0x1f
    "00011111", -- 7429 - 0x1d05  :   31 - 0x1f
    "00111111", -- 7430 - 0x1d06  :   63 - 0x3f
    "00111111", -- 7431 - 0x1d07  :   63 - 0x3f
    "00010111", -- 7432 - 0x1d08  :   23 - 0x17
    "00010111", -- 7433 - 0x1d09  :   23 - 0x17
    "00101111", -- 7434 - 0x1d0a  :   47 - 0x2f
    "00101111", -- 7435 - 0x1d0b  :   47 - 0x2f
    "01011111", -- 7436 - 0x1d0c  :   95 - 0x5f
    "01011111", -- 7437 - 0x1d0d  :   95 - 0x5f
    "00111111", -- 7438 - 0x1d0e  :   63 - 0x3f
    "00111111", -- 7439 - 0x1d0f  :   63 - 0x3f
    "11111111", -- 7440 - 0x1d10  :  255 - 0xff -- Background 0xd1
    "11001111", -- 7441 - 0x1d11  :  207 - 0xcf
    "11001111", -- 7442 - 0x1d12  :  207 - 0xcf
    "11111011", -- 7443 - 0x1d13  :  251 - 0xfb
    "11110111", -- 7444 - 0x1d14  :  247 - 0xf7
    "11100111", -- 7445 - 0x1d15  :  231 - 0xe7
    "11111111", -- 7446 - 0x1d16  :  255 - 0xff
    "11111111", -- 7447 - 0x1d17  :  255 - 0xff
    "11111111", -- 7448 - 0x1d18  :  255 - 0xff
    "11001111", -- 7449 - 0x1d19  :  207 - 0xcf
    "11001111", -- 7450 - 0x1d1a  :  207 - 0xcf
    "11111011", -- 7451 - 0x1d1b  :  251 - 0xfb
    "11110111", -- 7452 - 0x1d1c  :  247 - 0xf7
    "11100111", -- 7453 - 0x1d1d  :  231 - 0xe7
    "11111111", -- 7454 - 0x1d1e  :  255 - 0xff
    "11111111", -- 7455 - 0x1d1f  :  255 - 0xff
    "00011000", -- 7456 - 0x1d20  :   24 - 0x18 -- Background 0xd2
    "00001000", -- 7457 - 0x1d21  :    8 - 0x8
    "10001000", -- 7458 - 0x1d22  :  136 - 0x88
    "10000000", -- 7459 - 0x1d23  :  128 - 0x80
    "01000000", -- 7460 - 0x1d24  :   64 - 0x40
    "01000000", -- 7461 - 0x1d25  :   64 - 0x40
    "10100000", -- 7462 - 0x1d26  :  160 - 0xa0
    "10100000", -- 7463 - 0x1d27  :  160 - 0xa0
    "01000010", -- 7464 - 0x1d28  :   66 - 0x42
    "01100010", -- 7465 - 0x1d29  :   98 - 0x62
    "10100010", -- 7466 - 0x1d2a  :  162 - 0xa2
    "10110010", -- 7467 - 0x1d2b  :  178 - 0xb2
    "01010010", -- 7468 - 0x1d2c  :   82 - 0x52
    "01011010", -- 7469 - 0x1d2d  :   90 - 0x5a
    "10101010", -- 7470 - 0x1d2e  :  170 - 0xaa
    "10101100", -- 7471 - 0x1d2f  :  172 - 0xac
    "11111111", -- 7472 - 0x1d30  :  255 - 0xff -- Background 0xd3
    "11111111", -- 7473 - 0x1d31  :  255 - 0xff
    "11111111", -- 7474 - 0x1d32  :  255 - 0xff
    "11111111", -- 7475 - 0x1d33  :  255 - 0xff
    "11111101", -- 7476 - 0x1d34  :  253 - 0xfd
    "11111101", -- 7477 - 0x1d35  :  253 - 0xfd
    "11111101", -- 7478 - 0x1d36  :  253 - 0xfd
    "11111101", -- 7479 - 0x1d37  :  253 - 0xfd
    "11111111", -- 7480 - 0x1d38  :  255 - 0xff
    "11111111", -- 7481 - 0x1d39  :  255 - 0xff
    "11111111", -- 7482 - 0x1d3a  :  255 - 0xff
    "11111111", -- 7483 - 0x1d3b  :  255 - 0xff
    "11111101", -- 7484 - 0x1d3c  :  253 - 0xfd
    "11111101", -- 7485 - 0x1d3d  :  253 - 0xfd
    "11111101", -- 7486 - 0x1d3e  :  253 - 0xfd
    "11111101", -- 7487 - 0x1d3f  :  253 - 0xfd
    "11000111", -- 7488 - 0x1d40  :  199 - 0xc7 -- Background 0xd4
    "11110111", -- 7489 - 0x1d41  :  247 - 0xf7
    "11110000", -- 7490 - 0x1d42  :  240 - 0xf0
    "11111000", -- 7491 - 0x1d43  :  248 - 0xf8
    "11111000", -- 7492 - 0x1d44  :  248 - 0xf8
    "11111111", -- 7493 - 0x1d45  :  255 - 0xff
    "11111111", -- 7494 - 0x1d46  :  255 - 0xff
    "11111111", -- 7495 - 0x1d47  :  255 - 0xff
    "00000111", -- 7496 - 0x1d48  :    7 - 0x7
    "00000111", -- 7497 - 0x1d49  :    7 - 0x7
    "00000000", -- 7498 - 0x1d4a  :    0 - 0x0
    "00000011", -- 7499 - 0x1d4b  :    3 - 0x3
    "00000000", -- 7500 - 0x1d4c  :    0 - 0x0
    "00000000", -- 7501 - 0x1d4d  :    0 - 0x0
    "00000000", -- 7502 - 0x1d4e  :    0 - 0x0
    "00000000", -- 7503 - 0x1d4f  :    0 - 0x0
    "11111000", -- 7504 - 0x1d50  :  248 - 0xf8 -- Background 0xd5
    "11111000", -- 7505 - 0x1d51  :  248 - 0xf8
    "00000000", -- 7506 - 0x1d52  :    0 - 0x0
    "00000000", -- 7507 - 0x1d53  :    0 - 0x0
    "00000000", -- 7508 - 0x1d54  :    0 - 0x0
    "11111111", -- 7509 - 0x1d55  :  255 - 0xff
    "11111111", -- 7510 - 0x1d56  :  255 - 0xff
    "11111111", -- 7511 - 0x1d57  :  255 - 0xff
    "11111010", -- 7512 - 0x1d58  :  250 - 0xfa
    "11111010", -- 7513 - 0x1d59  :  250 - 0xfa
    "00000010", -- 7514 - 0x1d5a  :    2 - 0x2
    "11111110", -- 7515 - 0x1d5b  :  254 - 0xfe
    "00000000", -- 7516 - 0x1d5c  :    0 - 0x0
    "00000000", -- 7517 - 0x1d5d  :    0 - 0x0
    "00000000", -- 7518 - 0x1d5e  :    0 - 0x0
    "00000000", -- 7519 - 0x1d5f  :    0 - 0x0
    "10001111", -- 7520 - 0x1d60  :  143 - 0x8f -- Background 0xd6
    "11101111", -- 7521 - 0x1d61  :  239 - 0xef
    "11000000", -- 7522 - 0x1d62  :  192 - 0xc0
    "11110000", -- 7523 - 0x1d63  :  240 - 0xf0
    "11100000", -- 7524 - 0x1d64  :  224 - 0xe0
    "11111111", -- 7525 - 0x1d65  :  255 - 0xff
    "11111111", -- 7526 - 0x1d66  :  255 - 0xff
    "11111111", -- 7527 - 0x1d67  :  255 - 0xff
    "00001111", -- 7528 - 0x1d68  :   15 - 0xf
    "00001111", -- 7529 - 0x1d69  :   15 - 0xf
    "00000000", -- 7530 - 0x1d6a  :    0 - 0x0
    "00000111", -- 7531 - 0x1d6b  :    7 - 0x7
    "00000000", -- 7532 - 0x1d6c  :    0 - 0x0
    "00000000", -- 7533 - 0x1d6d  :    0 - 0x0
    "00000000", -- 7534 - 0x1d6e  :    0 - 0x0
    "00000000", -- 7535 - 0x1d6f  :    0 - 0x0
    "11111111", -- 7536 - 0x1d70  :  255 - 0xff -- Background 0xd7
    "11111111", -- 7537 - 0x1d71  :  255 - 0xff
    "00000000", -- 7538 - 0x1d72  :    0 - 0x0
    "00000000", -- 7539 - 0x1d73  :    0 - 0x0
    "00000000", -- 7540 - 0x1d74  :    0 - 0x0
    "11111111", -- 7541 - 0x1d75  :  255 - 0xff
    "11111111", -- 7542 - 0x1d76  :  255 - 0xff
    "11111111", -- 7543 - 0x1d77  :  255 - 0xff
    "11111111", -- 7544 - 0x1d78  :  255 - 0xff
    "11111111", -- 7545 - 0x1d79  :  255 - 0xff
    "00000000", -- 7546 - 0x1d7a  :    0 - 0x0
    "11111111", -- 7547 - 0x1d7b  :  255 - 0xff
    "00000000", -- 7548 - 0x1d7c  :    0 - 0x0
    "00000000", -- 7549 - 0x1d7d  :    0 - 0x0
    "00000000", -- 7550 - 0x1d7e  :    0 - 0x0
    "00000000", -- 7551 - 0x1d7f  :    0 - 0x0
    "11000011", -- 7552 - 0x1d80  :  195 - 0xc3 -- Background 0xd8
    "11111111", -- 7553 - 0x1d81  :  255 - 0xff
    "00000000", -- 7554 - 0x1d82  :    0 - 0x0
    "00000000", -- 7555 - 0x1d83  :    0 - 0x0
    "00000000", -- 7556 - 0x1d84  :    0 - 0x0
    "11111111", -- 7557 - 0x1d85  :  255 - 0xff
    "11111111", -- 7558 - 0x1d86  :  255 - 0xff
    "11111111", -- 7559 - 0x1d87  :  255 - 0xff
    "11000011", -- 7560 - 0x1d88  :  195 - 0xc3
    "11111111", -- 7561 - 0x1d89  :  255 - 0xff
    "00000000", -- 7562 - 0x1d8a  :    0 - 0x0
    "11111111", -- 7563 - 0x1d8b  :  255 - 0xff
    "00000000", -- 7564 - 0x1d8c  :    0 - 0x0
    "00000000", -- 7565 - 0x1d8d  :    0 - 0x0
    "00000000", -- 7566 - 0x1d8e  :    0 - 0x0
    "00000000", -- 7567 - 0x1d8f  :    0 - 0x0
    "00000011", -- 7568 - 0x1d90  :    3 - 0x3 -- Background 0xd9
    "10000001", -- 7569 - 0x1d91  :  129 - 0x81
    "00000000", -- 7570 - 0x1d92  :    0 - 0x0
    "00000000", -- 7571 - 0x1d93  :    0 - 0x0
    "00000011", -- 7572 - 0x1d94  :    3 - 0x3
    "11111111", -- 7573 - 0x1d95  :  255 - 0xff
    "11111111", -- 7574 - 0x1d96  :  255 - 0xff
    "11111111", -- 7575 - 0x1d97  :  255 - 0xff
    "01101011", -- 7576 - 0x1d98  :  107 - 0x6b
    "10110101", -- 7577 - 0x1d99  :  181 - 0xb5
    "00110110", -- 7578 - 0x1d9a  :   54 - 0x36
    "11111000", -- 7579 - 0x1d9b  :  248 - 0xf8
    "00000000", -- 7580 - 0x1d9c  :    0 - 0x0
    "00000000", -- 7581 - 0x1d9d  :    0 - 0x0
    "00000000", -- 7582 - 0x1d9e  :    0 - 0x0
    "00000000", -- 7583 - 0x1d9f  :    0 - 0x0
    "11111111", -- 7584 - 0x1da0  :  255 - 0xff -- Background 0xda
    "11111111", -- 7585 - 0x1da1  :  255 - 0xff
    "01111110", -- 7586 - 0x1da2  :  126 - 0x7e
    "00000000", -- 7587 - 0x1da3  :    0 - 0x0
    "00000000", -- 7588 - 0x1da4  :    0 - 0x0
    "11100000", -- 7589 - 0x1da5  :  224 - 0xe0
    "11111111", -- 7590 - 0x1da6  :  255 - 0xff
    "11111111", -- 7591 - 0x1da7  :  255 - 0xff
    "11111111", -- 7592 - 0x1da8  :  255 - 0xff
    "11111111", -- 7593 - 0x1da9  :  255 - 0xff
    "01111110", -- 7594 - 0x1daa  :  126 - 0x7e
    "10000001", -- 7595 - 0x1dab  :  129 - 0x81
    "00011111", -- 7596 - 0x1dac  :   31 - 0x1f
    "00000000", -- 7597 - 0x1dad  :    0 - 0x0
    "00000000", -- 7598 - 0x1dae  :    0 - 0x0
    "00000000", -- 7599 - 0x1daf  :    0 - 0x0
    "01100001", -- 7600 - 0x1db0  :   97 - 0x61 -- Background 0xdb
    "11000011", -- 7601 - 0x1db1  :  195 - 0xc3
    "00000111", -- 7602 - 0x1db2  :    7 - 0x7
    "00001111", -- 7603 - 0x1db3  :   15 - 0xf
    "00011111", -- 7604 - 0x1db4  :   31 - 0x1f
    "01111111", -- 7605 - 0x1db5  :  127 - 0x7f
    "11111111", -- 7606 - 0x1db6  :  255 - 0xff
    "11111111", -- 7607 - 0x1db7  :  255 - 0xff
    "01101100", -- 7608 - 0x1db8  :  108 - 0x6c
    "11011000", -- 7609 - 0x1db9  :  216 - 0xd8
    "00110000", -- 7610 - 0x1dba  :   48 - 0x30
    "11100000", -- 7611 - 0x1dbb  :  224 - 0xe0
    "10000000", -- 7612 - 0x1dbc  :  128 - 0x80
    "00000000", -- 7613 - 0x1dbd  :    0 - 0x0
    "00000000", -- 7614 - 0x1dbe  :    0 - 0x0
    "00000000", -- 7615 - 0x1dbf  :    0 - 0x0
    "00011111", -- 7616 - 0x1dc0  :   31 - 0x1f -- Background 0xdc
    "11011111", -- 7617 - 0x1dc1  :  223 - 0xdf
    "11000000", -- 7618 - 0x1dc2  :  192 - 0xc0
    "11110000", -- 7619 - 0x1dc3  :  240 - 0xf0
    "11110000", -- 7620 - 0x1dc4  :  240 - 0xf0
    "11111111", -- 7621 - 0x1dc5  :  255 - 0xff
    "11111111", -- 7622 - 0x1dc6  :  255 - 0xff
    "11111111", -- 7623 - 0x1dc7  :  255 - 0xff
    "00011111", -- 7624 - 0x1dc8  :   31 - 0x1f
    "00011111", -- 7625 - 0x1dc9  :   31 - 0x1f
    "00000000", -- 7626 - 0x1dca  :    0 - 0x0
    "00000111", -- 7627 - 0x1dcb  :    7 - 0x7
    "00000000", -- 7628 - 0x1dcc  :    0 - 0x0
    "00000000", -- 7629 - 0x1dcd  :    0 - 0x0
    "00000000", -- 7630 - 0x1dce  :    0 - 0x0
    "00000000", -- 7631 - 0x1dcf  :    0 - 0x0
    "10000100", -- 7632 - 0x1dd0  :  132 - 0x84 -- Background 0xdd
    "11111100", -- 7633 - 0x1dd1  :  252 - 0xfc
    "00000000", -- 7634 - 0x1dd2  :    0 - 0x0
    "00000000", -- 7635 - 0x1dd3  :    0 - 0x0
    "00000000", -- 7636 - 0x1dd4  :    0 - 0x0
    "11111111", -- 7637 - 0x1dd5  :  255 - 0xff
    "11111111", -- 7638 - 0x1dd6  :  255 - 0xff
    "11111111", -- 7639 - 0x1dd7  :  255 - 0xff
    "10000101", -- 7640 - 0x1dd8  :  133 - 0x85
    "11111101", -- 7641 - 0x1dd9  :  253 - 0xfd
    "00000001", -- 7642 - 0x1dda  :    1 - 0x1
    "11111111", -- 7643 - 0x1ddb  :  255 - 0xff
    "00000000", -- 7644 - 0x1ddc  :    0 - 0x0
    "00000000", -- 7645 - 0x1ddd  :    0 - 0x0
    "00000000", -- 7646 - 0x1dde  :    0 - 0x0
    "00000000", -- 7647 - 0x1ddf  :    0 - 0x0
    "01111111", -- 7648 - 0x1de0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 7649 - 0x1de1  :  127 - 0x7f
    "00000000", -- 7650 - 0x1de2  :    0 - 0x0
    "00000000", -- 7651 - 0x1de3  :    0 - 0x0
    "00000000", -- 7652 - 0x1de4  :    0 - 0x0
    "11111111", -- 7653 - 0x1de5  :  255 - 0xff
    "11111111", -- 7654 - 0x1de6  :  255 - 0xff
    "11111111", -- 7655 - 0x1de7  :  255 - 0xff
    "01111111", -- 7656 - 0x1de8  :  127 - 0x7f
    "01111111", -- 7657 - 0x1de9  :  127 - 0x7f
    "00000000", -- 7658 - 0x1dea  :    0 - 0x0
    "01011111", -- 7659 - 0x1deb  :   95 - 0x5f
    "00000000", -- 7660 - 0x1dec  :    0 - 0x0
    "00000000", -- 7661 - 0x1ded  :    0 - 0x0
    "00000000", -- 7662 - 0x1dee  :    0 - 0x0
    "00000000", -- 7663 - 0x1def  :    0 - 0x0
    "11111100", -- 7664 - 0x1df0  :  252 - 0xfc -- Background 0xdf
    "11111111", -- 7665 - 0x1df1  :  255 - 0xff
    "00000000", -- 7666 - 0x1df2  :    0 - 0x0
    "00000000", -- 7667 - 0x1df3  :    0 - 0x0
    "00000000", -- 7668 - 0x1df4  :    0 - 0x0
    "11111111", -- 7669 - 0x1df5  :  255 - 0xff
    "11111111", -- 7670 - 0x1df6  :  255 - 0xff
    "11111111", -- 7671 - 0x1df7  :  255 - 0xff
    "11111100", -- 7672 - 0x1df8  :  252 - 0xfc
    "11111111", -- 7673 - 0x1df9  :  255 - 0xff
    "00000000", -- 7674 - 0x1dfa  :    0 - 0x0
    "11111111", -- 7675 - 0x1dfb  :  255 - 0xff
    "00000000", -- 7676 - 0x1dfc  :    0 - 0x0
    "00000000", -- 7677 - 0x1dfd  :    0 - 0x0
    "00000000", -- 7678 - 0x1dfe  :    0 - 0x0
    "00000000", -- 7679 - 0x1dff  :    0 - 0x0
    "00110000", -- 7680 - 0x1e00  :   48 - 0x30 -- Background 0xe0
    "11110000", -- 7681 - 0x1e01  :  240 - 0xf0
    "00000000", -- 7682 - 0x1e02  :    0 - 0x0
    "00000000", -- 7683 - 0x1e03  :    0 - 0x0
    "00000000", -- 7684 - 0x1e04  :    0 - 0x0
    "11111111", -- 7685 - 0x1e05  :  255 - 0xff
    "11111111", -- 7686 - 0x1e06  :  255 - 0xff
    "11111111", -- 7687 - 0x1e07  :  255 - 0xff
    "00110100", -- 7688 - 0x1e08  :   52 - 0x34
    "11110110", -- 7689 - 0x1e09  :  246 - 0xf6
    "00000010", -- 7690 - 0x1e0a  :    2 - 0x2
    "11111111", -- 7691 - 0x1e0b  :  255 - 0xff
    "00000000", -- 7692 - 0x1e0c  :    0 - 0x0
    "00000000", -- 7693 - 0x1e0d  :    0 - 0x0
    "00000000", -- 7694 - 0x1e0e  :    0 - 0x0
    "00000000", -- 7695 - 0x1e0f  :    0 - 0x0
    "11111111", -- 7696 - 0x1e10  :  255 - 0xff -- Background 0xe1
    "11111111", -- 7697 - 0x1e11  :  255 - 0xff
    "00000000", -- 7698 - 0x1e12  :    0 - 0x0
    "00000000", -- 7699 - 0x1e13  :    0 - 0x0
    "00000000", -- 7700 - 0x1e14  :    0 - 0x0
    "11111111", -- 7701 - 0x1e15  :  255 - 0xff
    "11111111", -- 7702 - 0x1e16  :  255 - 0xff
    "11111111", -- 7703 - 0x1e17  :  255 - 0xff
    "11111111", -- 7704 - 0x1e18  :  255 - 0xff
    "11111111", -- 7705 - 0x1e19  :  255 - 0xff
    "00000000", -- 7706 - 0x1e1a  :    0 - 0x0
    "01111111", -- 7707 - 0x1e1b  :  127 - 0x7f
    "00000000", -- 7708 - 0x1e1c  :    0 - 0x0
    "00000000", -- 7709 - 0x1e1d  :    0 - 0x0
    "00000000", -- 7710 - 0x1e1e  :    0 - 0x0
    "00000000", -- 7711 - 0x1e1f  :    0 - 0x0
    "11100001", -- 7712 - 0x1e20  :  225 - 0xe1 -- Background 0xe2
    "11111111", -- 7713 - 0x1e21  :  255 - 0xff
    "00000000", -- 7714 - 0x1e22  :    0 - 0x0
    "00000000", -- 7715 - 0x1e23  :    0 - 0x0
    "00000000", -- 7716 - 0x1e24  :    0 - 0x0
    "11111111", -- 7717 - 0x1e25  :  255 - 0xff
    "11111111", -- 7718 - 0x1e26  :  255 - 0xff
    "11111111", -- 7719 - 0x1e27  :  255 - 0xff
    "11100001", -- 7720 - 0x1e28  :  225 - 0xe1
    "11111111", -- 7721 - 0x1e29  :  255 - 0xff
    "00000000", -- 7722 - 0x1e2a  :    0 - 0x0
    "11111111", -- 7723 - 0x1e2b  :  255 - 0xff
    "00000000", -- 7724 - 0x1e2c  :    0 - 0x0
    "00000000", -- 7725 - 0x1e2d  :    0 - 0x0
    "00000000", -- 7726 - 0x1e2e  :    0 - 0x0
    "00000000", -- 7727 - 0x1e2f  :    0 - 0x0
    "00011111", -- 7728 - 0x1e30  :   31 - 0x1f -- Background 0xe3
    "00011111", -- 7729 - 0x1e31  :   31 - 0x1f
    "00011111", -- 7730 - 0x1e32  :   31 - 0x1f
    "00011111", -- 7731 - 0x1e33  :   31 - 0x1f
    "00011111", -- 7732 - 0x1e34  :   31 - 0x1f
    "11111111", -- 7733 - 0x1e35  :  255 - 0xff
    "11111111", -- 7734 - 0x1e36  :  255 - 0xff
    "11111111", -- 7735 - 0x1e37  :  255 - 0xff
    "01000000", -- 7736 - 0x1e38  :   64 - 0x40
    "01000000", -- 7737 - 0x1e39  :   64 - 0x40
    "01000000", -- 7738 - 0x1e3a  :   64 - 0x40
    "11000000", -- 7739 - 0x1e3b  :  192 - 0xc0
    "00000000", -- 7740 - 0x1e3c  :    0 - 0x0
    "00000000", -- 7741 - 0x1e3d  :    0 - 0x0
    "00000000", -- 7742 - 0x1e3e  :    0 - 0x0
    "00000000", -- 7743 - 0x1e3f  :    0 - 0x0
    "00000000", -- 7744 - 0x1e40  :    0 - 0x0 -- Background 0xe4
    "00011111", -- 7745 - 0x1e41  :   31 - 0x1f
    "00111111", -- 7746 - 0x1e42  :   63 - 0x3f
    "01111000", -- 7747 - 0x1e43  :  120 - 0x78
    "01110111", -- 7748 - 0x1e44  :  119 - 0x77
    "01101111", -- 7749 - 0x1e45  :  111 - 0x6f
    "01101111", -- 7750 - 0x1e46  :  111 - 0x6f
    "01101111", -- 7751 - 0x1e47  :  111 - 0x6f
    "00000000", -- 7752 - 0x1e48  :    0 - 0x0
    "00000000", -- 7753 - 0x1e49  :    0 - 0x0
    "00000000", -- 7754 - 0x1e4a  :    0 - 0x0
    "00000000", -- 7755 - 0x1e4b  :    0 - 0x0
    "00000111", -- 7756 - 0x1e4c  :    7 - 0x7
    "00001111", -- 7757 - 0x1e4d  :   15 - 0xf
    "00001111", -- 7758 - 0x1e4e  :   15 - 0xf
    "00001111", -- 7759 - 0x1e4f  :   15 - 0xf
    "00000000", -- 7760 - 0x1e50  :    0 - 0x0 -- Background 0xe5
    "11111000", -- 7761 - 0x1e51  :  248 - 0xf8
    "11111100", -- 7762 - 0x1e52  :  252 - 0xfc
    "00011110", -- 7763 - 0x1e53  :   30 - 0x1e
    "11101110", -- 7764 - 0x1e54  :  238 - 0xee
    "11110110", -- 7765 - 0x1e55  :  246 - 0xf6
    "11110110", -- 7766 - 0x1e56  :  246 - 0xf6
    "11110110", -- 7767 - 0x1e57  :  246 - 0xf6
    "00000000", -- 7768 - 0x1e58  :    0 - 0x0
    "00000000", -- 7769 - 0x1e59  :    0 - 0x0
    "00000000", -- 7770 - 0x1e5a  :    0 - 0x0
    "00000000", -- 7771 - 0x1e5b  :    0 - 0x0
    "11100000", -- 7772 - 0x1e5c  :  224 - 0xe0
    "11110000", -- 7773 - 0x1e5d  :  240 - 0xf0
    "11110000", -- 7774 - 0x1e5e  :  240 - 0xf0
    "11110000", -- 7775 - 0x1e5f  :  240 - 0xf0
    "11110110", -- 7776 - 0x1e60  :  246 - 0xf6 -- Background 0xe6
    "11110110", -- 7777 - 0x1e61  :  246 - 0xf6
    "11110110", -- 7778 - 0x1e62  :  246 - 0xf6
    "11101110", -- 7779 - 0x1e63  :  238 - 0xee
    "00011110", -- 7780 - 0x1e64  :   30 - 0x1e
    "11111100", -- 7781 - 0x1e65  :  252 - 0xfc
    "11111000", -- 7782 - 0x1e66  :  248 - 0xf8
    "00000000", -- 7783 - 0x1e67  :    0 - 0x0
    "11110000", -- 7784 - 0x1e68  :  240 - 0xf0
    "11110000", -- 7785 - 0x1e69  :  240 - 0xf0
    "11110000", -- 7786 - 0x1e6a  :  240 - 0xf0
    "11100000", -- 7787 - 0x1e6b  :  224 - 0xe0
    "00000000", -- 7788 - 0x1e6c  :    0 - 0x0
    "00000000", -- 7789 - 0x1e6d  :    0 - 0x0
    "00000000", -- 7790 - 0x1e6e  :    0 - 0x0
    "00000000", -- 7791 - 0x1e6f  :    0 - 0x0
    "01101111", -- 7792 - 0x1e70  :  111 - 0x6f -- Background 0xe7
    "01101111", -- 7793 - 0x1e71  :  111 - 0x6f
    "01101111", -- 7794 - 0x1e72  :  111 - 0x6f
    "01110111", -- 7795 - 0x1e73  :  119 - 0x77
    "01111000", -- 7796 - 0x1e74  :  120 - 0x78
    "00111111", -- 7797 - 0x1e75  :   63 - 0x3f
    "00011111", -- 7798 - 0x1e76  :   31 - 0x1f
    "00000000", -- 7799 - 0x1e77  :    0 - 0x0
    "00001111", -- 7800 - 0x1e78  :   15 - 0xf
    "00001111", -- 7801 - 0x1e79  :   15 - 0xf
    "00001111", -- 7802 - 0x1e7a  :   15 - 0xf
    "00000111", -- 7803 - 0x1e7b  :    7 - 0x7
    "00000000", -- 7804 - 0x1e7c  :    0 - 0x0
    "00000000", -- 7805 - 0x1e7d  :    0 - 0x0
    "00000000", -- 7806 - 0x1e7e  :    0 - 0x0
    "00000000", -- 7807 - 0x1e7f  :    0 - 0x0
    "00000000", -- 7808 - 0x1e80  :    0 - 0x0 -- Background 0xe8
    "11111111", -- 7809 - 0x1e81  :  255 - 0xff
    "11111111", -- 7810 - 0x1e82  :  255 - 0xff
    "00000000", -- 7811 - 0x1e83  :    0 - 0x0
    "11111111", -- 7812 - 0x1e84  :  255 - 0xff
    "11111111", -- 7813 - 0x1e85  :  255 - 0xff
    "11111111", -- 7814 - 0x1e86  :  255 - 0xff
    "11111111", -- 7815 - 0x1e87  :  255 - 0xff
    "00000000", -- 7816 - 0x1e88  :    0 - 0x0
    "00000000", -- 7817 - 0x1e89  :    0 - 0x0
    "00000000", -- 7818 - 0x1e8a  :    0 - 0x0
    "00000000", -- 7819 - 0x1e8b  :    0 - 0x0
    "11111111", -- 7820 - 0x1e8c  :  255 - 0xff
    "11111111", -- 7821 - 0x1e8d  :  255 - 0xff
    "11111111", -- 7822 - 0x1e8e  :  255 - 0xff
    "11111111", -- 7823 - 0x1e8f  :  255 - 0xff
    "11110110", -- 7824 - 0x1e90  :  246 - 0xf6 -- Background 0xe9
    "11110110", -- 7825 - 0x1e91  :  246 - 0xf6
    "11110110", -- 7826 - 0x1e92  :  246 - 0xf6
    "11110110", -- 7827 - 0x1e93  :  246 - 0xf6
    "11110110", -- 7828 - 0x1e94  :  246 - 0xf6
    "11110110", -- 7829 - 0x1e95  :  246 - 0xf6
    "11110110", -- 7830 - 0x1e96  :  246 - 0xf6
    "11110110", -- 7831 - 0x1e97  :  246 - 0xf6
    "11110000", -- 7832 - 0x1e98  :  240 - 0xf0
    "11110000", -- 7833 - 0x1e99  :  240 - 0xf0
    "11110000", -- 7834 - 0x1e9a  :  240 - 0xf0
    "11110000", -- 7835 - 0x1e9b  :  240 - 0xf0
    "11110000", -- 7836 - 0x1e9c  :  240 - 0xf0
    "11110000", -- 7837 - 0x1e9d  :  240 - 0xf0
    "11110000", -- 7838 - 0x1e9e  :  240 - 0xf0
    "11110000", -- 7839 - 0x1e9f  :  240 - 0xf0
    "11111111", -- 7840 - 0x1ea0  :  255 - 0xff -- Background 0xea
    "11111111", -- 7841 - 0x1ea1  :  255 - 0xff
    "11111111", -- 7842 - 0x1ea2  :  255 - 0xff
    "11111111", -- 7843 - 0x1ea3  :  255 - 0xff
    "00000000", -- 7844 - 0x1ea4  :    0 - 0x0
    "11111111", -- 7845 - 0x1ea5  :  255 - 0xff
    "11111111", -- 7846 - 0x1ea6  :  255 - 0xff
    "00000000", -- 7847 - 0x1ea7  :    0 - 0x0
    "11111111", -- 7848 - 0x1ea8  :  255 - 0xff
    "11111111", -- 7849 - 0x1ea9  :  255 - 0xff
    "11111111", -- 7850 - 0x1eaa  :  255 - 0xff
    "11111111", -- 7851 - 0x1eab  :  255 - 0xff
    "00000000", -- 7852 - 0x1eac  :    0 - 0x0
    "00000000", -- 7853 - 0x1ead  :    0 - 0x0
    "00000000", -- 7854 - 0x1eae  :    0 - 0x0
    "00000000", -- 7855 - 0x1eaf  :    0 - 0x0
    "01101111", -- 7856 - 0x1eb0  :  111 - 0x6f -- Background 0xeb
    "01101111", -- 7857 - 0x1eb1  :  111 - 0x6f
    "01101111", -- 7858 - 0x1eb2  :  111 - 0x6f
    "01101111", -- 7859 - 0x1eb3  :  111 - 0x6f
    "01101111", -- 7860 - 0x1eb4  :  111 - 0x6f
    "01101111", -- 7861 - 0x1eb5  :  111 - 0x6f
    "01101111", -- 7862 - 0x1eb6  :  111 - 0x6f
    "01101111", -- 7863 - 0x1eb7  :  111 - 0x6f
    "00001111", -- 7864 - 0x1eb8  :   15 - 0xf
    "00001111", -- 7865 - 0x1eb9  :   15 - 0xf
    "00001111", -- 7866 - 0x1eba  :   15 - 0xf
    "00001111", -- 7867 - 0x1ebb  :   15 - 0xf
    "00001111", -- 7868 - 0x1ebc  :   15 - 0xf
    "00001111", -- 7869 - 0x1ebd  :   15 - 0xf
    "00001111", -- 7870 - 0x1ebe  :   15 - 0xf
    "00001111", -- 7871 - 0x1ebf  :   15 - 0xf
    "00000000", -- 7872 - 0x1ec0  :    0 - 0x0 -- Background 0xec
    "00000000", -- 7873 - 0x1ec1  :    0 - 0x0
    "00000000", -- 7874 - 0x1ec2  :    0 - 0x0
    "00000000", -- 7875 - 0x1ec3  :    0 - 0x0
    "00000000", -- 7876 - 0x1ec4  :    0 - 0x0
    "00000000", -- 7877 - 0x1ec5  :    0 - 0x0
    "00000000", -- 7878 - 0x1ec6  :    0 - 0x0
    "00000000", -- 7879 - 0x1ec7  :    0 - 0x0
    "00000000", -- 7880 - 0x1ec8  :    0 - 0x0
    "00000000", -- 7881 - 0x1ec9  :    0 - 0x0
    "00000000", -- 7882 - 0x1eca  :    0 - 0x0
    "00000000", -- 7883 - 0x1ecb  :    0 - 0x0
    "00000000", -- 7884 - 0x1ecc  :    0 - 0x0
    "00000000", -- 7885 - 0x1ecd  :    0 - 0x0
    "00000000", -- 7886 - 0x1ece  :    0 - 0x0
    "00000000", -- 7887 - 0x1ecf  :    0 - 0x0
    "00000000", -- 7888 - 0x1ed0  :    0 - 0x0 -- Background 0xed
    "00000000", -- 7889 - 0x1ed1  :    0 - 0x0
    "00000000", -- 7890 - 0x1ed2  :    0 - 0x0
    "00000000", -- 7891 - 0x1ed3  :    0 - 0x0
    "00000000", -- 7892 - 0x1ed4  :    0 - 0x0
    "00000000", -- 7893 - 0x1ed5  :    0 - 0x0
    "00000000", -- 7894 - 0x1ed6  :    0 - 0x0
    "00000000", -- 7895 - 0x1ed7  :    0 - 0x0
    "00000000", -- 7896 - 0x1ed8  :    0 - 0x0
    "00000000", -- 7897 - 0x1ed9  :    0 - 0x0
    "00000000", -- 7898 - 0x1eda  :    0 - 0x0
    "00000000", -- 7899 - 0x1edb  :    0 - 0x0
    "00000000", -- 7900 - 0x1edc  :    0 - 0x0
    "00000000", -- 7901 - 0x1edd  :    0 - 0x0
    "00000000", -- 7902 - 0x1ede  :    0 - 0x0
    "00000000", -- 7903 - 0x1edf  :    0 - 0x0
    "00000000", -- 7904 - 0x1ee0  :    0 - 0x0 -- Background 0xee
    "00000000", -- 7905 - 0x1ee1  :    0 - 0x0
    "00000000", -- 7906 - 0x1ee2  :    0 - 0x0
    "00000000", -- 7907 - 0x1ee3  :    0 - 0x0
    "00000000", -- 7908 - 0x1ee4  :    0 - 0x0
    "00000000", -- 7909 - 0x1ee5  :    0 - 0x0
    "00000000", -- 7910 - 0x1ee6  :    0 - 0x0
    "00000000", -- 7911 - 0x1ee7  :    0 - 0x0
    "00000000", -- 7912 - 0x1ee8  :    0 - 0x0
    "00000000", -- 7913 - 0x1ee9  :    0 - 0x0
    "00000000", -- 7914 - 0x1eea  :    0 - 0x0
    "00000000", -- 7915 - 0x1eeb  :    0 - 0x0
    "00000000", -- 7916 - 0x1eec  :    0 - 0x0
    "00000000", -- 7917 - 0x1eed  :    0 - 0x0
    "00000000", -- 7918 - 0x1eee  :    0 - 0x0
    "00000000", -- 7919 - 0x1eef  :    0 - 0x0
    "00000000", -- 7920 - 0x1ef0  :    0 - 0x0 -- Background 0xef
    "00000000", -- 7921 - 0x1ef1  :    0 - 0x0
    "00000000", -- 7922 - 0x1ef2  :    0 - 0x0
    "00000000", -- 7923 - 0x1ef3  :    0 - 0x0
    "00000000", -- 7924 - 0x1ef4  :    0 - 0x0
    "00000000", -- 7925 - 0x1ef5  :    0 - 0x0
    "00000000", -- 7926 - 0x1ef6  :    0 - 0x0
    "00000000", -- 7927 - 0x1ef7  :    0 - 0x0
    "00000000", -- 7928 - 0x1ef8  :    0 - 0x0
    "00000000", -- 7929 - 0x1ef9  :    0 - 0x0
    "00000000", -- 7930 - 0x1efa  :    0 - 0x0
    "00000000", -- 7931 - 0x1efb  :    0 - 0x0
    "00000000", -- 7932 - 0x1efc  :    0 - 0x0
    "00000000", -- 7933 - 0x1efd  :    0 - 0x0
    "00000000", -- 7934 - 0x1efe  :    0 - 0x0
    "00000000", -- 7935 - 0x1eff  :    0 - 0x0
    "11111111", -- 7936 - 0x1f00  :  255 - 0xff -- Background 0xf0
    "11111111", -- 7937 - 0x1f01  :  255 - 0xff
    "11111111", -- 7938 - 0x1f02  :  255 - 0xff
    "11111111", -- 7939 - 0x1f03  :  255 - 0xff
    "11111111", -- 7940 - 0x1f04  :  255 - 0xff
    "11111111", -- 7941 - 0x1f05  :  255 - 0xff
    "11111111", -- 7942 - 0x1f06  :  255 - 0xff
    "11111111", -- 7943 - 0x1f07  :  255 - 0xff
    "11111111", -- 7944 - 0x1f08  :  255 - 0xff
    "11111111", -- 7945 - 0x1f09  :  255 - 0xff
    "11111111", -- 7946 - 0x1f0a  :  255 - 0xff
    "11111111", -- 7947 - 0x1f0b  :  255 - 0xff
    "11111111", -- 7948 - 0x1f0c  :  255 - 0xff
    "11111111", -- 7949 - 0x1f0d  :  255 - 0xff
    "11111111", -- 7950 - 0x1f0e  :  255 - 0xff
    "11111111", -- 7951 - 0x1f0f  :  255 - 0xff
    "11111111", -- 7952 - 0x1f10  :  255 - 0xff -- Background 0xf1
    "11111111", -- 7953 - 0x1f11  :  255 - 0xff
    "11111111", -- 7954 - 0x1f12  :  255 - 0xff
    "11111111", -- 7955 - 0x1f13  :  255 - 0xff
    "11111111", -- 7956 - 0x1f14  :  255 - 0xff
    "11111111", -- 7957 - 0x1f15  :  255 - 0xff
    "11111111", -- 7958 - 0x1f16  :  255 - 0xff
    "11111111", -- 7959 - 0x1f17  :  255 - 0xff
    "11111111", -- 7960 - 0x1f18  :  255 - 0xff
    "11111111", -- 7961 - 0x1f19  :  255 - 0xff
    "11111111", -- 7962 - 0x1f1a  :  255 - 0xff
    "11111111", -- 7963 - 0x1f1b  :  255 - 0xff
    "11111111", -- 7964 - 0x1f1c  :  255 - 0xff
    "11111111", -- 7965 - 0x1f1d  :  255 - 0xff
    "11111111", -- 7966 - 0x1f1e  :  255 - 0xff
    "11111111", -- 7967 - 0x1f1f  :  255 - 0xff
    "11111111", -- 7968 - 0x1f20  :  255 - 0xff -- Background 0xf2
    "11111111", -- 7969 - 0x1f21  :  255 - 0xff
    "11111111", -- 7970 - 0x1f22  :  255 - 0xff
    "11111111", -- 7971 - 0x1f23  :  255 - 0xff
    "11111111", -- 7972 - 0x1f24  :  255 - 0xff
    "11111111", -- 7973 - 0x1f25  :  255 - 0xff
    "11111111", -- 7974 - 0x1f26  :  255 - 0xff
    "11111111", -- 7975 - 0x1f27  :  255 - 0xff
    "11111111", -- 7976 - 0x1f28  :  255 - 0xff
    "11111111", -- 7977 - 0x1f29  :  255 - 0xff
    "11111111", -- 7978 - 0x1f2a  :  255 - 0xff
    "11111111", -- 7979 - 0x1f2b  :  255 - 0xff
    "11111111", -- 7980 - 0x1f2c  :  255 - 0xff
    "11111111", -- 7981 - 0x1f2d  :  255 - 0xff
    "11111111", -- 7982 - 0x1f2e  :  255 - 0xff
    "11111111", -- 7983 - 0x1f2f  :  255 - 0xff
    "11111111", -- 7984 - 0x1f30  :  255 - 0xff -- Background 0xf3
    "11111111", -- 7985 - 0x1f31  :  255 - 0xff
    "11111111", -- 7986 - 0x1f32  :  255 - 0xff
    "11111111", -- 7987 - 0x1f33  :  255 - 0xff
    "11111111", -- 7988 - 0x1f34  :  255 - 0xff
    "11111111", -- 7989 - 0x1f35  :  255 - 0xff
    "11111111", -- 7990 - 0x1f36  :  255 - 0xff
    "11111111", -- 7991 - 0x1f37  :  255 - 0xff
    "11111111", -- 7992 - 0x1f38  :  255 - 0xff
    "11111111", -- 7993 - 0x1f39  :  255 - 0xff
    "11111111", -- 7994 - 0x1f3a  :  255 - 0xff
    "11111111", -- 7995 - 0x1f3b  :  255 - 0xff
    "11111111", -- 7996 - 0x1f3c  :  255 - 0xff
    "11111111", -- 7997 - 0x1f3d  :  255 - 0xff
    "11111111", -- 7998 - 0x1f3e  :  255 - 0xff
    "11111111", -- 7999 - 0x1f3f  :  255 - 0xff
    "11111111", -- 8000 - 0x1f40  :  255 - 0xff -- Background 0xf4
    "11111111", -- 8001 - 0x1f41  :  255 - 0xff
    "11111111", -- 8002 - 0x1f42  :  255 - 0xff
    "11111111", -- 8003 - 0x1f43  :  255 - 0xff
    "11111111", -- 8004 - 0x1f44  :  255 - 0xff
    "11111111", -- 8005 - 0x1f45  :  255 - 0xff
    "11111111", -- 8006 - 0x1f46  :  255 - 0xff
    "11111111", -- 8007 - 0x1f47  :  255 - 0xff
    "11111111", -- 8008 - 0x1f48  :  255 - 0xff
    "11111111", -- 8009 - 0x1f49  :  255 - 0xff
    "11111111", -- 8010 - 0x1f4a  :  255 - 0xff
    "11111111", -- 8011 - 0x1f4b  :  255 - 0xff
    "11111111", -- 8012 - 0x1f4c  :  255 - 0xff
    "11111111", -- 8013 - 0x1f4d  :  255 - 0xff
    "11111111", -- 8014 - 0x1f4e  :  255 - 0xff
    "11111111", -- 8015 - 0x1f4f  :  255 - 0xff
    "11111111", -- 8016 - 0x1f50  :  255 - 0xff -- Background 0xf5
    "11111111", -- 8017 - 0x1f51  :  255 - 0xff
    "11111111", -- 8018 - 0x1f52  :  255 - 0xff
    "11111111", -- 8019 - 0x1f53  :  255 - 0xff
    "11111111", -- 8020 - 0x1f54  :  255 - 0xff
    "11111111", -- 8021 - 0x1f55  :  255 - 0xff
    "11111111", -- 8022 - 0x1f56  :  255 - 0xff
    "11111111", -- 8023 - 0x1f57  :  255 - 0xff
    "11111111", -- 8024 - 0x1f58  :  255 - 0xff
    "11111111", -- 8025 - 0x1f59  :  255 - 0xff
    "11111111", -- 8026 - 0x1f5a  :  255 - 0xff
    "11111111", -- 8027 - 0x1f5b  :  255 - 0xff
    "11111111", -- 8028 - 0x1f5c  :  255 - 0xff
    "11111111", -- 8029 - 0x1f5d  :  255 - 0xff
    "11111111", -- 8030 - 0x1f5e  :  255 - 0xff
    "11111111", -- 8031 - 0x1f5f  :  255 - 0xff
    "11111111", -- 8032 - 0x1f60  :  255 - 0xff -- Background 0xf6
    "11111111", -- 8033 - 0x1f61  :  255 - 0xff
    "11111111", -- 8034 - 0x1f62  :  255 - 0xff
    "11111111", -- 8035 - 0x1f63  :  255 - 0xff
    "11111111", -- 8036 - 0x1f64  :  255 - 0xff
    "11111111", -- 8037 - 0x1f65  :  255 - 0xff
    "11111111", -- 8038 - 0x1f66  :  255 - 0xff
    "11111111", -- 8039 - 0x1f67  :  255 - 0xff
    "11111111", -- 8040 - 0x1f68  :  255 - 0xff
    "11111111", -- 8041 - 0x1f69  :  255 - 0xff
    "11111111", -- 8042 - 0x1f6a  :  255 - 0xff
    "11111111", -- 8043 - 0x1f6b  :  255 - 0xff
    "11111111", -- 8044 - 0x1f6c  :  255 - 0xff
    "11111111", -- 8045 - 0x1f6d  :  255 - 0xff
    "11111111", -- 8046 - 0x1f6e  :  255 - 0xff
    "11111111", -- 8047 - 0x1f6f  :  255 - 0xff
    "11111111", -- 8048 - 0x1f70  :  255 - 0xff -- Background 0xf7
    "11111111", -- 8049 - 0x1f71  :  255 - 0xff
    "11111111", -- 8050 - 0x1f72  :  255 - 0xff
    "11111111", -- 8051 - 0x1f73  :  255 - 0xff
    "11111111", -- 8052 - 0x1f74  :  255 - 0xff
    "11111111", -- 8053 - 0x1f75  :  255 - 0xff
    "11111111", -- 8054 - 0x1f76  :  255 - 0xff
    "11111111", -- 8055 - 0x1f77  :  255 - 0xff
    "11111111", -- 8056 - 0x1f78  :  255 - 0xff
    "11111111", -- 8057 - 0x1f79  :  255 - 0xff
    "11111111", -- 8058 - 0x1f7a  :  255 - 0xff
    "11111111", -- 8059 - 0x1f7b  :  255 - 0xff
    "11111111", -- 8060 - 0x1f7c  :  255 - 0xff
    "11111111", -- 8061 - 0x1f7d  :  255 - 0xff
    "11111111", -- 8062 - 0x1f7e  :  255 - 0xff
    "11111111", -- 8063 - 0x1f7f  :  255 - 0xff
    "11111111", -- 8064 - 0x1f80  :  255 - 0xff -- Background 0xf8
    "11111111", -- 8065 - 0x1f81  :  255 - 0xff
    "11111111", -- 8066 - 0x1f82  :  255 - 0xff
    "11111111", -- 8067 - 0x1f83  :  255 - 0xff
    "11111111", -- 8068 - 0x1f84  :  255 - 0xff
    "11111111", -- 8069 - 0x1f85  :  255 - 0xff
    "11111111", -- 8070 - 0x1f86  :  255 - 0xff
    "11111111", -- 8071 - 0x1f87  :  255 - 0xff
    "11111111", -- 8072 - 0x1f88  :  255 - 0xff
    "11111111", -- 8073 - 0x1f89  :  255 - 0xff
    "11111111", -- 8074 - 0x1f8a  :  255 - 0xff
    "11111111", -- 8075 - 0x1f8b  :  255 - 0xff
    "11111111", -- 8076 - 0x1f8c  :  255 - 0xff
    "11111111", -- 8077 - 0x1f8d  :  255 - 0xff
    "11111111", -- 8078 - 0x1f8e  :  255 - 0xff
    "11111111", -- 8079 - 0x1f8f  :  255 - 0xff
    "11111111", -- 8080 - 0x1f90  :  255 - 0xff -- Background 0xf9
    "11111111", -- 8081 - 0x1f91  :  255 - 0xff
    "11111111", -- 8082 - 0x1f92  :  255 - 0xff
    "11111111", -- 8083 - 0x1f93  :  255 - 0xff
    "11111111", -- 8084 - 0x1f94  :  255 - 0xff
    "11111111", -- 8085 - 0x1f95  :  255 - 0xff
    "11111111", -- 8086 - 0x1f96  :  255 - 0xff
    "11111111", -- 8087 - 0x1f97  :  255 - 0xff
    "11111111", -- 8088 - 0x1f98  :  255 - 0xff
    "11111111", -- 8089 - 0x1f99  :  255 - 0xff
    "11111111", -- 8090 - 0x1f9a  :  255 - 0xff
    "11111111", -- 8091 - 0x1f9b  :  255 - 0xff
    "11111111", -- 8092 - 0x1f9c  :  255 - 0xff
    "11111111", -- 8093 - 0x1f9d  :  255 - 0xff
    "11111111", -- 8094 - 0x1f9e  :  255 - 0xff
    "11111111", -- 8095 - 0x1f9f  :  255 - 0xff
    "11111111", -- 8096 - 0x1fa0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 8097 - 0x1fa1  :  255 - 0xff
    "11111111", -- 8098 - 0x1fa2  :  255 - 0xff
    "11111111", -- 8099 - 0x1fa3  :  255 - 0xff
    "11111111", -- 8100 - 0x1fa4  :  255 - 0xff
    "11111111", -- 8101 - 0x1fa5  :  255 - 0xff
    "11111111", -- 8102 - 0x1fa6  :  255 - 0xff
    "11111111", -- 8103 - 0x1fa7  :  255 - 0xff
    "11111111", -- 8104 - 0x1fa8  :  255 - 0xff
    "11111111", -- 8105 - 0x1fa9  :  255 - 0xff
    "11111111", -- 8106 - 0x1faa  :  255 - 0xff
    "11111111", -- 8107 - 0x1fab  :  255 - 0xff
    "11111111", -- 8108 - 0x1fac  :  255 - 0xff
    "11111111", -- 8109 - 0x1fad  :  255 - 0xff
    "11111111", -- 8110 - 0x1fae  :  255 - 0xff
    "11111111", -- 8111 - 0x1faf  :  255 - 0xff
    "11111111", -- 8112 - 0x1fb0  :  255 - 0xff -- Background 0xfb
    "11111111", -- 8113 - 0x1fb1  :  255 - 0xff
    "11111111", -- 8114 - 0x1fb2  :  255 - 0xff
    "11111111", -- 8115 - 0x1fb3  :  255 - 0xff
    "11111111", -- 8116 - 0x1fb4  :  255 - 0xff
    "11111111", -- 8117 - 0x1fb5  :  255 - 0xff
    "11111111", -- 8118 - 0x1fb6  :  255 - 0xff
    "11111111", -- 8119 - 0x1fb7  :  255 - 0xff
    "11111111", -- 8120 - 0x1fb8  :  255 - 0xff
    "11111111", -- 8121 - 0x1fb9  :  255 - 0xff
    "11111111", -- 8122 - 0x1fba  :  255 - 0xff
    "11111111", -- 8123 - 0x1fbb  :  255 - 0xff
    "11111111", -- 8124 - 0x1fbc  :  255 - 0xff
    "11111111", -- 8125 - 0x1fbd  :  255 - 0xff
    "11111111", -- 8126 - 0x1fbe  :  255 - 0xff
    "11111111", -- 8127 - 0x1fbf  :  255 - 0xff
    "11111111", -- 8128 - 0x1fc0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 8129 - 0x1fc1  :  255 - 0xff
    "11111111", -- 8130 - 0x1fc2  :  255 - 0xff
    "11111111", -- 8131 - 0x1fc3  :  255 - 0xff
    "11111111", -- 8132 - 0x1fc4  :  255 - 0xff
    "11111111", -- 8133 - 0x1fc5  :  255 - 0xff
    "11111111", -- 8134 - 0x1fc6  :  255 - 0xff
    "11111111", -- 8135 - 0x1fc7  :  255 - 0xff
    "11111111", -- 8136 - 0x1fc8  :  255 - 0xff
    "11111111", -- 8137 - 0x1fc9  :  255 - 0xff
    "11111111", -- 8138 - 0x1fca  :  255 - 0xff
    "11111111", -- 8139 - 0x1fcb  :  255 - 0xff
    "11111111", -- 8140 - 0x1fcc  :  255 - 0xff
    "11111111", -- 8141 - 0x1fcd  :  255 - 0xff
    "11111111", -- 8142 - 0x1fce  :  255 - 0xff
    "11111111", -- 8143 - 0x1fcf  :  255 - 0xff
    "11111111", -- 8144 - 0x1fd0  :  255 - 0xff -- Background 0xfd
    "11111111", -- 8145 - 0x1fd1  :  255 - 0xff
    "11111111", -- 8146 - 0x1fd2  :  255 - 0xff
    "11111111", -- 8147 - 0x1fd3  :  255 - 0xff
    "11111111", -- 8148 - 0x1fd4  :  255 - 0xff
    "11111111", -- 8149 - 0x1fd5  :  255 - 0xff
    "11111111", -- 8150 - 0x1fd6  :  255 - 0xff
    "11111111", -- 8151 - 0x1fd7  :  255 - 0xff
    "11111111", -- 8152 - 0x1fd8  :  255 - 0xff
    "11111111", -- 8153 - 0x1fd9  :  255 - 0xff
    "11111111", -- 8154 - 0x1fda  :  255 - 0xff
    "11111111", -- 8155 - 0x1fdb  :  255 - 0xff
    "11111111", -- 8156 - 0x1fdc  :  255 - 0xff
    "11111111", -- 8157 - 0x1fdd  :  255 - 0xff
    "11111111", -- 8158 - 0x1fde  :  255 - 0xff
    "11111111", -- 8159 - 0x1fdf  :  255 - 0xff
    "11111111", -- 8160 - 0x1fe0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 8161 - 0x1fe1  :  255 - 0xff
    "11111111", -- 8162 - 0x1fe2  :  255 - 0xff
    "11111111", -- 8163 - 0x1fe3  :  255 - 0xff
    "11111111", -- 8164 - 0x1fe4  :  255 - 0xff
    "11111111", -- 8165 - 0x1fe5  :  255 - 0xff
    "11111111", -- 8166 - 0x1fe6  :  255 - 0xff
    "11111111", -- 8167 - 0x1fe7  :  255 - 0xff
    "11111111", -- 8168 - 0x1fe8  :  255 - 0xff
    "11111111", -- 8169 - 0x1fe9  :  255 - 0xff
    "11111111", -- 8170 - 0x1fea  :  255 - 0xff
    "11111111", -- 8171 - 0x1feb  :  255 - 0xff
    "11111111", -- 8172 - 0x1fec  :  255 - 0xff
    "11111111", -- 8173 - 0x1fed  :  255 - 0xff
    "11111111", -- 8174 - 0x1fee  :  255 - 0xff
    "11111111", -- 8175 - 0x1fef  :  255 - 0xff
    "11111111", -- 8176 - 0x1ff0  :  255 - 0xff -- Background 0xff
    "11111111", -- 8177 - 0x1ff1  :  255 - 0xff
    "11111111", -- 8178 - 0x1ff2  :  255 - 0xff
    "11111111", -- 8179 - 0x1ff3  :  255 - 0xff
    "11111111", -- 8180 - 0x1ff4  :  255 - 0xff
    "11111111", -- 8181 - 0x1ff5  :  255 - 0xff
    "11111111", -- 8182 - 0x1ff6  :  255 - 0xff
    "11111111", -- 8183 - 0x1ff7  :  255 - 0xff
    "11111111", -- 8184 - 0x1ff8  :  255 - 0xff
    "11111111", -- 8185 - 0x1ff9  :  255 - 0xff
    "11111111", -- 8186 - 0x1ffa  :  255 - 0xff
    "11111111", -- 8187 - 0x1ffb  :  255 - 0xff
    "11111111", -- 8188 - 0x1ffc  :  255 - 0xff
    "11111111", -- 8189 - 0x1ffd  :  255 - 0xff
    "11111111", -- 8190 - 0x1ffe  :  255 - 0xff
    "11111111"  -- 8191 - 0x1fff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
