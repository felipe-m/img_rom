--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: pacman_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_PACMAN_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_PACMAN_00;

architecture BEHAVIORAL of ROM_NTABLE_PACMAN_00 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00100000", --    0 -  0x0  :   32 - 0x20 -- line 0x0
    "00100000", --    1 -  0x1  :   32 - 0x20
    "00100000", --    2 -  0x2  :   32 - 0x20
    "00100000", --    3 -  0x3  :   32 - 0x20
    "00100000", --    4 -  0x4  :   32 - 0x20
    "00100000", --    5 -  0x5  :   32 - 0x20
    "00100000", --    6 -  0x6  :   32 - 0x20
    "00100000", --    7 -  0x7  :   32 - 0x20
    "00100000", --    8 -  0x8  :   32 - 0x20
    "00100000", --    9 -  0x9  :   32 - 0x20
    "00100000", --   10 -  0xa  :   32 - 0x20
    "00100000", --   11 -  0xb  :   32 - 0x20
    "00100000", --   12 -  0xc  :   32 - 0x20
    "00100000", --   13 -  0xd  :   32 - 0x20
    "00100000", --   14 -  0xe  :   32 - 0x20
    "00100000", --   15 -  0xf  :   32 - 0x20
    "00100000", --   16 - 0x10  :   32 - 0x20
    "00100000", --   17 - 0x11  :   32 - 0x20
    "00100000", --   18 - 0x12  :   32 - 0x20
    "00100000", --   19 - 0x13  :   32 - 0x20
    "00100000", --   20 - 0x14  :   32 - 0x20
    "00100000", --   21 - 0x15  :   32 - 0x20
    "00100000", --   22 - 0x16  :   32 - 0x20
    "00100000", --   23 - 0x17  :   32 - 0x20
    "00100000", --   24 - 0x18  :   32 - 0x20
    "00100000", --   25 - 0x19  :   32 - 0x20
    "00100000", --   26 - 0x1a  :   32 - 0x20
    "00100000", --   27 - 0x1b  :   32 - 0x20
    "00100000", --   28 - 0x1c  :   32 - 0x20
    "00100000", --   29 - 0x1d  :   32 - 0x20
    "00100000", --   30 - 0x1e  :   32 - 0x20
    "00100000", --   31 - 0x1f  :   32 - 0x20
    "00100000", --   32 - 0x20  :   32 - 0x20 -- line 0x1
    "00100000", --   33 - 0x21  :   32 - 0x20
    "00100000", --   34 - 0x22  :   32 - 0x20
    "00100000", --   35 - 0x23  :   32 - 0x20
    "00100000", --   36 - 0x24  :   32 - 0x20
    "00100000", --   37 - 0x25  :   32 - 0x20
    "00100000", --   38 - 0x26  :   32 - 0x20
    "00100000", --   39 - 0x27  :   32 - 0x20
    "00100000", --   40 - 0x28  :   32 - 0x20
    "00100000", --   41 - 0x29  :   32 - 0x20
    "00100000", --   42 - 0x2a  :   32 - 0x20
    "00100000", --   43 - 0x2b  :   32 - 0x20
    "00100000", --   44 - 0x2c  :   32 - 0x20
    "00100000", --   45 - 0x2d  :   32 - 0x20
    "00100000", --   46 - 0x2e  :   32 - 0x20
    "00100000", --   47 - 0x2f  :   32 - 0x20
    "00100000", --   48 - 0x30  :   32 - 0x20
    "00100000", --   49 - 0x31  :   32 - 0x20
    "00100000", --   50 - 0x32  :   32 - 0x20
    "00100000", --   51 - 0x33  :   32 - 0x20
    "00100000", --   52 - 0x34  :   32 - 0x20
    "00100000", --   53 - 0x35  :   32 - 0x20
    "00100000", --   54 - 0x36  :   32 - 0x20
    "00100000", --   55 - 0x37  :   32 - 0x20
    "00100000", --   56 - 0x38  :   32 - 0x20
    "00100000", --   57 - 0x39  :   32 - 0x20
    "00100000", --   58 - 0x3a  :   32 - 0x20
    "00100000", --   59 - 0x3b  :   32 - 0x20
    "00100000", --   60 - 0x3c  :   32 - 0x20
    "00100000", --   61 - 0x3d  :   32 - 0x20
    "00100000", --   62 - 0x3e  :   32 - 0x20
    "00100000", --   63 - 0x3f  :   32 - 0x20
    "00101101", --   64 - 0x40  :   45 - 0x2d -- line 0x2
    "00011111", --   65 - 0x41  :   31 - 0x1f
    "00010000", --   66 - 0x42  :   16 - 0x10
    "00010000", --   67 - 0x43  :   16 - 0x10
    "00010000", --   68 - 0x44  :   16 - 0x10
    "00010000", --   69 - 0x45  :   16 - 0x10
    "00010000", --   70 - 0x46  :   16 - 0x10
    "00010000", --   71 - 0x47  :   16 - 0x10
    "00010000", --   72 - 0x48  :   16 - 0x10
    "00010000", --   73 - 0x49  :   16 - 0x10
    "00010000", --   74 - 0x4a  :   16 - 0x10
    "00010011", --   75 - 0x4b  :   19 - 0x13
    "00010000", --   76 - 0x4c  :   16 - 0x10
    "00010000", --   77 - 0x4d  :   16 - 0x10
    "00010000", --   78 - 0x4e  :   16 - 0x10
    "00010000", --   79 - 0x4f  :   16 - 0x10
    "00010000", --   80 - 0x50  :   16 - 0x10
    "00010000", --   81 - 0x51  :   16 - 0x10
    "00010000", --   82 - 0x52  :   16 - 0x10
    "00010000", --   83 - 0x53  :   16 - 0x10
    "00010000", --   84 - 0x54  :   16 - 0x10
    "00011101", --   85 - 0x55  :   29 - 0x1d
    "00100000", --   86 - 0x56  :   32 - 0x20
    "00100000", --   87 - 0x57  :   32 - 0x20
    "00100000", --   88 - 0x58  :   32 - 0x20
    "00100000", --   89 - 0x59  :   32 - 0x20
    "00100000", --   90 - 0x5a  :   32 - 0x20
    "00100000", --   91 - 0x5b  :   32 - 0x20
    "00100000", --   92 - 0x5c  :   32 - 0x20
    "00100000", --   93 - 0x5d  :   32 - 0x20
    "00100000", --   94 - 0x5e  :   32 - 0x20
    "00100000", --   95 - 0x5f  :   32 - 0x20
    "00101101", --   96 - 0x60  :   45 - 0x2d -- line 0x3
    "00010001", --   97 - 0x61  :   17 - 0x11
    "00000011", --   98 - 0x62  :    3 - 0x3
    "00000011", --   99 - 0x63  :    3 - 0x3
    "00000011", --  100 - 0x64  :    3 - 0x3
    "00000011", --  101 - 0x65  :    3 - 0x3
    "00000011", --  102 - 0x66  :    3 - 0x3
    "00000011", --  103 - 0x67  :    3 - 0x3
    "00000011", --  104 - 0x68  :    3 - 0x3
    "00000011", --  105 - 0x69  :    3 - 0x3
    "00000011", --  106 - 0x6a  :    3 - 0x3
    "00010001", --  107 - 0x6b  :   17 - 0x11
    "00000011", --  108 - 0x6c  :    3 - 0x3
    "00000011", --  109 - 0x6d  :    3 - 0x3
    "00000011", --  110 - 0x6e  :    3 - 0x3
    "00000011", --  111 - 0x6f  :    3 - 0x3
    "00000011", --  112 - 0x70  :    3 - 0x3
    "00000011", --  113 - 0x71  :    3 - 0x3
    "00000011", --  114 - 0x72  :    3 - 0x3
    "00000011", --  115 - 0x73  :    3 - 0x3
    "00000011", --  116 - 0x74  :    3 - 0x3
    "00010001", --  117 - 0x75  :   17 - 0x11
    "10110100", --  118 - 0x76  :  180 - 0xb4
    "10110101", --  119 - 0x77  :  181 - 0xb5
    "10110110", --  120 - 0x78  :  182 - 0xb6
    "10110111", --  121 - 0x79  :  183 - 0xb7
    "10111000", --  122 - 0x7a  :  184 - 0xb8
    "10111001", --  123 - 0x7b  :  185 - 0xb9
    "10111010", --  124 - 0x7c  :  186 - 0xba
    "10111011", --  125 - 0x7d  :  187 - 0xbb
    "00100000", --  126 - 0x7e  :   32 - 0x20
    "00100000", --  127 - 0x7f  :   32 - 0x20
    "00101101", --  128 - 0x80  :   45 - 0x2d -- line 0x4
    "00010001", --  129 - 0x81  :   17 - 0x11
    "00000011", --  130 - 0x82  :    3 - 0x3
    "00011111", --  131 - 0x83  :   31 - 0x1f
    "00010000", --  132 - 0x84  :   16 - 0x10
    "00011101", --  133 - 0x85  :   29 - 0x1d
    "00000011", --  134 - 0x86  :    3 - 0x3
    "00011111", --  135 - 0x87  :   31 - 0x1f
    "00010000", --  136 - 0x88  :   16 - 0x10
    "00011101", --  137 - 0x89  :   29 - 0x1d
    "00000011", --  138 - 0x8a  :    3 - 0x3
    "00010001", --  139 - 0x8b  :   17 - 0x11
    "00000011", --  140 - 0x8c  :    3 - 0x3
    "00011111", --  141 - 0x8d  :   31 - 0x1f
    "00010000", --  142 - 0x8e  :   16 - 0x10
    "00011101", --  143 - 0x8f  :   29 - 0x1d
    "00000011", --  144 - 0x90  :    3 - 0x3
    "00011111", --  145 - 0x91  :   31 - 0x1f
    "00010000", --  146 - 0x92  :   16 - 0x10
    "00011101", --  147 - 0x93  :   29 - 0x1d
    "00000011", --  148 - 0x94  :    3 - 0x3
    "00010001", --  149 - 0x95  :   17 - 0x11
    "00100000", --  150 - 0x96  :   32 - 0x20
    "00100000", --  151 - 0x97  :   32 - 0x20
    "00100000", --  152 - 0x98  :   32 - 0x20
    "00100000", --  153 - 0x99  :   32 - 0x20
    "00100000", --  154 - 0x9a  :   32 - 0x20
    "00100000", --  155 - 0x9b  :   32 - 0x20
    "00100000", --  156 - 0x9c  :   32 - 0x20
    "00100000", --  157 - 0x9d  :   32 - 0x20
    "00100000", --  158 - 0x9e  :   32 - 0x20
    "00100000", --  159 - 0x9f  :   32 - 0x20
    "00101101", --  160 - 0xa0  :   45 - 0x2d -- line 0x5
    "00010001", --  161 - 0xa1  :   17 - 0x11
    "00000001", --  162 - 0xa2  :    1 - 0x1
    "00010001", --  163 - 0xa3  :   17 - 0x11
    "00100000", --  164 - 0xa4  :   32 - 0x20
    "00010001", --  165 - 0xa5  :   17 - 0x11
    "00000011", --  166 - 0xa6  :    3 - 0x3
    "00010001", --  167 - 0xa7  :   17 - 0x11
    "00100000", --  168 - 0xa8  :   32 - 0x20
    "00010001", --  169 - 0xa9  :   17 - 0x11
    "00000011", --  170 - 0xaa  :    3 - 0x3
    "00010001", --  171 - 0xab  :   17 - 0x11
    "00000011", --  172 - 0xac  :    3 - 0x3
    "00010001", --  173 - 0xad  :   17 - 0x11
    "00100000", --  174 - 0xae  :   32 - 0x20
    "00010001", --  175 - 0xaf  :   17 - 0x11
    "00000011", --  176 - 0xb0  :    3 - 0x3
    "00010001", --  177 - 0xb1  :   17 - 0x11
    "00100000", --  178 - 0xb2  :   32 - 0x20
    "00010001", --  179 - 0xb3  :   17 - 0x11
    "00000001", --  180 - 0xb4  :    1 - 0x1
    "00010001", --  181 - 0xb5  :   17 - 0x11
    "00100000", --  182 - 0xb6  :   32 - 0x20
    "00100000", --  183 - 0xb7  :   32 - 0x20
    "00110001", --  184 - 0xb8  :   49 - 0x31
    "00110000", --  185 - 0xb9  :   48 - 0x30
    "00110000", --  186 - 0xba  :   48 - 0x30
    "00110000", --  187 - 0xbb  :   48 - 0x30
    "00110000", --  188 - 0xbc  :   48 - 0x30
    "00100000", --  189 - 0xbd  :   32 - 0x20
    "00100000", --  190 - 0xbe  :   32 - 0x20
    "00100000", --  191 - 0xbf  :   32 - 0x20
    "00101101", --  192 - 0xc0  :   45 - 0x2d -- line 0x6
    "00010001", --  193 - 0xc1  :   17 - 0x11
    "00000011", --  194 - 0xc2  :    3 - 0x3
    "00011110", --  195 - 0xc3  :   30 - 0x1e
    "00010000", --  196 - 0xc4  :   16 - 0x10
    "00011100", --  197 - 0xc5  :   28 - 0x1c
    "00000011", --  198 - 0xc6  :    3 - 0x3
    "00011110", --  199 - 0xc7  :   30 - 0x1e
    "00010000", --  200 - 0xc8  :   16 - 0x10
    "00011100", --  201 - 0xc9  :   28 - 0x1c
    "00000011", --  202 - 0xca  :    3 - 0x3
    "00011010", --  203 - 0xcb  :   26 - 0x1a
    "00000011", --  204 - 0xcc  :    3 - 0x3
    "00011110", --  205 - 0xcd  :   30 - 0x1e
    "00010000", --  206 - 0xce  :   16 - 0x10
    "00011100", --  207 - 0xcf  :   28 - 0x1c
    "00000011", --  208 - 0xd0  :    3 - 0x3
    "00011110", --  209 - 0xd1  :   30 - 0x1e
    "00010000", --  210 - 0xd2  :   16 - 0x10
    "00011100", --  211 - 0xd3  :   28 - 0x1c
    "00000011", --  212 - 0xd4  :    3 - 0x3
    "00010001", --  213 - 0xd5  :   17 - 0x11
    "00100000", --  214 - 0xd6  :   32 - 0x20
    "00100000", --  215 - 0xd7  :   32 - 0x20
    "00100000", --  216 - 0xd8  :   32 - 0x20
    "00100000", --  217 - 0xd9  :   32 - 0x20
    "00100000", --  218 - 0xda  :   32 - 0x20
    "00100000", --  219 - 0xdb  :   32 - 0x20
    "00100000", --  220 - 0xdc  :   32 - 0x20
    "00100000", --  221 - 0xdd  :   32 - 0x20
    "00100000", --  222 - 0xde  :   32 - 0x20
    "00100000", --  223 - 0xdf  :   32 - 0x20
    "00101101", --  224 - 0xe0  :   45 - 0x2d -- line 0x7
    "00010001", --  225 - 0xe1  :   17 - 0x11
    "00000011", --  226 - 0xe2  :    3 - 0x3
    "00000011", --  227 - 0xe3  :    3 - 0x3
    "00000011", --  228 - 0xe4  :    3 - 0x3
    "00000011", --  229 - 0xe5  :    3 - 0x3
    "00000011", --  230 - 0xe6  :    3 - 0x3
    "00000011", --  231 - 0xe7  :    3 - 0x3
    "00000011", --  232 - 0xe8  :    3 - 0x3
    "00000011", --  233 - 0xe9  :    3 - 0x3
    "00000011", --  234 - 0xea  :    3 - 0x3
    "00000011", --  235 - 0xeb  :    3 - 0x3
    "00000011", --  236 - 0xec  :    3 - 0x3
    "00000011", --  237 - 0xed  :    3 - 0x3
    "00000011", --  238 - 0xee  :    3 - 0x3
    "00000011", --  239 - 0xef  :    3 - 0x3
    "00000011", --  240 - 0xf0  :    3 - 0x3
    "00000011", --  241 - 0xf1  :    3 - 0x3
    "00000011", --  242 - 0xf2  :    3 - 0x3
    "00000011", --  243 - 0xf3  :    3 - 0x3
    "00000011", --  244 - 0xf4  :    3 - 0x3
    "00010001", --  245 - 0xf5  :   17 - 0x11
    "00100000", --  246 - 0xf6  :   32 - 0x20
    "00100000", --  247 - 0xf7  :   32 - 0x20
    "00100000", --  248 - 0xf8  :   32 - 0x20
    "00100000", --  249 - 0xf9  :   32 - 0x20
    "00100000", --  250 - 0xfa  :   32 - 0x20
    "00100000", --  251 - 0xfb  :   32 - 0x20
    "00100000", --  252 - 0xfc  :   32 - 0x20
    "00100000", --  253 - 0xfd  :   32 - 0x20
    "00100000", --  254 - 0xfe  :   32 - 0x20
    "00100000", --  255 - 0xff  :   32 - 0x20
    "00101101", --  256 - 0x100  :   45 - 0x2d -- line 0x8
    "00010001", --  257 - 0x101  :   17 - 0x11
    "00000011", --  258 - 0x102  :    3 - 0x3
    "00011111", --  259 - 0x103  :   31 - 0x1f
    "00010000", --  260 - 0x104  :   16 - 0x10
    "00011101", --  261 - 0x105  :   29 - 0x1d
    "00000011", --  262 - 0x106  :    3 - 0x3
    "00011011", --  263 - 0x107  :   27 - 0x1b
    "00000011", --  264 - 0x108  :    3 - 0x3
    "00011111", --  265 - 0x109  :   31 - 0x1f
    "00010000", --  266 - 0x10a  :   16 - 0x10
    "00010000", --  267 - 0x10b  :   16 - 0x10
    "00010000", --  268 - 0x10c  :   16 - 0x10
    "00011101", --  269 - 0x10d  :   29 - 0x1d
    "00000011", --  270 - 0x10e  :    3 - 0x3
    "00011011", --  271 - 0x10f  :   27 - 0x1b
    "00000011", --  272 - 0x110  :    3 - 0x3
    "00011111", --  273 - 0x111  :   31 - 0x1f
    "00010000", --  274 - 0x112  :   16 - 0x10
    "00011101", --  275 - 0x113  :   29 - 0x1d
    "00000011", --  276 - 0x114  :    3 - 0x3
    "00010001", --  277 - 0x115  :   17 - 0x11
    "00100000", --  278 - 0x116  :   32 - 0x20
    "00100000", --  279 - 0x117  :   32 - 0x20
    "00100000", --  280 - 0x118  :   32 - 0x20
    "00100000", --  281 - 0x119  :   32 - 0x20
    "00100000", --  282 - 0x11a  :   32 - 0x20
    "00100000", --  283 - 0x11b  :   32 - 0x20
    "00100000", --  284 - 0x11c  :   32 - 0x20
    "00100000", --  285 - 0x11d  :   32 - 0x20
    "00100000", --  286 - 0x11e  :   32 - 0x20
    "00100000", --  287 - 0x11f  :   32 - 0x20
    "00101101", --  288 - 0x120  :   45 - 0x2d -- line 0x9
    "00010001", --  289 - 0x121  :   17 - 0x11
    "00000011", --  290 - 0x122  :    3 - 0x3
    "00011110", --  291 - 0x123  :   30 - 0x1e
    "00010000", --  292 - 0x124  :   16 - 0x10
    "00011100", --  293 - 0x125  :   28 - 0x1c
    "00000011", --  294 - 0x126  :    3 - 0x3
    "00010001", --  295 - 0x127  :   17 - 0x11
    "00000011", --  296 - 0x128  :    3 - 0x3
    "00011110", --  297 - 0x129  :   30 - 0x1e
    "00010000", --  298 - 0x12a  :   16 - 0x10
    "00010011", --  299 - 0x12b  :   19 - 0x13
    "00010000", --  300 - 0x12c  :   16 - 0x10
    "00011100", --  301 - 0x12d  :   28 - 0x1c
    "00000011", --  302 - 0x12e  :    3 - 0x3
    "00010001", --  303 - 0x12f  :   17 - 0x11
    "00000011", --  304 - 0x130  :    3 - 0x3
    "00011110", --  305 - 0x131  :   30 - 0x1e
    "00010000", --  306 - 0x132  :   16 - 0x10
    "00011100", --  307 - 0x133  :   28 - 0x1c
    "00000011", --  308 - 0x134  :    3 - 0x3
    "00010001", --  309 - 0x135  :   17 - 0x11
    "00100000", --  310 - 0x136  :   32 - 0x20
    "00100000", --  311 - 0x137  :   32 - 0x20
    "00100000", --  312 - 0x138  :   32 - 0x20
    "00100000", --  313 - 0x139  :   32 - 0x20
    "00100000", --  314 - 0x13a  :   32 - 0x20
    "00110000", --  315 - 0x13b  :   48 - 0x30
    "00110000", --  316 - 0x13c  :   48 - 0x30
    "00100000", --  317 - 0x13d  :   32 - 0x20
    "00100000", --  318 - 0x13e  :   32 - 0x20
    "00100000", --  319 - 0x13f  :   32 - 0x20
    "00101101", --  320 - 0x140  :   45 - 0x2d -- line 0xa
    "00010001", --  321 - 0x141  :   17 - 0x11
    "00000011", --  322 - 0x142  :    3 - 0x3
    "00000011", --  323 - 0x143  :    3 - 0x3
    "00000011", --  324 - 0x144  :    3 - 0x3
    "00000011", --  325 - 0x145  :    3 - 0x3
    "00000011", --  326 - 0x146  :    3 - 0x3
    "00010001", --  327 - 0x147  :   17 - 0x11
    "00000011", --  328 - 0x148  :    3 - 0x3
    "00000011", --  329 - 0x149  :    3 - 0x3
    "00000011", --  330 - 0x14a  :    3 - 0x3
    "00010001", --  331 - 0x14b  :   17 - 0x11
    "00000011", --  332 - 0x14c  :    3 - 0x3
    "00000011", --  333 - 0x14d  :    3 - 0x3
    "00000011", --  334 - 0x14e  :    3 - 0x3
    "00010001", --  335 - 0x14f  :   17 - 0x11
    "00000011", --  336 - 0x150  :    3 - 0x3
    "00000011", --  337 - 0x151  :    3 - 0x3
    "00000011", --  338 - 0x152  :    3 - 0x3
    "00000011", --  339 - 0x153  :    3 - 0x3
    "00000011", --  340 - 0x154  :    3 - 0x3
    "00010001", --  341 - 0x155  :   17 - 0x11
    "00100000", --  342 - 0x156  :   32 - 0x20
    "00100000", --  343 - 0x157  :   32 - 0x20
    "00100000", --  344 - 0x158  :   32 - 0x20
    "00100000", --  345 - 0x159  :   32 - 0x20
    "00100000", --  346 - 0x15a  :   32 - 0x20
    "00100000", --  347 - 0x15b  :   32 - 0x20
    "00100000", --  348 - 0x15c  :   32 - 0x20
    "00100000", --  349 - 0x15d  :   32 - 0x20
    "00100000", --  350 - 0x15e  :   32 - 0x20
    "00100000", --  351 - 0x15f  :   32 - 0x20
    "00101101", --  352 - 0x160  :   45 - 0x2d -- line 0xb
    "00011110", --  353 - 0x161  :   30 - 0x1e
    "00010000", --  354 - 0x162  :   16 - 0x10
    "00010000", --  355 - 0x163  :   16 - 0x10
    "00010000", --  356 - 0x164  :   16 - 0x10
    "00011101", --  357 - 0x165  :   29 - 0x1d
    "00000011", --  358 - 0x166  :    3 - 0x3
    "00010101", --  359 - 0x167  :   21 - 0x15
    "00010000", --  360 - 0x168  :   16 - 0x10
    "00011000", --  361 - 0x169  :   24 - 0x18
    "00001000", --  362 - 0x16a  :    8 - 0x8
    "00011010", --  363 - 0x16b  :   26 - 0x1a
    "00001000", --  364 - 0x16c  :    8 - 0x8
    "00011001", --  365 - 0x16d  :   25 - 0x19
    "00010000", --  366 - 0x16e  :   16 - 0x10
    "00010100", --  367 - 0x16f  :   20 - 0x14
    "00000011", --  368 - 0x170  :    3 - 0x3
    "00011111", --  369 - 0x171  :   31 - 0x1f
    "00010000", --  370 - 0x172  :   16 - 0x10
    "00010000", --  371 - 0x173  :   16 - 0x10
    "00010000", --  372 - 0x174  :   16 - 0x10
    "00011100", --  373 - 0x175  :   28 - 0x1c
    "00100000", --  374 - 0x176  :   32 - 0x20
    "00100000", --  375 - 0x177  :   32 - 0x20
    "00100000", --  376 - 0x178  :   32 - 0x20
    "00100000", --  377 - 0x179  :   32 - 0x20
    "00100000", --  378 - 0x17a  :   32 - 0x20
    "00100000", --  379 - 0x17b  :   32 - 0x20
    "00100000", --  380 - 0x17c  :   32 - 0x20
    "00100000", --  381 - 0x17d  :   32 - 0x20
    "00100000", --  382 - 0x17e  :   32 - 0x20
    "00100000", --  383 - 0x17f  :   32 - 0x20
    "00101101", --  384 - 0x180  :   45 - 0x2d -- line 0xc
    "00100000", --  385 - 0x181  :   32 - 0x20
    "00100000", --  386 - 0x182  :   32 - 0x20
    "00100000", --  387 - 0x183  :   32 - 0x20
    "00100000", --  388 - 0x184  :   32 - 0x20
    "00010001", --  389 - 0x185  :   17 - 0x11
    "00000011", --  390 - 0x186  :    3 - 0x3
    "00010001", --  391 - 0x187  :   17 - 0x11
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00010001", --  399 - 0x18f  :   17 - 0x11
    "00000011", --  400 - 0x190  :    3 - 0x3
    "00010001", --  401 - 0x191  :   17 - 0x11
    "00100000", --  402 - 0x192  :   32 - 0x20
    "00100000", --  403 - 0x193  :   32 - 0x20
    "00100000", --  404 - 0x194  :   32 - 0x20
    "00100000", --  405 - 0x195  :   32 - 0x20
    "00100000", --  406 - 0x196  :   32 - 0x20
    "00100000", --  407 - 0x197  :   32 - 0x20
    "00100000", --  408 - 0x198  :   32 - 0x20
    "00100000", --  409 - 0x199  :   32 - 0x20
    "00100000", --  410 - 0x19a  :   32 - 0x20
    "00100000", --  411 - 0x19b  :   32 - 0x20
    "00100000", --  412 - 0x19c  :   32 - 0x20
    "00100000", --  413 - 0x19d  :   32 - 0x20
    "00100000", --  414 - 0x19e  :   32 - 0x20
    "00100000", --  415 - 0x19f  :   32 - 0x20
    "00101101", --  416 - 0x1a0  :   45 - 0x2d -- line 0xd
    "00100000", --  417 - 0x1a1  :   32 - 0x20
    "00100000", --  418 - 0x1a2  :   32 - 0x20
    "00100000", --  419 - 0x1a3  :   32 - 0x20
    "00100000", --  420 - 0x1a4  :   32 - 0x20
    "00010001", --  421 - 0x1a5  :   17 - 0x11
    "00000011", --  422 - 0x1a6  :    3 - 0x3
    "00010001", --  423 - 0x1a7  :   17 - 0x11
    "00000000", --  424 - 0x1a8  :    0 - 0x0
    "00011111", --  425 - 0x1a9  :   31 - 0x1f
    "00010111", --  426 - 0x1aa  :   23 - 0x17
    "00101100", --  427 - 0x1ab  :   44 - 0x2c
    "00010110", --  428 - 0x1ac  :   22 - 0x16
    "00011101", --  429 - 0x1ad  :   29 - 0x1d
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00010001", --  431 - 0x1af  :   17 - 0x11
    "00000011", --  432 - 0x1b0  :    3 - 0x3
    "00010001", --  433 - 0x1b1  :   17 - 0x11
    "00100000", --  434 - 0x1b2  :   32 - 0x20
    "00100000", --  435 - 0x1b3  :   32 - 0x20
    "00100000", --  436 - 0x1b4  :   32 - 0x20
    "00100000", --  437 - 0x1b5  :   32 - 0x20
    "00100000", --  438 - 0x1b6  :   32 - 0x20
    "00100000", --  439 - 0x1b7  :   32 - 0x20
    "00100000", --  440 - 0x1b8  :   32 - 0x20
    "00100000", --  441 - 0x1b9  :   32 - 0x20
    "00100000", --  442 - 0x1ba  :   32 - 0x20
    "00100000", --  443 - 0x1bb  :   32 - 0x20
    "00100000", --  444 - 0x1bc  :   32 - 0x20
    "00100000", --  445 - 0x1bd  :   32 - 0x20
    "00100000", --  446 - 0x1be  :   32 - 0x20
    "00100000", --  447 - 0x1bf  :   32 - 0x20
    "00101101", --  448 - 0x1c0  :   45 - 0x2d -- line 0xe
    "00100010", --  449 - 0x1c1  :   34 - 0x22
    "00010000", --  450 - 0x1c2  :   16 - 0x10
    "00010000", --  451 - 0x1c3  :   16 - 0x10
    "00010000", --  452 - 0x1c4  :   16 - 0x10
    "00011100", --  453 - 0x1c5  :   28 - 0x1c
    "00000011", --  454 - 0x1c6  :    3 - 0x3
    "00011010", --  455 - 0x1c7  :   26 - 0x1a
    "00000000", --  456 - 0x1c8  :    0 - 0x0
    "00010001", --  457 - 0x1c9  :   17 - 0x11
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00010001", --  461 - 0x1cd  :   17 - 0x11
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00011010", --  463 - 0x1cf  :   26 - 0x1a
    "00000011", --  464 - 0x1d0  :    3 - 0x3
    "00011110", --  465 - 0x1d1  :   30 - 0x1e
    "00010000", --  466 - 0x1d2  :   16 - 0x10
    "00010000", --  467 - 0x1d3  :   16 - 0x10
    "00010000", --  468 - 0x1d4  :   16 - 0x10
    "00100001", --  469 - 0x1d5  :   33 - 0x21
    "00101101", --  470 - 0x1d6  :   45 - 0x2d
    "00101101", --  471 - 0x1d7  :   45 - 0x2d
    "00101101", --  472 - 0x1d8  :   45 - 0x2d
    "00101101", --  473 - 0x1d9  :   45 - 0x2d
    "00101101", --  474 - 0x1da  :   45 - 0x2d
    "00101101", --  475 - 0x1db  :   45 - 0x2d
    "00101101", --  476 - 0x1dc  :   45 - 0x2d
    "00101101", --  477 - 0x1dd  :   45 - 0x2d
    "00100000", --  478 - 0x1de  :   32 - 0x20
    "00100000", --  479 - 0x1df  :   32 - 0x20
    "00000100", --  480 - 0x1e0  :    4 - 0x4 -- line 0xf
    "00000110", --  481 - 0x1e1  :    6 - 0x6
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000011", --  486 - 0x1e6  :    3 - 0x3
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "00010001", --  489 - 0x1e9  :   17 - 0x11
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00010001", --  493 - 0x1ed  :   17 - 0x11
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000011", --  496 - 0x1f0  :    3 - 0x3
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000101", --  501 - 0x1f5  :    5 - 0x5
    "00000100", --  502 - 0x1f6  :    4 - 0x4
    "00000100", --  503 - 0x1f7  :    4 - 0x4
    "00000100", --  504 - 0x1f8  :    4 - 0x4
    "00000100", --  505 - 0x1f9  :    4 - 0x4
    "00000100", --  506 - 0x1fa  :    4 - 0x4
    "00000100", --  507 - 0x1fb  :    4 - 0x4
    "00000100", --  508 - 0x1fc  :    4 - 0x4
    "00000100", --  509 - 0x1fd  :    4 - 0x4
    "00100000", --  510 - 0x1fe  :   32 - 0x20
    "00100000", --  511 - 0x1ff  :   32 - 0x20
    "00101101", --  512 - 0x200  :   45 - 0x2d -- line 0x10
    "00100010", --  513 - 0x201  :   34 - 0x22
    "00010000", --  514 - 0x202  :   16 - 0x10
    "00010000", --  515 - 0x203  :   16 - 0x10
    "00010000", --  516 - 0x204  :   16 - 0x10
    "00011101", --  517 - 0x205  :   29 - 0x1d
    "00000011", --  518 - 0x206  :    3 - 0x3
    "00011011", --  519 - 0x207  :   27 - 0x1b
    "00000000", --  520 - 0x208  :    0 - 0x0
    "00011110", --  521 - 0x209  :   30 - 0x1e
    "00010000", --  522 - 0x20a  :   16 - 0x10
    "00010000", --  523 - 0x20b  :   16 - 0x10
    "00010000", --  524 - 0x20c  :   16 - 0x10
    "00011100", --  525 - 0x20d  :   28 - 0x1c
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00011011", --  527 - 0x20f  :   27 - 0x1b
    "00000011", --  528 - 0x210  :    3 - 0x3
    "00011111", --  529 - 0x211  :   31 - 0x1f
    "00010000", --  530 - 0x212  :   16 - 0x10
    "00010000", --  531 - 0x213  :   16 - 0x10
    "00010000", --  532 - 0x214  :   16 - 0x10
    "00100001", --  533 - 0x215  :   33 - 0x21
    "00101101", --  534 - 0x216  :   45 - 0x2d
    "00101101", --  535 - 0x217  :   45 - 0x2d
    "00101101", --  536 - 0x218  :   45 - 0x2d
    "00101101", --  537 - 0x219  :   45 - 0x2d
    "00101101", --  538 - 0x21a  :   45 - 0x2d
    "00101101", --  539 - 0x21b  :   45 - 0x2d
    "00101101", --  540 - 0x21c  :   45 - 0x2d
    "00101101", --  541 - 0x21d  :   45 - 0x2d
    "00100000", --  542 - 0x21e  :   32 - 0x20
    "00100000", --  543 - 0x21f  :   32 - 0x20
    "00101101", --  544 - 0x220  :   45 - 0x2d -- line 0x11
    "00100000", --  545 - 0x221  :   32 - 0x20
    "00100000", --  546 - 0x222  :   32 - 0x20
    "00100000", --  547 - 0x223  :   32 - 0x20
    "00100000", --  548 - 0x224  :   32 - 0x20
    "00010001", --  549 - 0x225  :   17 - 0x11
    "00000011", --  550 - 0x226  :    3 - 0x3
    "00010001", --  551 - 0x227  :   17 - 0x11
    "00000000", --  552 - 0x228  :    0 - 0x0
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00010001", --  559 - 0x22f  :   17 - 0x11
    "00000011", --  560 - 0x230  :    3 - 0x3
    "00010001", --  561 - 0x231  :   17 - 0x11
    "00100000", --  562 - 0x232  :   32 - 0x20
    "00100000", --  563 - 0x233  :   32 - 0x20
    "00100000", --  564 - 0x234  :   32 - 0x20
    "00100000", --  565 - 0x235  :   32 - 0x20
    "00100000", --  566 - 0x236  :   32 - 0x20
    "00100000", --  567 - 0x237  :   32 - 0x20
    "00100000", --  568 - 0x238  :   32 - 0x20
    "00100000", --  569 - 0x239  :   32 - 0x20
    "00100000", --  570 - 0x23a  :   32 - 0x20
    "00100000", --  571 - 0x23b  :   32 - 0x20
    "00100000", --  572 - 0x23c  :   32 - 0x20
    "00100000", --  573 - 0x23d  :   32 - 0x20
    "00100000", --  574 - 0x23e  :   32 - 0x20
    "00100000", --  575 - 0x23f  :   32 - 0x20
    "00101101", --  576 - 0x240  :   45 - 0x2d -- line 0x12
    "00100000", --  577 - 0x241  :   32 - 0x20
    "00100000", --  578 - 0x242  :   32 - 0x20
    "00100000", --  579 - 0x243  :   32 - 0x20
    "00100000", --  580 - 0x244  :   32 - 0x20
    "00010001", --  581 - 0x245  :   17 - 0x11
    "00000011", --  582 - 0x246  :    3 - 0x3
    "00010001", --  583 - 0x247  :   17 - 0x11
    "00000000", --  584 - 0x248  :    0 - 0x0
    "00011111", --  585 - 0x249  :   31 - 0x1f
    "00010000", --  586 - 0x24a  :   16 - 0x10
    "00010000", --  587 - 0x24b  :   16 - 0x10
    "00010000", --  588 - 0x24c  :   16 - 0x10
    "00011101", --  589 - 0x24d  :   29 - 0x1d
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00010001", --  591 - 0x24f  :   17 - 0x11
    "00000011", --  592 - 0x250  :    3 - 0x3
    "00010001", --  593 - 0x251  :   17 - 0x11
    "00100000", --  594 - 0x252  :   32 - 0x20
    "00100000", --  595 - 0x253  :   32 - 0x20
    "00100000", --  596 - 0x254  :   32 - 0x20
    "00100000", --  597 - 0x255  :   32 - 0x20
    "01100000", --  598 - 0x256  :   96 - 0x60
    "01100001", --  599 - 0x257  :   97 - 0x61
    "00100000", --  600 - 0x258  :   32 - 0x20
    "00100000", --  601 - 0x259  :   32 - 0x20
    "00100000", --  602 - 0x25a  :   32 - 0x20
    "00100000", --  603 - 0x25b  :   32 - 0x20
    "00101101", --  604 - 0x25c  :   45 - 0x2d
    "00101101", --  605 - 0x25d  :   45 - 0x2d
    "00100000", --  606 - 0x25e  :   32 - 0x20
    "00100000", --  607 - 0x25f  :   32 - 0x20
    "00101101", --  608 - 0x260  :   45 - 0x2d -- line 0x13
    "00011111", --  609 - 0x261  :   31 - 0x1f
    "00010000", --  610 - 0x262  :   16 - 0x10
    "00010000", --  611 - 0x263  :   16 - 0x10
    "00010000", --  612 - 0x264  :   16 - 0x10
    "00011100", --  613 - 0x265  :   28 - 0x1c
    "00000011", --  614 - 0x266  :    3 - 0x3
    "00011010", --  615 - 0x267  :   26 - 0x1a
    "00000000", --  616 - 0x268  :    0 - 0x0
    "00011110", --  617 - 0x269  :   30 - 0x1e
    "00010000", --  618 - 0x26a  :   16 - 0x10
    "00010011", --  619 - 0x26b  :   19 - 0x13
    "00010000", --  620 - 0x26c  :   16 - 0x10
    "00011100", --  621 - 0x26d  :   28 - 0x1c
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00011010", --  623 - 0x26f  :   26 - 0x1a
    "00000011", --  624 - 0x270  :    3 - 0x3
    "00011110", --  625 - 0x271  :   30 - 0x1e
    "00010000", --  626 - 0x272  :   16 - 0x10
    "00010000", --  627 - 0x273  :   16 - 0x10
    "00010000", --  628 - 0x274  :   16 - 0x10
    "00011101", --  629 - 0x275  :   29 - 0x1d
    "01100010", --  630 - 0x276  :   98 - 0x62
    "01100011", --  631 - 0x277  :   99 - 0x63
    "00100000", --  632 - 0x278  :   32 - 0x20
    "00100000", --  633 - 0x279  :   32 - 0x20
    "00100000", --  634 - 0x27a  :   32 - 0x20
    "00100000", --  635 - 0x27b  :   32 - 0x20
    "00101101", --  636 - 0x27c  :   45 - 0x2d
    "00101101", --  637 - 0x27d  :   45 - 0x2d
    "00100000", --  638 - 0x27e  :   32 - 0x20
    "00100000", --  639 - 0x27f  :   32 - 0x20
    "00101101", --  640 - 0x280  :   45 - 0x2d -- line 0x14
    "00010001", --  641 - 0x281  :   17 - 0x11
    "00000011", --  642 - 0x282  :    3 - 0x3
    "00000011", --  643 - 0x283  :    3 - 0x3
    "00000011", --  644 - 0x284  :    3 - 0x3
    "00000011", --  645 - 0x285  :    3 - 0x3
    "00000011", --  646 - 0x286  :    3 - 0x3
    "00000011", --  647 - 0x287  :    3 - 0x3
    "00000011", --  648 - 0x288  :    3 - 0x3
    "00000011", --  649 - 0x289  :    3 - 0x3
    "00000011", --  650 - 0x28a  :    3 - 0x3
    "00010001", --  651 - 0x28b  :   17 - 0x11
    "00000011", --  652 - 0x28c  :    3 - 0x3
    "00000011", --  653 - 0x28d  :    3 - 0x3
    "00000011", --  654 - 0x28e  :    3 - 0x3
    "00000011", --  655 - 0x28f  :    3 - 0x3
    "00000011", --  656 - 0x290  :    3 - 0x3
    "00000011", --  657 - 0x291  :    3 - 0x3
    "00000011", --  658 - 0x292  :    3 - 0x3
    "00000011", --  659 - 0x293  :    3 - 0x3
    "00000011", --  660 - 0x294  :    3 - 0x3
    "00010001", --  661 - 0x295  :   17 - 0x11
    "00100000", --  662 - 0x296  :   32 - 0x20
    "00100000", --  663 - 0x297  :   32 - 0x20
    "00100000", --  664 - 0x298  :   32 - 0x20
    "00100000", --  665 - 0x299  :   32 - 0x20
    "00100000", --  666 - 0x29a  :   32 - 0x20
    "00100000", --  667 - 0x29b  :   32 - 0x20
    "00101101", --  668 - 0x29c  :   45 - 0x2d
    "00101101", --  669 - 0x29d  :   45 - 0x2d
    "00100000", --  670 - 0x29e  :   32 - 0x20
    "00100000", --  671 - 0x29f  :   32 - 0x20
    "00101101", --  672 - 0x2a0  :   45 - 0x2d -- line 0x15
    "00010001", --  673 - 0x2a1  :   17 - 0x11
    "00000011", --  674 - 0x2a2  :    3 - 0x3
    "00011001", --  675 - 0x2a3  :   25 - 0x19
    "00010000", --  676 - 0x2a4  :   16 - 0x10
    "00011101", --  677 - 0x2a5  :   29 - 0x1d
    "00000011", --  678 - 0x2a6  :    3 - 0x3
    "00011001", --  679 - 0x2a7  :   25 - 0x19
    "00010000", --  680 - 0x2a8  :   16 - 0x10
    "00011000", --  681 - 0x2a9  :   24 - 0x18
    "00001001", --  682 - 0x2aa  :    9 - 0x9
    "00011010", --  683 - 0x2ab  :   26 - 0x1a
    "00001001", --  684 - 0x2ac  :    9 - 0x9
    "00011001", --  685 - 0x2ad  :   25 - 0x19
    "00010000", --  686 - 0x2ae  :   16 - 0x10
    "00011000", --  687 - 0x2af  :   24 - 0x18
    "00000011", --  688 - 0x2b0  :    3 - 0x3
    "00011111", --  689 - 0x2b1  :   31 - 0x1f
    "00010000", --  690 - 0x2b2  :   16 - 0x10
    "00011000", --  691 - 0x2b3  :   24 - 0x18
    "00000011", --  692 - 0x2b4  :    3 - 0x3
    "00010001", --  693 - 0x2b5  :   17 - 0x11
    "00100000", --  694 - 0x2b6  :   32 - 0x20
    "00100000", --  695 - 0x2b7  :   32 - 0x20
    "00100000", --  696 - 0x2b8  :   32 - 0x20
    "00100000", --  697 - 0x2b9  :   32 - 0x20
    "00100000", --  698 - 0x2ba  :   32 - 0x20
    "00100000", --  699 - 0x2bb  :   32 - 0x20
    "00101101", --  700 - 0x2bc  :   45 - 0x2d
    "00101101", --  701 - 0x2bd  :   45 - 0x2d
    "00100000", --  702 - 0x2be  :   32 - 0x20
    "00100000", --  703 - 0x2bf  :   32 - 0x20
    "00101101", --  704 - 0x2c0  :   45 - 0x2d -- line 0x16
    "00010001", --  705 - 0x2c1  :   17 - 0x11
    "00000001", --  706 - 0x2c2  :    1 - 0x1
    "00000011", --  707 - 0x2c3  :    3 - 0x3
    "00000011", --  708 - 0x2c4  :    3 - 0x3
    "00010001", --  709 - 0x2c5  :   17 - 0x11
    "00000011", --  710 - 0x2c6  :    3 - 0x3
    "00000011", --  711 - 0x2c7  :    3 - 0x3
    "00000011", --  712 - 0x2c8  :    3 - 0x3
    "00000011", --  713 - 0x2c9  :    3 - 0x3
    "00000011", --  714 - 0x2ca  :    3 - 0x3
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000011", --  716 - 0x2cc  :    3 - 0x3
    "00000011", --  717 - 0x2cd  :    3 - 0x3
    "00000011", --  718 - 0x2ce  :    3 - 0x3
    "00000011", --  719 - 0x2cf  :    3 - 0x3
    "00000011", --  720 - 0x2d0  :    3 - 0x3
    "00010001", --  721 - 0x2d1  :   17 - 0x11
    "00000011", --  722 - 0x2d2  :    3 - 0x3
    "00000011", --  723 - 0x2d3  :    3 - 0x3
    "00000001", --  724 - 0x2d4  :    1 - 0x1
    "00010001", --  725 - 0x2d5  :   17 - 0x11
    "00100000", --  726 - 0x2d6  :   32 - 0x20
    "00100000", --  727 - 0x2d7  :   32 - 0x20
    "00100000", --  728 - 0x2d8  :   32 - 0x20
    "00100000", --  729 - 0x2d9  :   32 - 0x20
    "00100000", --  730 - 0x2da  :   32 - 0x20
    "00100000", --  731 - 0x2db  :   32 - 0x20
    "00101101", --  732 - 0x2dc  :   45 - 0x2d
    "00101101", --  733 - 0x2dd  :   45 - 0x2d
    "00100000", --  734 - 0x2de  :   32 - 0x20
    "00100000", --  735 - 0x2df  :   32 - 0x20
    "00101101", --  736 - 0x2e0  :   45 - 0x2d -- line 0x17
    "00010101", --  737 - 0x2e1  :   21 - 0x15
    "00010000", --  738 - 0x2e2  :   16 - 0x10
    "00011101", --  739 - 0x2e3  :   29 - 0x1d
    "00000011", --  740 - 0x2e4  :    3 - 0x3
    "00010001", --  741 - 0x2e5  :   17 - 0x11
    "00000011", --  742 - 0x2e6  :    3 - 0x3
    "00011011", --  743 - 0x2e7  :   27 - 0x1b
    "00000011", --  744 - 0x2e8  :    3 - 0x3
    "00011111", --  745 - 0x2e9  :   31 - 0x1f
    "00010000", --  746 - 0x2ea  :   16 - 0x10
    "00010000", --  747 - 0x2eb  :   16 - 0x10
    "00010000", --  748 - 0x2ec  :   16 - 0x10
    "00011101", --  749 - 0x2ed  :   29 - 0x1d
    "00000011", --  750 - 0x2ee  :    3 - 0x3
    "00011011", --  751 - 0x2ef  :   27 - 0x1b
    "00000011", --  752 - 0x2f0  :    3 - 0x3
    "00010001", --  753 - 0x2f1  :   17 - 0x11
    "00000011", --  754 - 0x2f2  :    3 - 0x3
    "00011111", --  755 - 0x2f3  :   31 - 0x1f
    "00010000", --  756 - 0x2f4  :   16 - 0x10
    "00010100", --  757 - 0x2f5  :   20 - 0x14
    "00100000", --  758 - 0x2f6  :   32 - 0x20
    "00100000", --  759 - 0x2f7  :   32 - 0x20
    "00100000", --  760 - 0x2f8  :   32 - 0x20
    "00100000", --  761 - 0x2f9  :   32 - 0x20
    "00100000", --  762 - 0x2fa  :   32 - 0x20
    "00100000", --  763 - 0x2fb  :   32 - 0x20
    "00101101", --  764 - 0x2fc  :   45 - 0x2d
    "00101101", --  765 - 0x2fd  :   45 - 0x2d
    "00100000", --  766 - 0x2fe  :   32 - 0x20
    "00100000", --  767 - 0x2ff  :   32 - 0x20
    "00101101", --  768 - 0x300  :   45 - 0x2d -- line 0x18
    "00010101", --  769 - 0x301  :   21 - 0x15
    "00010000", --  770 - 0x302  :   16 - 0x10
    "00011100", --  771 - 0x303  :   28 - 0x1c
    "00000011", --  772 - 0x304  :    3 - 0x3
    "00011010", --  773 - 0x305  :   26 - 0x1a
    "00000011", --  774 - 0x306  :    3 - 0x3
    "00010001", --  775 - 0x307  :   17 - 0x11
    "00000011", --  776 - 0x308  :    3 - 0x3
    "00011110", --  777 - 0x309  :   30 - 0x1e
    "00010000", --  778 - 0x30a  :   16 - 0x10
    "00010011", --  779 - 0x30b  :   19 - 0x13
    "00010000", --  780 - 0x30c  :   16 - 0x10
    "00011100", --  781 - 0x30d  :   28 - 0x1c
    "00000011", --  782 - 0x30e  :    3 - 0x3
    "00010001", --  783 - 0x30f  :   17 - 0x11
    "00000011", --  784 - 0x310  :    3 - 0x3
    "00011010", --  785 - 0x311  :   26 - 0x1a
    "00000011", --  786 - 0x312  :    3 - 0x3
    "00011110", --  787 - 0x313  :   30 - 0x1e
    "00010000", --  788 - 0x314  :   16 - 0x10
    "00010100", --  789 - 0x315  :   20 - 0x14
    "00100000", --  790 - 0x316  :   32 - 0x20
    "00111100", --  791 - 0x317  :   60 - 0x3c
    "00111101", --  792 - 0x318  :   61 - 0x3d
    "00111100", --  793 - 0x319  :   60 - 0x3c
    "00111101", --  794 - 0x31a  :   61 - 0x3d
    "00101101", --  795 - 0x31b  :   45 - 0x2d
    "00101101", --  796 - 0x31c  :   45 - 0x2d
    "00101101", --  797 - 0x31d  :   45 - 0x2d
    "00100000", --  798 - 0x31e  :   32 - 0x20
    "00100000", --  799 - 0x31f  :   32 - 0x20
    "00101101", --  800 - 0x320  :   45 - 0x2d -- line 0x19
    "00010001", --  801 - 0x321  :   17 - 0x11
    "00000011", --  802 - 0x322  :    3 - 0x3
    "00000011", --  803 - 0x323  :    3 - 0x3
    "00000011", --  804 - 0x324  :    3 - 0x3
    "00000011", --  805 - 0x325  :    3 - 0x3
    "00000011", --  806 - 0x326  :    3 - 0x3
    "00010001", --  807 - 0x327  :   17 - 0x11
    "00000011", --  808 - 0x328  :    3 - 0x3
    "00000011", --  809 - 0x329  :    3 - 0x3
    "00000011", --  810 - 0x32a  :    3 - 0x3
    "00010001", --  811 - 0x32b  :   17 - 0x11
    "00000011", --  812 - 0x32c  :    3 - 0x3
    "00000011", --  813 - 0x32d  :    3 - 0x3
    "00000011", --  814 - 0x32e  :    3 - 0x3
    "00010001", --  815 - 0x32f  :   17 - 0x11
    "00000011", --  816 - 0x330  :    3 - 0x3
    "00000011", --  817 - 0x331  :    3 - 0x3
    "00000011", --  818 - 0x332  :    3 - 0x3
    "00000011", --  819 - 0x333  :    3 - 0x3
    "00000011", --  820 - 0x334  :    3 - 0x3
    "00010001", --  821 - 0x335  :   17 - 0x11
    "00100000", --  822 - 0x336  :   32 - 0x20
    "00111110", --  823 - 0x337  :   62 - 0x3e
    "00111111", --  824 - 0x338  :   63 - 0x3f
    "00111110", --  825 - 0x339  :   62 - 0x3e
    "00111111", --  826 - 0x33a  :   63 - 0x3f
    "00101101", --  827 - 0x33b  :   45 - 0x2d
    "00101101", --  828 - 0x33c  :   45 - 0x2d
    "00101101", --  829 - 0x33d  :   45 - 0x2d
    "00100000", --  830 - 0x33e  :   32 - 0x20
    "00100000", --  831 - 0x33f  :   32 - 0x20
    "00101101", --  832 - 0x340  :   45 - 0x2d -- line 0x1a
    "00010001", --  833 - 0x341  :   17 - 0x11
    "00000011", --  834 - 0x342  :    3 - 0x3
    "00011001", --  835 - 0x343  :   25 - 0x19
    "00010000", --  836 - 0x344  :   16 - 0x10
    "00010000", --  837 - 0x345  :   16 - 0x10
    "00010000", --  838 - 0x346  :   16 - 0x10
    "00010010", --  839 - 0x347  :   18 - 0x12
    "00010000", --  840 - 0x348  :   16 - 0x10
    "00011000", --  841 - 0x349  :   24 - 0x18
    "00000011", --  842 - 0x34a  :    3 - 0x3
    "00011010", --  843 - 0x34b  :   26 - 0x1a
    "00000011", --  844 - 0x34c  :    3 - 0x3
    "00011001", --  845 - 0x34d  :   25 - 0x19
    "00010000", --  846 - 0x34e  :   16 - 0x10
    "00010010", --  847 - 0x34f  :   18 - 0x12
    "00010000", --  848 - 0x350  :   16 - 0x10
    "00010000", --  849 - 0x351  :   16 - 0x10
    "00010000", --  850 - 0x352  :   16 - 0x10
    "00011000", --  851 - 0x353  :   24 - 0x18
    "00000011", --  852 - 0x354  :    3 - 0x3
    "00010001", --  853 - 0x355  :   17 - 0x11
    "00100000", --  854 - 0x356  :   32 - 0x20
    "00100000", --  855 - 0x357  :   32 - 0x20
    "00100000", --  856 - 0x358  :   32 - 0x20
    "00100000", --  857 - 0x359  :   32 - 0x20
    "00100000", --  858 - 0x35a  :   32 - 0x20
    "00100000", --  859 - 0x35b  :   32 - 0x20
    "00101101", --  860 - 0x35c  :   45 - 0x2d
    "00101101", --  861 - 0x35d  :   45 - 0x2d
    "00100000", --  862 - 0x35e  :   32 - 0x20
    "00100000", --  863 - 0x35f  :   32 - 0x20
    "00101101", --  864 - 0x360  :   45 - 0x2d -- line 0x1b
    "00010001", --  865 - 0x361  :   17 - 0x11
    "00000011", --  866 - 0x362  :    3 - 0x3
    "00000011", --  867 - 0x363  :    3 - 0x3
    "00000011", --  868 - 0x364  :    3 - 0x3
    "00000011", --  869 - 0x365  :    3 - 0x3
    "00000011", --  870 - 0x366  :    3 - 0x3
    "00000011", --  871 - 0x367  :    3 - 0x3
    "00000011", --  872 - 0x368  :    3 - 0x3
    "00000011", --  873 - 0x369  :    3 - 0x3
    "00000011", --  874 - 0x36a  :    3 - 0x3
    "00000011", --  875 - 0x36b  :    3 - 0x3
    "00000011", --  876 - 0x36c  :    3 - 0x3
    "00000011", --  877 - 0x36d  :    3 - 0x3
    "00000011", --  878 - 0x36e  :    3 - 0x3
    "00000011", --  879 - 0x36f  :    3 - 0x3
    "00000011", --  880 - 0x370  :    3 - 0x3
    "00000011", --  881 - 0x371  :    3 - 0x3
    "00000011", --  882 - 0x372  :    3 - 0x3
    "00000011", --  883 - 0x373  :    3 - 0x3
    "00000011", --  884 - 0x374  :    3 - 0x3
    "00010001", --  885 - 0x375  :   17 - 0x11
    "00100000", --  886 - 0x376  :   32 - 0x20
    "00100000", --  887 - 0x377  :   32 - 0x20
    "00100000", --  888 - 0x378  :   32 - 0x20
    "00100000", --  889 - 0x379  :   32 - 0x20
    "00100000", --  890 - 0x37a  :   32 - 0x20
    "00100000", --  891 - 0x37b  :   32 - 0x20
    "00101101", --  892 - 0x37c  :   45 - 0x2d
    "00101101", --  893 - 0x37d  :   45 - 0x2d
    "00100000", --  894 - 0x37e  :   32 - 0x20
    "00100000", --  895 - 0x37f  :   32 - 0x20
    "00101101", --  896 - 0x380  :   45 - 0x2d -- line 0x1c
    "00011110", --  897 - 0x381  :   30 - 0x1e
    "00010000", --  898 - 0x382  :   16 - 0x10
    "00010000", --  899 - 0x383  :   16 - 0x10
    "00010000", --  900 - 0x384  :   16 - 0x10
    "00010000", --  901 - 0x385  :   16 - 0x10
    "00010000", --  902 - 0x386  :   16 - 0x10
    "00010000", --  903 - 0x387  :   16 - 0x10
    "00010000", --  904 - 0x388  :   16 - 0x10
    "00010000", --  905 - 0x389  :   16 - 0x10
    "00010000", --  906 - 0x38a  :   16 - 0x10
    "00010000", --  907 - 0x38b  :   16 - 0x10
    "00010000", --  908 - 0x38c  :   16 - 0x10
    "00010000", --  909 - 0x38d  :   16 - 0x10
    "00010000", --  910 - 0x38e  :   16 - 0x10
    "00010000", --  911 - 0x38f  :   16 - 0x10
    "00010000", --  912 - 0x390  :   16 - 0x10
    "00010000", --  913 - 0x391  :   16 - 0x10
    "00010000", --  914 - 0x392  :   16 - 0x10
    "00010000", --  915 - 0x393  :   16 - 0x10
    "00010000", --  916 - 0x394  :   16 - 0x10
    "00011100", --  917 - 0x395  :   28 - 0x1c
    "00100000", --  918 - 0x396  :   32 - 0x20
    "00100000", --  919 - 0x397  :   32 - 0x20
    "00100000", --  920 - 0x398  :   32 - 0x20
    "00100000", --  921 - 0x399  :   32 - 0x20
    "00100000", --  922 - 0x39a  :   32 - 0x20
    "00100000", --  923 - 0x39b  :   32 - 0x20
    "00100000", --  924 - 0x39c  :   32 - 0x20
    "00100000", --  925 - 0x39d  :   32 - 0x20
    "00100000", --  926 - 0x39e  :   32 - 0x20
    "00100000", --  927 - 0x39f  :   32 - 0x20
    "00100000", --  928 - 0x3a0  :   32 - 0x20 -- line 0x1d
    "00100000", --  929 - 0x3a1  :   32 - 0x20
    "00100000", --  930 - 0x3a2  :   32 - 0x20
    "00100000", --  931 - 0x3a3  :   32 - 0x20
    "00100000", --  932 - 0x3a4  :   32 - 0x20
    "00100000", --  933 - 0x3a5  :   32 - 0x20
    "00100000", --  934 - 0x3a6  :   32 - 0x20
    "00100000", --  935 - 0x3a7  :   32 - 0x20
    "00100000", --  936 - 0x3a8  :   32 - 0x20
    "00100000", --  937 - 0x3a9  :   32 - 0x20
    "00100000", --  938 - 0x3aa  :   32 - 0x20
    "00100000", --  939 - 0x3ab  :   32 - 0x20
    "00100000", --  940 - 0x3ac  :   32 - 0x20
    "00100000", --  941 - 0x3ad  :   32 - 0x20
    "00100000", --  942 - 0x3ae  :   32 - 0x20
    "00100000", --  943 - 0x3af  :   32 - 0x20
    "00100000", --  944 - 0x3b0  :   32 - 0x20
    "00100000", --  945 - 0x3b1  :   32 - 0x20
    "00100000", --  946 - 0x3b2  :   32 - 0x20
    "00100000", --  947 - 0x3b3  :   32 - 0x20
    "00100000", --  948 - 0x3b4  :   32 - 0x20
    "00100000", --  949 - 0x3b5  :   32 - 0x20
    "00100000", --  950 - 0x3b6  :   32 - 0x20
    "00100000", --  951 - 0x3b7  :   32 - 0x20
    "00100000", --  952 - 0x3b8  :   32 - 0x20
    "00100000", --  953 - 0x3b9  :   32 - 0x20
    "00100000", --  954 - 0x3ba  :   32 - 0x20
    "00100000", --  955 - 0x3bb  :   32 - 0x20
    "00100000", --  956 - 0x3bc  :   32 - 0x20
    "00100000", --  957 - 0x3bd  :   32 - 0x20
    "00100000", --  958 - 0x3be  :   32 - 0x20
    "00100000", --  959 - 0x3bf  :   32 - 0x20
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "01010101", --  961 - 0x3c1  :   85 - 0x55
    "01010101", --  962 - 0x3c2  :   85 - 0x55
    "01010101", --  963 - 0x3c3  :   85 - 0x55
    "01010101", --  964 - 0x3c4  :   85 - 0x55
    "00010001", --  965 - 0x3c5  :   17 - 0x11
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "01010101", --  968 - 0x3c8  :   85 - 0x55
    "01010101", --  969 - 0x3c9  :   85 - 0x55
    "01010101", --  970 - 0x3ca  :   85 - 0x55
    "01010101", --  971 - 0x3cb  :   85 - 0x55
    "01010101", --  972 - 0x3cc  :   85 - 0x55
    "00010001", --  973 - 0x3cd  :   17 - 0x11
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "01010101", --  977 - 0x3d1  :   85 - 0x55
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "00010001", --  981 - 0x3d5  :   17 - 0x11
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010001", --  989 - 0x3dd  :   81 - 0x51
    "01010000", --  990 - 0x3de  :   80 - 0x50
    "01010000", --  991 - 0x3df  :   80 - 0x50
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "10010101", --  997 - 0x3e5  :  149 - 0x95
    "00000101", --  998 - 0x3e6  :    5 - 0x5
    "00000101", --  999 - 0x3e7  :    5 - 0x5
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "01010101", -- 1002 - 0x3ea  :   85 - 0x55
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "00010001", -- 1005 - 0x3ed  :   17 - 0x11
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "01010101", -- 1010 - 0x3f2  :   85 - 0x55
    "01010101", -- 1011 - 0x3f3  :   85 - 0x55
    "01010101", -- 1012 - 0x3f4  :   85 - 0x55
    "01010101", -- 1013 - 0x3f5  :   85 - 0x55
    "01010101", -- 1014 - 0x3f6  :   85 - 0x55
    "01010101", -- 1015 - 0x3f7  :   85 - 0x55
    "01010101", -- 1016 - 0x3f8  :   85 - 0x55
    "01010101", -- 1017 - 0x3f9  :   85 - 0x55
    "01010101", -- 1018 - 0x3fa  :   85 - 0x55
    "01010101", -- 1019 - 0x3fb  :   85 - 0x55
    "01010101", -- 1020 - 0x3fc  :   85 - 0x55
    "01010101", -- 1021 - 0x3fd  :   85 - 0x55
    "01010101", -- 1022 - 0x3fe  :   85 - 0x55
    "01010101"  -- 1023 - 0x3ff  :   85 - 0x55
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
