--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_color0 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_color0;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00001111", --    1 -  0x1  :   15 - 0xf
    "00000100", --    2 -  0x2  :    4 - 0x4
    "00000011", --    3 -  0x3  :    3 - 0x3
    "00000011", --    4 -  0x4  :    3 - 0x3
    "00000011", --    5 -  0x5  :    3 - 0x3
    "00000100", --    6 -  0x6  :    4 - 0x4
    "00111010", --    7 -  0x7  :   58 - 0x3a
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "11000110", --   10 -  0xa  :  198 - 0xc6
    "11001011", --   11 -  0xb  :  203 - 0xcb
    "11011100", --   12 -  0xc  :  220 - 0xdc
    "00111010", --   13 -  0xd  :   58 - 0x3a
    "10011010", --   14 -  0xe  :  154 - 0x9a
    "10000001", --   15 -  0xf  :  129 - 0x81
    "01000101", --   16 - 0x10  :   69 - 0x45 -- Sprite 0x2
    "10000111", --   17 - 0x11  :  135 - 0x87
    "10000011", --   18 - 0x12  :  131 - 0x83
    "10000001", --   19 - 0x13  :  129 - 0x81
    "10000001", --   20 - 0x14  :  129 - 0x81
    "10000001", --   21 - 0x15  :  129 - 0x81
    "01000001", --   22 - 0x16  :   65 - 0x41
    "00100001", --   23 - 0x17  :   33 - 0x21
    "01111111", --   24 - 0x18  :  127 - 0x7f -- Sprite 0x3
    "01111110", --   25 - 0x19  :  126 - 0x7e
    "11111100", --   26 - 0x1a  :  252 - 0xfc
    "00111000", --   27 - 0x1b  :   56 - 0x38
    "00011000", --   28 - 0x1c  :   24 - 0x18
    "10001100", --   29 - 0x1d  :  140 - 0x8c
    "11000100", --   30 - 0x1e  :  196 - 0xc4
    "11111100", --   31 - 0x1f  :  252 - 0xfc
    "00100011", --   32 - 0x20  :   35 - 0x23 -- Sprite 0x4
    "00100011", --   33 - 0x21  :   35 - 0x23
    "00100001", --   34 - 0x22  :   33 - 0x21
    "00100000", --   35 - 0x23  :   32 - 0x20
    "00010011", --   36 - 0x24  :   19 - 0x13
    "00001100", --   37 - 0x25  :   12 - 0xc
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "11111100", --   40 - 0x28  :  252 - 0xfc -- Sprite 0x5
    "11111100", --   41 - 0x29  :  252 - 0xfc
    "11111100", --   42 - 0x2a  :  252 - 0xfc
    "11111100", --   43 - 0x2b  :  252 - 0xfc
    "10010000", --   44 - 0x2c  :  144 - 0x90
    "10010000", --   45 - 0x2d  :  144 - 0x90
    "10001000", --   46 - 0x2e  :  136 - 0x88
    "11111000", --   47 - 0x2f  :  248 - 0xf8
    "00100011", --   48 - 0x30  :   35 - 0x23 -- Sprite 0x6
    "00100011", --   49 - 0x31  :   35 - 0x23
    "00100001", --   50 - 0x32  :   33 - 0x21
    "00100000", --   51 - 0x33  :   32 - 0x20
    "00010011", --   52 - 0x34  :   19 - 0x13
    "00001101", --   53 - 0x35  :   13 - 0xd
    "00000010", --   54 - 0x36  :    2 - 0x2
    "00000001", --   55 - 0x37  :    1 - 0x1
    "11111100", --   56 - 0x38  :  252 - 0xfc -- Sprite 0x7
    "11111100", --   57 - 0x39  :  252 - 0xfc
    "11111100", --   58 - 0x3a  :  252 - 0xfc
    "11111100", --   59 - 0x3b  :  252 - 0xfc
    "10100100", --   60 - 0x3c  :  164 - 0xa4
    "00100100", --   61 - 0x3d  :   36 - 0x24
    "01010010", --   62 - 0x3e  :   82 - 0x52
    "11101110", --   63 - 0x3f  :  238 - 0xee
    "00100011", --   64 - 0x40  :   35 - 0x23 -- Sprite 0x8
    "00100011", --   65 - 0x41  :   35 - 0x23
    "00100001", --   66 - 0x42  :   33 - 0x21
    "00100000", --   67 - 0x43  :   32 - 0x20
    "00010011", --   68 - 0x44  :   19 - 0x13
    "00001101", --   69 - 0x45  :   13 - 0xd
    "00000001", --   70 - 0x46  :    1 - 0x1
    "00000001", --   71 - 0x47  :    1 - 0x1
    "11111110", --   72 - 0x48  :  254 - 0xfe -- Sprite 0x9
    "11111110", --   73 - 0x49  :  254 - 0xfe
    "11111110", --   74 - 0x4a  :  254 - 0xfe
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "10010001", --   76 - 0x4c  :  145 - 0x91
    "00101111", --   77 - 0x4d  :   47 - 0x2f
    "01000000", --   78 - 0x4e  :   64 - 0x40
    "11100000", --   79 - 0x4f  :  224 - 0xe0
    "00100011", --   80 - 0x50  :   35 - 0x23 -- Sprite 0xa
    "00100011", --   81 - 0x51  :   35 - 0x23
    "00100001", --   82 - 0x52  :   33 - 0x21
    "00100000", --   83 - 0x53  :   32 - 0x20
    "00010011", --   84 - 0x54  :   19 - 0x13
    "00001110", --   85 - 0x55  :   14 - 0xe
    "00000001", --   86 - 0x56  :    1 - 0x1
    "00000000", --   87 - 0x57  :    0 - 0x0
    "11111110", --   88 - 0x58  :  254 - 0xfe -- Sprite 0xb
    "11111110", --   89 - 0x59  :  254 - 0xfe
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111100", --   91 - 0x5b  :  252 - 0xfc
    "00100100", --   92 - 0x5c  :   36 - 0x24
    "00100010", --   93 - 0x5d  :   34 - 0x22
    "11010010", --   94 - 0x5e  :  210 - 0xd2
    "00001111", --   95 - 0x5f  :   15 - 0xf
    "01111111", --   96 - 0x60  :  127 - 0x7f -- Sprite 0xc
    "01111110", --   97 - 0x61  :  126 - 0x7e
    "11111100", --   98 - 0x62  :  252 - 0xfc
    "00000010", --   99 - 0x63  :    2 - 0x2
    "00000100", --  100 - 0x64  :    4 - 0x4
    "11111100", --  101 - 0x65  :  252 - 0xfc
    "11111100", --  102 - 0x66  :  252 - 0xfc
    "11111110", --  103 - 0x67  :  254 - 0xfe
    "01000101", --  104 - 0x68  :   69 - 0x45 -- Sprite 0xd
    "10000111", --  105 - 0x69  :  135 - 0x87
    "10000011", --  106 - 0x6a  :  131 - 0x83
    "10000010", --  107 - 0x6b  :  130 - 0x82
    "10000010", --  108 - 0x6c  :  130 - 0x82
    "10000100", --  109 - 0x6d  :  132 - 0x84
    "01000100", --  110 - 0x6e  :   68 - 0x44
    "00100100", --  111 - 0x6f  :   36 - 0x24
    "01111111", --  112 - 0x70  :  127 - 0x7f -- Sprite 0xe
    "01111110", --  113 - 0x71  :  126 - 0x7e
    "11111100", --  114 - 0x72  :  252 - 0xfc
    "11111000", --  115 - 0x73  :  248 - 0xf8
    "01111000", --  116 - 0x74  :  120 - 0x78
    "01111100", --  117 - 0x75  :  124 - 0x7c
    "11111100", --  118 - 0x76  :  252 - 0xfc
    "11111110", --  119 - 0x77  :  254 - 0xfe
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Sprite 0xf
    "00001111", --  121 - 0x79  :   15 - 0xf
    "00000100", --  122 - 0x7a  :    4 - 0x4
    "00000011", --  123 - 0x7b  :    3 - 0x3
    "00000011", --  124 - 0x7c  :    3 - 0x3
    "00000011", --  125 - 0x7d  :    3 - 0x3
    "00000100", --  126 - 0x7e  :    4 - 0x4
    "00000010", --  127 - 0x7f  :    2 - 0x2
    "00000111", --  128 - 0x80  :    7 - 0x7 -- Sprite 0x10
    "00001100", --  129 - 0x81  :   12 - 0xc
    "00010000", --  130 - 0x82  :   16 - 0x10
    "00010000", --  131 - 0x83  :   16 - 0x10
    "00010000", --  132 - 0x84  :   16 - 0x10
    "00100000", --  133 - 0x85  :   32 - 0x20
    "00100000", --  134 - 0x86  :   32 - 0x20
    "00100001", --  135 - 0x87  :   33 - 0x21
    "11111111", --  136 - 0x88  :  255 - 0xff -- Sprite 0x11
    "01111110", --  137 - 0x89  :  126 - 0x7e
    "01111100", --  138 - 0x8a  :  124 - 0x7c
    "01111000", --  139 - 0x8b  :  120 - 0x78
    "01011000", --  140 - 0x8c  :   88 - 0x58
    "10001100", --  141 - 0x8d  :  140 - 0x8c
    "11000100", --  142 - 0x8e  :  196 - 0xc4
    "11111100", --  143 - 0x8f  :  252 - 0xfc
    "00100011", --  144 - 0x90  :   35 - 0x23 -- Sprite 0x12
    "00100011", --  145 - 0x91  :   35 - 0x23
    "00100001", --  146 - 0x92  :   33 - 0x21
    "00100000", --  147 - 0x93  :   32 - 0x20
    "00010011", --  148 - 0x94  :   19 - 0x13
    "00001100", --  149 - 0x95  :   12 - 0xc
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000001", --  152 - 0x98  :    1 - 0x1 -- Sprite 0x13
    "00000001", --  153 - 0x99  :    1 - 0x1
    "00000011", --  154 - 0x9a  :    3 - 0x3
    "00000100", --  155 - 0x9b  :    4 - 0x4
    "00001000", --  156 - 0x9c  :    8 - 0x8
    "00010000", --  157 - 0x9d  :   16 - 0x10
    "00010000", --  158 - 0x9e  :   16 - 0x10
    "00100000", --  159 - 0x9f  :   32 - 0x20
    "01111111", --  160 - 0xa0  :  127 - 0x7f -- Sprite 0x14
    "11111110", --  161 - 0xa1  :  254 - 0xfe
    "00000110", --  162 - 0xa2  :    6 - 0x6
    "00000001", --  163 - 0xa3  :    1 - 0x1
    "00000001", --  164 - 0xa4  :    1 - 0x1
    "00000001", --  165 - 0xa5  :    1 - 0x1
    "00000111", --  166 - 0xa6  :    7 - 0x7
    "11111110", --  167 - 0xa7  :  254 - 0xfe
    "00000101", --  168 - 0xa8  :    5 - 0x5 -- Sprite 0x15
    "00000101", --  169 - 0xa9  :    5 - 0x5
    "00000111", --  170 - 0xaa  :    7 - 0x7
    "00000100", --  171 - 0xab  :    4 - 0x4
    "00000100", --  172 - 0xac  :    4 - 0x4
    "00001111", --  173 - 0xad  :   15 - 0xf
    "00110000", --  174 - 0xae  :   48 - 0x30
    "01000000", --  175 - 0xaf  :   64 - 0x40
    "11111100", --  176 - 0xb0  :  252 - 0xfc -- Sprite 0x16
    "11111000", --  177 - 0xb1  :  248 - 0xf8
    "11110000", --  178 - 0xb2  :  240 - 0xf0
    "11100000", --  179 - 0xb3  :  224 - 0xe0
    "01100000", --  180 - 0xb4  :   96 - 0x60
    "11110000", --  181 - 0xb5  :  240 - 0xf0
    "00011100", --  182 - 0xb6  :   28 - 0x1c
    "00000010", --  183 - 0xb7  :    2 - 0x2
    "10000000", --  184 - 0xb8  :  128 - 0x80 -- Sprite 0x17
    "10000000", --  185 - 0xb9  :  128 - 0x80
    "10000000", --  186 - 0xba  :  128 - 0x80
    "10000011", --  187 - 0xbb  :  131 - 0x83
    "01001111", --  188 - 0xbc  :   79 - 0x4f
    "00110010", --  189 - 0xbd  :   50 - 0x32
    "00000010", --  190 - 0xbe  :    2 - 0x2
    "00000011", --  191 - 0xbf  :    3 - 0x3
    "00000010", --  192 - 0xc0  :    2 - 0x2 -- Sprite 0x18
    "00000001", --  193 - 0xc1  :    1 - 0x1
    "00000010", --  194 - 0xc2  :    2 - 0x2
    "11111100", --  195 - 0xc3  :  252 - 0xfc
    "11000000", --  196 - 0xc4  :  192 - 0xc0
    "01000000", --  197 - 0xc5  :   64 - 0x40
    "00100000", --  198 - 0xc6  :   32 - 0x20
    "11100000", --  199 - 0xc7  :  224 - 0xe0
    "00001011", --  200 - 0xc8  :   11 - 0xb -- Sprite 0x19
    "00001011", --  201 - 0xc9  :   11 - 0xb
    "00001111", --  202 - 0xca  :   15 - 0xf
    "00001001", --  203 - 0xcb  :    9 - 0x9
    "00001000", --  204 - 0xcc  :    8 - 0x8
    "00001001", --  205 - 0xcd  :    9 - 0x9
    "00001111", --  206 - 0xce  :   15 - 0xf
    "00110000", --  207 - 0xcf  :   48 - 0x30
    "11111000", --  208 - 0xd0  :  248 - 0xf8 -- Sprite 0x1a
    "11110000", --  209 - 0xd1  :  240 - 0xf0
    "11100000", --  210 - 0xd2  :  224 - 0xe0
    "11000000", --  211 - 0xd3  :  192 - 0xc0
    "11000000", --  212 - 0xd4  :  192 - 0xc0
    "11000000", --  213 - 0xd5  :  192 - 0xc0
    "11111000", --  214 - 0xd6  :  248 - 0xf8
    "00011111", --  215 - 0xd7  :   31 - 0x1f
    "01000000", --  216 - 0xd8  :   64 - 0x40 -- Sprite 0x1b
    "01000000", --  217 - 0xd9  :   64 - 0x40
    "10000000", --  218 - 0xda  :  128 - 0x80
    "10000000", --  219 - 0xdb  :  128 - 0x80
    "01000000", --  220 - 0xdc  :   64 - 0x40
    "00111111", --  221 - 0xdd  :   63 - 0x3f
    "00000100", --  222 - 0xde  :    4 - 0x4
    "00000111", --  223 - 0xdf  :    7 - 0x7
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0x1c
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "01000000", --  230 - 0xe6  :   64 - 0x40
    "11000000", --  231 - 0xe7  :  192 - 0xc0
    "11000000", --  232 - 0xe8  :  192 - 0xc0 -- Sprite 0x1d
    "00100000", --  233 - 0xe9  :   32 - 0x20
    "00100000", --  234 - 0xea  :   32 - 0x20
    "00100000", --  235 - 0xeb  :   32 - 0x20
    "01000000", --  236 - 0xec  :   64 - 0x40
    "10000000", --  237 - 0xed  :  128 - 0x80
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "01111111", --  240 - 0xf0  :  127 - 0x7f -- Sprite 0x1e
    "01100010", --  241 - 0xf1  :   98 - 0x62
    "11000100", --  242 - 0xf2  :  196 - 0xc4
    "00011000", --  243 - 0xf3  :   24 - 0x18
    "00111100", --  244 - 0xf4  :   60 - 0x3c
    "11111110", --  245 - 0xf5  :  254 - 0xfe
    "11111110", --  246 - 0xf6  :  254 - 0xfe
    "11111110", --  247 - 0xf7  :  254 - 0xfe
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Sprite 0x1f
    "00111000", --  249 - 0xf9  :   56 - 0x38
    "11000110", --  250 - 0xfa  :  198 - 0xc6
    "11001011", --  251 - 0xfb  :  203 - 0xcb
    "11011100", --  252 - 0xfc  :  220 - 0xdc
    "00111010", --  253 - 0xfd  :   58 - 0x3a
    "10011010", --  254 - 0xfe  :  154 - 0x9a
    "11100001", --  255 - 0xff  :  225 - 0xe1
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00011100", --  257 - 0x101  :   28 - 0x1c
    "00010011", --  258 - 0x102  :   19 - 0x13
    "00001000", --  259 - 0x103  :    8 - 0x8
    "00010000", --  260 - 0x104  :   16 - 0x10
    "00001000", --  261 - 0x105  :    8 - 0x8
    "00010000", --  262 - 0x106  :   16 - 0x10
    "00010000", --  263 - 0x107  :   16 - 0x10
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00111000", --  265 - 0x109  :   56 - 0x38
    "11001000", --  266 - 0x10a  :  200 - 0xc8
    "00010000", --  267 - 0x10b  :   16 - 0x10
    "00001000", --  268 - 0x10c  :    8 - 0x8
    "00010000", --  269 - 0x10d  :   16 - 0x10
    "00001000", --  270 - 0x10e  :    8 - 0x8
    "00001000", --  271 - 0x10f  :    8 - 0x8
    "00001000", --  272 - 0x110  :    8 - 0x8 -- Sprite 0x22
    "00011100", --  273 - 0x111  :   28 - 0x1c
    "00100111", --  274 - 0x112  :   39 - 0x27
    "00101111", --  275 - 0x113  :   47 - 0x2f
    "00011111", --  276 - 0x114  :   31 - 0x1f
    "00001111", --  277 - 0x115  :   15 - 0xf
    "00001111", --  278 - 0x116  :   15 - 0xf
    "00001111", --  279 - 0x117  :   15 - 0xf
    "00010000", --  280 - 0x118  :   16 - 0x10 -- Sprite 0x23
    "00111100", --  281 - 0x119  :   60 - 0x3c
    "11000010", --  282 - 0x11a  :  194 - 0xc2
    "10000010", --  283 - 0x11b  :  130 - 0x82
    "10000010", --  284 - 0x11c  :  130 - 0x82
    "10000010", --  285 - 0x11d  :  130 - 0x82
    "00010010", --  286 - 0x11e  :   18 - 0x12
    "00011100", --  287 - 0x11f  :   28 - 0x1c
    "00001111", --  288 - 0x120  :   15 - 0xf -- Sprite 0x24
    "00001110", --  289 - 0x121  :   14 - 0xe
    "00010100", --  290 - 0x122  :   20 - 0x14
    "00010100", --  291 - 0x123  :   20 - 0x14
    "00010010", --  292 - 0x124  :   18 - 0x12
    "00100101", --  293 - 0x125  :   37 - 0x25
    "01000100", --  294 - 0x126  :   68 - 0x44
    "00111000", --  295 - 0x127  :   56 - 0x38
    "00010000", --  296 - 0x128  :   16 - 0x10 -- Sprite 0x25
    "00010000", --  297 - 0x129  :   16 - 0x10
    "00010000", --  298 - 0x12a  :   16 - 0x10
    "00101100", --  299 - 0x12b  :   44 - 0x2c
    "01000100", --  300 - 0x12c  :   68 - 0x44
    "11000100", --  301 - 0x12d  :  196 - 0xc4
    "00111000", --  302 - 0x12e  :   56 - 0x38
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Sprite 0x27
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00100000", --  328 - 0x148  :   32 - 0x20 -- Sprite 0x29
    "00100000", --  329 - 0x149  :   32 - 0x20
    "00100000", --  330 - 0x14a  :   32 - 0x20
    "00100000", --  331 - 0x14b  :   32 - 0x20
    "00010011", --  332 - 0x14c  :   19 - 0x13
    "00001101", --  333 - 0x14d  :   13 - 0xd
    "00000010", --  334 - 0x14e  :    2 - 0x2
    "00000001", --  335 - 0x14f  :    1 - 0x1
    "00100000", --  336 - 0x150  :   32 - 0x20 -- Sprite 0x2a
    "00100000", --  337 - 0x151  :   32 - 0x20
    "00100000", --  338 - 0x152  :   32 - 0x20
    "00100000", --  339 - 0x153  :   32 - 0x20
    "00010011", --  340 - 0x154  :   19 - 0x13
    "00001101", --  341 - 0x155  :   13 - 0xd
    "00000001", --  342 - 0x156  :    1 - 0x1
    "00000001", --  343 - 0x157  :    1 - 0x1
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Sprite 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00111100", --  360 - 0x168  :   60 - 0x3c -- Sprite 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "10000001", --  362 - 0x16a  :  129 - 0x81
    "10011001", --  363 - 0x16b  :  153 - 0x99
    "10011001", --  364 - 0x16c  :  153 - 0x99
    "10000001", --  365 - 0x16d  :  129 - 0x81
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00111100", --  367 - 0x16f  :   60 - 0x3c
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "10011111", --  376 - 0x178  :  159 - 0x9f -- Sprite 0x2f
    "10011110", --  377 - 0x179  :  158 - 0x9e
    "10011100", --  378 - 0x17a  :  156 - 0x9c
    "00011000", --  379 - 0x17b  :   24 - 0x18
    "00111000", --  380 - 0x17c  :   56 - 0x38
    "11111100", --  381 - 0x17d  :  252 - 0xfc
    "11111100", --  382 - 0x17e  :  252 - 0xfc
    "11111100", --  383 - 0x17f  :  252 - 0xfc
    "01111111", --  384 - 0x180  :  127 - 0x7f -- Sprite 0x30
    "01111110", --  385 - 0x181  :  126 - 0x7e
    "11111100", --  386 - 0x182  :  252 - 0xfc
    "00111000", --  387 - 0x183  :   56 - 0x38
    "00111000", --  388 - 0x184  :   56 - 0x38
    "00000100", --  389 - 0x185  :    4 - 0x4
    "10000100", --  390 - 0x186  :  132 - 0x84
    "11111100", --  391 - 0x187  :  252 - 0xfc
    "01111111", --  392 - 0x188  :  127 - 0x7f -- Sprite 0x31
    "01111110", --  393 - 0x189  :  126 - 0x7e
    "11111100", --  394 - 0x18a  :  252 - 0xfc
    "00111000", --  395 - 0x18b  :   56 - 0x38
    "00111000", --  396 - 0x18c  :   56 - 0x38
    "00011100", --  397 - 0x18d  :   28 - 0x1c
    "10000100", --  398 - 0x18e  :  132 - 0x84
    "11000100", --  399 - 0x18f  :  196 - 0xc4
    "01111111", --  400 - 0x190  :  127 - 0x7f -- Sprite 0x32
    "01111110", --  401 - 0x191  :  126 - 0x7e
    "11111100", --  402 - 0x192  :  252 - 0xfc
    "00111000", --  403 - 0x193  :   56 - 0x38
    "00100100", --  404 - 0x194  :   36 - 0x24
    "00000100", --  405 - 0x195  :    4 - 0x4
    "10011100", --  406 - 0x196  :  156 - 0x9c
    "11111100", --  407 - 0x197  :  252 - 0xfc
    "00100011", --  408 - 0x198  :   35 - 0x23 -- Sprite 0x33
    "00100011", --  409 - 0x199  :   35 - 0x23
    "00100001", --  410 - 0x19a  :   33 - 0x21
    "00100000", --  411 - 0x19b  :   32 - 0x20
    "00010011", --  412 - 0x19c  :   19 - 0x13
    "00001101", --  413 - 0x19d  :   13 - 0xd
    "00000001", --  414 - 0x19e  :    1 - 0x1
    "00000001", --  415 - 0x19f  :    1 - 0x1
    "11111100", --  416 - 0x1a0  :  252 - 0xfc -- Sprite 0x34
    "11111100", --  417 - 0x1a1  :  252 - 0xfc
    "11111100", --  418 - 0x1a2  :  252 - 0xfc
    "11111100", --  419 - 0x1a3  :  252 - 0xfc
    "10100100", --  420 - 0x1a4  :  164 - 0xa4
    "00100100", --  421 - 0x1a5  :   36 - 0x24
    "00010010", --  422 - 0x1a6  :   18 - 0x12
    "11101110", --  423 - 0x1a7  :  238 - 0xee
    "00100011", --  424 - 0x1a8  :   35 - 0x23 -- Sprite 0x35
    "00100011", --  425 - 0x1a9  :   35 - 0x23
    "00100001", --  426 - 0x1aa  :   33 - 0x21
    "00100000", --  427 - 0x1ab  :   32 - 0x20
    "00010011", --  428 - 0x1ac  :   19 - 0x13
    "00001110", --  429 - 0x1ad  :   14 - 0xe
    "00000010", --  430 - 0x1ae  :    2 - 0x2
    "00000001", --  431 - 0x1af  :    1 - 0x1
    "11111100", --  432 - 0x1b0  :  252 - 0xfc -- Sprite 0x36
    "11111100", --  433 - 0x1b1  :  252 - 0xfc
    "11111100", --  434 - 0x1b2  :  252 - 0xfc
    "11111100", --  435 - 0x1b3  :  252 - 0xfc
    "10100110", --  436 - 0x1b4  :  166 - 0xa6
    "00110001", --  437 - 0x1b5  :   49 - 0x31
    "01001001", --  438 - 0x1b6  :   73 - 0x49
    "11000110", --  439 - 0x1b7  :  198 - 0xc6
    "11111100", --  440 - 0x1b8  :  252 - 0xfc -- Sprite 0x37
    "11111100", --  441 - 0x1b9  :  252 - 0xfc
    "11111100", --  442 - 0x1ba  :  252 - 0xfc
    "11111100", --  443 - 0x1bb  :  252 - 0xfc
    "10100100", --  444 - 0x1bc  :  164 - 0xa4
    "00100100", --  445 - 0x1bd  :   36 - 0x24
    "00010010", --  446 - 0x1be  :   18 - 0x12
    "11101110", --  447 - 0x1bf  :  238 - 0xee
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x40
    "00111110", --  513 - 0x201  :   62 - 0x3e
    "01111111", --  514 - 0x202  :  127 - 0x7f
    "01111111", --  515 - 0x203  :  127 - 0x7f
    "01111111", --  516 - 0x204  :  127 - 0x7f
    "01111111", --  517 - 0x205  :  127 - 0x7f
    "01111111", --  518 - 0x206  :  127 - 0x7f
    "00111110", --  519 - 0x207  :   62 - 0x3e
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Sprite 0x41
    "00111100", --  521 - 0x209  :   60 - 0x3c
    "00011100", --  522 - 0x20a  :   28 - 0x1c
    "00011100", --  523 - 0x20b  :   28 - 0x1c
    "00011100", --  524 - 0x20c  :   28 - 0x1c
    "00011100", --  525 - 0x20d  :   28 - 0x1c
    "00011100", --  526 - 0x20e  :   28 - 0x1c
    "00011100", --  527 - 0x20f  :   28 - 0x1c
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x42
    "01111100", --  529 - 0x211  :  124 - 0x7c
    "01111111", --  530 - 0x212  :  127 - 0x7f
    "01100111", --  531 - 0x213  :  103 - 0x67
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "01111110", --  533 - 0x215  :  126 - 0x7e
    "01111111", --  534 - 0x216  :  127 - 0x7f
    "01111111", --  535 - 0x217  :  127 - 0x7f
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Sprite 0x43
    "01111110", --  537 - 0x219  :  126 - 0x7e
    "01111111", --  538 - 0x21a  :  127 - 0x7f
    "01111111", --  539 - 0x21b  :  127 - 0x7f
    "00011111", --  540 - 0x21c  :   31 - 0x1f
    "01110111", --  541 - 0x21d  :  119 - 0x77
    "01111111", --  542 - 0x21e  :  127 - 0x7f
    "01111110", --  543 - 0x21f  :  126 - 0x7e
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x44
    "00001110", --  545 - 0x221  :   14 - 0xe
    "00011110", --  546 - 0x222  :   30 - 0x1e
    "00111110", --  547 - 0x223  :   62 - 0x3e
    "01111110", --  548 - 0x224  :  126 - 0x7e
    "01111111", --  549 - 0x225  :  127 - 0x7f
    "01111110", --  550 - 0x226  :  126 - 0x7e
    "00001100", --  551 - 0x227  :   12 - 0xc
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Sprite 0x45
    "01111111", --  553 - 0x229  :  127 - 0x7f
    "01111111", --  554 - 0x22a  :  127 - 0x7f
    "01111111", --  555 - 0x22b  :  127 - 0x7f
    "01111111", --  556 - 0x22c  :  127 - 0x7f
    "01110111", --  557 - 0x22d  :  119 - 0x77
    "01111111", --  558 - 0x22e  :  127 - 0x7f
    "01111110", --  559 - 0x22f  :  126 - 0x7e
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Sprite 0x46
    "00111110", --  561 - 0x231  :   62 - 0x3e
    "01111110", --  562 - 0x232  :  126 - 0x7e
    "01111111", --  563 - 0x233  :  127 - 0x7f
    "01111111", --  564 - 0x234  :  127 - 0x7f
    "01110111", --  565 - 0x235  :  119 - 0x77
    "01111111", --  566 - 0x236  :  127 - 0x7f
    "00111110", --  567 - 0x237  :   62 - 0x3e
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Sprite 0x47
    "01111110", --  569 - 0x239  :  126 - 0x7e
    "01111110", --  570 - 0x23a  :  126 - 0x7e
    "00011110", --  571 - 0x23b  :   30 - 0x1e
    "00011100", --  572 - 0x23c  :   28 - 0x1c
    "00111100", --  573 - 0x23d  :   60 - 0x3c
    "00111000", --  574 - 0x23e  :   56 - 0x38
    "00111000", --  575 - 0x23f  :   56 - 0x38
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x48
    "00111110", --  577 - 0x241  :   62 - 0x3e
    "01111111", --  578 - 0x242  :  127 - 0x7f
    "01111111", --  579 - 0x243  :  127 - 0x7f
    "01111111", --  580 - 0x244  :  127 - 0x7f
    "01111111", --  581 - 0x245  :  127 - 0x7f
    "01111111", --  582 - 0x246  :  127 - 0x7f
    "00111110", --  583 - 0x247  :   62 - 0x3e
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Sprite 0x49
    "00111110", --  585 - 0x249  :   62 - 0x3e
    "01111111", --  586 - 0x24a  :  127 - 0x7f
    "01110111", --  587 - 0x24b  :  119 - 0x77
    "01111111", --  588 - 0x24c  :  127 - 0x7f
    "01111111", --  589 - 0x24d  :  127 - 0x7f
    "00111111", --  590 - 0x24e  :   63 - 0x3f
    "00111110", --  591 - 0x24f  :   62 - 0x3e
    "11111111", --  592 - 0x250  :  255 - 0xff -- Sprite 0x4a
    "10011001", --  593 - 0x251  :  153 - 0x99
    "10011001", --  594 - 0x252  :  153 - 0x99
    "10011001", --  595 - 0x253  :  153 - 0x99
    "10011001", --  596 - 0x254  :  153 - 0x99
    "10011001", --  597 - 0x255  :  153 - 0x99
    "10011001", --  598 - 0x256  :  153 - 0x99
    "11111111", --  599 - 0x257  :  255 - 0xff
    "11110000", --  600 - 0x258  :  240 - 0xf0 -- Sprite 0x4b
    "10010000", --  601 - 0x259  :  144 - 0x90
    "10010000", --  602 - 0x25a  :  144 - 0x90
    "10010000", --  603 - 0x25b  :  144 - 0x90
    "10010000", --  604 - 0x25c  :  144 - 0x90
    "10010000", --  605 - 0x25d  :  144 - 0x90
    "10010000", --  606 - 0x25e  :  144 - 0x90
    "11110000", --  607 - 0x25f  :  240 - 0xf0
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x4c
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111111", --  614 - 0x266  :  255 - 0xff
    "11111111", --  615 - 0x267  :  255 - 0xff
    "11111111", --  616 - 0x268  :  255 - 0xff -- Sprite 0x4d
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11111111", --  620 - 0x26c  :  255 - 0xff
    "11111111", --  621 - 0x26d  :  255 - 0xff
    "11111111", --  622 - 0x26e  :  255 - 0xff
    "11111111", --  623 - 0x26f  :  255 - 0xff
    "11111111", --  624 - 0x270  :  255 - 0xff -- Sprite 0x4e
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11111111", --  626 - 0x272  :  255 - 0xff
    "11111111", --  627 - 0x273  :  255 - 0xff
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111111", --  629 - 0x275  :  255 - 0xff
    "11111111", --  630 - 0x276  :  255 - 0xff
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11111111", --  632 - 0x278  :  255 - 0xff -- Sprite 0x4f
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11111111", --  634 - 0x27a  :  255 - 0xff
    "11111111", --  635 - 0x27b  :  255 - 0xff
    "11111111", --  636 - 0x27c  :  255 - 0xff
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11111111", --  638 - 0x27e  :  255 - 0xff
    "11111111", --  639 - 0x27f  :  255 - 0xff
    "00010000", --  640 - 0x280  :   16 - 0x10 -- Sprite 0x50
    "00101000", --  641 - 0x281  :   40 - 0x28
    "11101110", --  642 - 0x282  :  238 - 0xee
    "10000010", --  643 - 0x283  :  130 - 0x82
    "01000100", --  644 - 0x284  :   68 - 0x44
    "01000100", --  645 - 0x285  :   68 - 0x44
    "10010010", --  646 - 0x286  :  146 - 0x92
    "11101110", --  647 - 0x287  :  238 - 0xee
    "00010000", --  648 - 0x288  :   16 - 0x10 -- Sprite 0x51
    "00101000", --  649 - 0x289  :   40 - 0x28
    "11101110", --  650 - 0x28a  :  238 - 0xee
    "10000010", --  651 - 0x28b  :  130 - 0x82
    "01000100", --  652 - 0x28c  :   68 - 0x44
    "01000100", --  653 - 0x28d  :   68 - 0x44
    "10010010", --  654 - 0x28e  :  146 - 0x92
    "11101110", --  655 - 0x28f  :  238 - 0xee
    "00010000", --  656 - 0x290  :   16 - 0x10 -- Sprite 0x52
    "00111000", --  657 - 0x291  :   56 - 0x38
    "11111110", --  658 - 0x292  :  254 - 0xfe
    "11111110", --  659 - 0x293  :  254 - 0xfe
    "01111100", --  660 - 0x294  :  124 - 0x7c
    "01111100", --  661 - 0x295  :  124 - 0x7c
    "11111110", --  662 - 0x296  :  254 - 0xfe
    "11101110", --  663 - 0x297  :  238 - 0xee
    "11111111", --  664 - 0x298  :  255 - 0xff -- Sprite 0x53
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111111", --  668 - 0x29c  :  255 - 0xff
    "11111111", --  669 - 0x29d  :  255 - 0xff
    "11111111", --  670 - 0x29e  :  255 - 0xff
    "11111111", --  671 - 0x29f  :  255 - 0xff
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Sprite 0x55
    "11111111", --  681 - 0x2a9  :  255 - 0xff
    "11111111", --  682 - 0x2aa  :  255 - 0xff
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11111111", --  684 - 0x2ac  :  255 - 0xff
    "11111111", --  685 - 0x2ad  :  255 - 0xff
    "11111111", --  686 - 0x2ae  :  255 - 0xff
    "11111111", --  687 - 0x2af  :  255 - 0xff
    "00101010", --  688 - 0x2b0  :   42 - 0x2a -- Sprite 0x56
    "01000101", --  689 - 0x2b1  :   69 - 0x45
    "00001000", --  690 - 0x2b2  :    8 - 0x8
    "00010101", --  691 - 0x2b3  :   21 - 0x15
    "00100000", --  692 - 0x2b4  :   32 - 0x20
    "01000101", --  693 - 0x2b5  :   69 - 0x45
    "10101000", --  694 - 0x2b6  :  168 - 0xa8
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00001000", --  696 - 0x2b8  :    8 - 0x8 -- Sprite 0x57
    "01010101", --  697 - 0x2b9  :   85 - 0x55
    "10100000", --  698 - 0x2ba  :  160 - 0xa0
    "00010000", --  699 - 0x2bb  :   16 - 0x10
    "10000000", --  700 - 0x2bc  :  128 - 0x80
    "00010100", --  701 - 0x2bd  :   20 - 0x14
    "00100010", --  702 - 0x2be  :   34 - 0x22
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Sprite 0x58
    "11010101", --  705 - 0x2c1  :  213 - 0xd5
    "10100000", --  706 - 0x2c2  :  160 - 0xa0
    "11010000", --  707 - 0x2c3  :  208 - 0xd0
    "10001111", --  708 - 0x2c4  :  143 - 0x8f
    "11001000", --  709 - 0x2c5  :  200 - 0xc8
    "10001000", --  710 - 0x2c6  :  136 - 0x88
    "11001000", --  711 - 0x2c7  :  200 - 0xc8
    "10001000", --  712 - 0x2c8  :  136 - 0x88 -- Sprite 0x59
    "11001000", --  713 - 0x2c9  :  200 - 0xc8
    "10001000", --  714 - 0x2ca  :  136 - 0x88
    "11001111", --  715 - 0x2cb  :  207 - 0xcf
    "10010000", --  716 - 0x2cc  :  144 - 0x90
    "11100000", --  717 - 0x2cd  :  224 - 0xe0
    "11101010", --  718 - 0x2ce  :  234 - 0xea
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Sprite 0x5a
    "01011011", --  721 - 0x2d1  :   91 - 0x5b
    "00000111", --  722 - 0x2d2  :    7 - 0x7
    "00001001", --  723 - 0x2d3  :    9 - 0x9
    "11110011", --  724 - 0x2d4  :  243 - 0xf3
    "00010001", --  725 - 0x2d5  :   17 - 0x11
    "00010011", --  726 - 0x2d6  :   19 - 0x13
    "00010001", --  727 - 0x2d7  :   17 - 0x11
    "00010011", --  728 - 0x2d8  :   19 - 0x13 -- Sprite 0x5b
    "00010001", --  729 - 0x2d9  :   17 - 0x11
    "00010011", --  730 - 0x2da  :   19 - 0x13
    "11110001", --  731 - 0x2db  :  241 - 0xf1
    "00001011", --  732 - 0x2dc  :   11 - 0xb
    "00000101", --  733 - 0x2dd  :    5 - 0x5
    "10101011", --  734 - 0x2de  :  171 - 0xab
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00011100", --  736 - 0x2e0  :   28 - 0x1c -- Sprite 0x5c
    "00100010", --  737 - 0x2e1  :   34 - 0x22
    "01000001", --  738 - 0x2e2  :   65 - 0x41
    "01000001", --  739 - 0x2e3  :   65 - 0x41
    "01000001", --  740 - 0x2e4  :   65 - 0x41
    "00100010", --  741 - 0x2e5  :   34 - 0x22
    "00100010", --  742 - 0x2e6  :   34 - 0x22
    "00011100", --  743 - 0x2e7  :   28 - 0x1c
    "00001000", --  744 - 0x2e8  :    8 - 0x8 -- Sprite 0x5d
    "00010000", --  745 - 0x2e9  :   16 - 0x10
    "00010000", --  746 - 0x2ea  :   16 - 0x10
    "00001000", --  747 - 0x2eb  :    8 - 0x8
    "00000100", --  748 - 0x2ec  :    4 - 0x4
    "00000100", --  749 - 0x2ed  :    4 - 0x4
    "00001000", --  750 - 0x2ee  :    8 - 0x8
    "00010000", --  751 - 0x2ef  :   16 - 0x10
    "00110110", --  752 - 0x2f0  :   54 - 0x36 -- Sprite 0x5e
    "01101011", --  753 - 0x2f1  :  107 - 0x6b
    "01001001", --  754 - 0x2f2  :   73 - 0x49
    "01000001", --  755 - 0x2f3  :   65 - 0x41
    "01000001", --  756 - 0x2f4  :   65 - 0x41
    "00100010", --  757 - 0x2f5  :   34 - 0x22
    "00010100", --  758 - 0x2f6  :   20 - 0x14
    "00001000", --  759 - 0x2f7  :    8 - 0x8
    "00111110", --  760 - 0x2f8  :   62 - 0x3e -- Sprite 0x5f
    "01101011", --  761 - 0x2f9  :  107 - 0x6b
    "00100010", --  762 - 0x2fa  :   34 - 0x22
    "01100011", --  763 - 0x2fb  :   99 - 0x63
    "00100010", --  764 - 0x2fc  :   34 - 0x22
    "01100011", --  765 - 0x2fd  :   99 - 0x63
    "00100010", --  766 - 0x2fe  :   34 - 0x22
    "01111111", --  767 - 0x2ff  :  127 - 0x7f
    "11111111", --  768 - 0x300  :  255 - 0xff -- Sprite 0x60
    "11111111", --  769 - 0x301  :  255 - 0xff
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11010101", --  772 - 0x304  :  213 - 0xd5
    "10101010", --  773 - 0x305  :  170 - 0xaa
    "11010101", --  774 - 0x306  :  213 - 0xd5
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff -- Sprite 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "01010101", --  780 - 0x30c  :   85 - 0x55
    "10101010", --  781 - 0x30d  :  170 - 0xaa
    "01010101", --  782 - 0x30e  :   85 - 0x55
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff -- Sprite 0x62
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "01010101", --  788 - 0x314  :   85 - 0x55
    "10101011", --  789 - 0x315  :  171 - 0xab
    "01010101", --  790 - 0x316  :   85 - 0x55
    "11111111", --  791 - 0x317  :  255 - 0xff
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Sprite 0x63
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000001", --  800 - 0x320  :    1 - 0x1 -- Sprite 0x64
    "00000001", --  801 - 0x321  :    1 - 0x1
    "00000011", --  802 - 0x322  :    3 - 0x3
    "00000011", --  803 - 0x323  :    3 - 0x3
    "00000110", --  804 - 0x324  :    6 - 0x6
    "00000110", --  805 - 0x325  :    6 - 0x6
    "00001100", --  806 - 0x326  :   12 - 0xc
    "00001100", --  807 - 0x327  :   12 - 0xc
    "00011000", --  808 - 0x328  :   24 - 0x18 -- Sprite 0x65
    "00011000", --  809 - 0x329  :   24 - 0x18
    "00110000", --  810 - 0x32a  :   48 - 0x30
    "00110000", --  811 - 0x32b  :   48 - 0x30
    "01100000", --  812 - 0x32c  :   96 - 0x60
    "01100000", --  813 - 0x32d  :   96 - 0x60
    "11101010", --  814 - 0x32e  :  234 - 0xea
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "10000000", --  816 - 0x330  :  128 - 0x80 -- Sprite 0x66
    "10000000", --  817 - 0x331  :  128 - 0x80
    "11000000", --  818 - 0x332  :  192 - 0xc0
    "01000000", --  819 - 0x333  :   64 - 0x40
    "10100000", --  820 - 0x334  :  160 - 0xa0
    "01100000", --  821 - 0x335  :   96 - 0x60
    "00110000", --  822 - 0x336  :   48 - 0x30
    "00010000", --  823 - 0x337  :   16 - 0x10
    "00101000", --  824 - 0x338  :   40 - 0x28 -- Sprite 0x67
    "00011000", --  825 - 0x339  :   24 - 0x18
    "00001100", --  826 - 0x33a  :   12 - 0xc
    "00010100", --  827 - 0x33b  :   20 - 0x14
    "00001010", --  828 - 0x33c  :   10 - 0xa
    "00000110", --  829 - 0x33d  :    6 - 0x6
    "10101011", --  830 - 0x33e  :  171 - 0xab
    "11111111", --  831 - 0x33f  :  255 - 0xff
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- Sprite 0x6f
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Sprite 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Sprite 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Sprite 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Sprite 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000011", -- 1024 - 0x400  :    3 - 0x3 -- Sprite 0x80
    "00001111", -- 1025 - 0x401  :   15 - 0xf
    "00011100", -- 1026 - 0x402  :   28 - 0x1c
    "00110000", -- 1027 - 0x403  :   48 - 0x30
    "00100000", -- 1028 - 0x404  :   32 - 0x20
    "01000000", -- 1029 - 0x405  :   64 - 0x40
    "01000000", -- 1030 - 0x406  :   64 - 0x40
    "01111111", -- 1031 - 0x407  :  127 - 0x7f
    "00000001", -- 1032 - 0x408  :    1 - 0x1 -- Sprite 0x81
    "00000001", -- 1033 - 0x409  :    1 - 0x1
    "00000001", -- 1034 - 0x40a  :    1 - 0x1
    "00000001", -- 1035 - 0x40b  :    1 - 0x1
    "00000001", -- 1036 - 0x40c  :    1 - 0x1
    "00000001", -- 1037 - 0x40d  :    1 - 0x1
    "00000011", -- 1038 - 0x40e  :    3 - 0x3
    "00000011", -- 1039 - 0x40f  :    3 - 0x3
    "11000000", -- 1040 - 0x410  :  192 - 0xc0 -- Sprite 0x82
    "11110000", -- 1041 - 0x411  :  240 - 0xf0
    "00111000", -- 1042 - 0x412  :   56 - 0x38
    "00001110", -- 1043 - 0x413  :   14 - 0xe
    "00011110", -- 1044 - 0x414  :   30 - 0x1e
    "00011110", -- 1045 - 0x415  :   30 - 0x1e
    "00000010", -- 1046 - 0x416  :    2 - 0x2
    "11111110", -- 1047 - 0x417  :  254 - 0xfe
    "10000000", -- 1048 - 0x418  :  128 - 0x80 -- Sprite 0x83
    "10000000", -- 1049 - 0x419  :  128 - 0x80
    "10000000", -- 1050 - 0x41a  :  128 - 0x80
    "10000000", -- 1051 - 0x41b  :  128 - 0x80
    "10000000", -- 1052 - 0x41c  :  128 - 0x80
    "11100000", -- 1053 - 0x41d  :  224 - 0xe0
    "00010000", -- 1054 - 0x41e  :   16 - 0x10
    "11110000", -- 1055 - 0x41f  :  240 - 0xf0
    "00000011", -- 1056 - 0x420  :    3 - 0x3 -- Sprite 0x84
    "00001111", -- 1057 - 0x421  :   15 - 0xf
    "00011100", -- 1058 - 0x422  :   28 - 0x1c
    "00110000", -- 1059 - 0x423  :   48 - 0x30
    "00100000", -- 1060 - 0x424  :   32 - 0x20
    "01000000", -- 1061 - 0x425  :   64 - 0x40
    "01000000", -- 1062 - 0x426  :   64 - 0x40
    "01111111", -- 1063 - 0x427  :  127 - 0x7f
    "00000011", -- 1064 - 0x428  :    3 - 0x3 -- Sprite 0x85
    "00000110", -- 1065 - 0x429  :    6 - 0x6
    "00000110", -- 1066 - 0x42a  :    6 - 0x6
    "00011100", -- 1067 - 0x42b  :   28 - 0x1c
    "00011000", -- 1068 - 0x42c  :   24 - 0x18
    "00110110", -- 1069 - 0x42d  :   54 - 0x36
    "00110001", -- 1070 - 0x42e  :   49 - 0x31
    "00001111", -- 1071 - 0x42f  :   15 - 0xf
    "11000000", -- 1072 - 0x430  :  192 - 0xc0 -- Sprite 0x86
    "11110000", -- 1073 - 0x431  :  240 - 0xf0
    "00111000", -- 1074 - 0x432  :   56 - 0x38
    "00001110", -- 1075 - 0x433  :   14 - 0xe
    "00011110", -- 1076 - 0x434  :   30 - 0x1e
    "00011110", -- 1077 - 0x435  :   30 - 0x1e
    "00000010", -- 1078 - 0x436  :    2 - 0x2
    "11111110", -- 1079 - 0x437  :  254 - 0xfe
    "11000000", -- 1080 - 0x438  :  192 - 0xc0 -- Sprite 0x87
    "01100000", -- 1081 - 0x439  :   96 - 0x60
    "01100000", -- 1082 - 0x43a  :   96 - 0x60
    "00110000", -- 1083 - 0x43b  :   48 - 0x30
    "00111110", -- 1084 - 0x43c  :   62 - 0x3e
    "00011001", -- 1085 - 0x43d  :   25 - 0x19
    "00110011", -- 1086 - 0x43e  :   51 - 0x33
    "00111100", -- 1087 - 0x43f  :   60 - 0x3c
    "00000011", -- 1088 - 0x440  :    3 - 0x3 -- Sprite 0x88
    "00000111", -- 1089 - 0x441  :    7 - 0x7
    "00000111", -- 1090 - 0x442  :    7 - 0x7
    "00001011", -- 1091 - 0x443  :   11 - 0xb
    "00010000", -- 1092 - 0x444  :   16 - 0x10
    "01100000", -- 1093 - 0x445  :   96 - 0x60
    "11110000", -- 1094 - 0x446  :  240 - 0xf0
    "11110000", -- 1095 - 0x447  :  240 - 0xf0
    "11110000", -- 1096 - 0x448  :  240 - 0xf0 -- Sprite 0x89
    "11110000", -- 1097 - 0x449  :  240 - 0xf0
    "01100000", -- 1098 - 0x44a  :   96 - 0x60
    "00010000", -- 1099 - 0x44b  :   16 - 0x10
    "00001011", -- 1100 - 0x44c  :   11 - 0xb
    "00000111", -- 1101 - 0x44d  :    7 - 0x7
    "00000111", -- 1102 - 0x44e  :    7 - 0x7
    "00000011", -- 1103 - 0x44f  :    3 - 0x3
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x8a
    "00011100", -- 1105 - 0x451  :   28 - 0x1c
    "00111111", -- 1106 - 0x452  :   63 - 0x3f
    "01111000", -- 1107 - 0x453  :  120 - 0x78
    "01110000", -- 1108 - 0x454  :  112 - 0x70
    "01100000", -- 1109 - 0x455  :   96 - 0x60
    "00100000", -- 1110 - 0x456  :   32 - 0x20
    "00100000", -- 1111 - 0x457  :   32 - 0x20
    "00100000", -- 1112 - 0x458  :   32 - 0x20 -- Sprite 0x8b
    "00100000", -- 1113 - 0x459  :   32 - 0x20
    "01100000", -- 1114 - 0x45a  :   96 - 0x60
    "01110000", -- 1115 - 0x45b  :  112 - 0x70
    "01111000", -- 1116 - 0x45c  :  120 - 0x78
    "00111111", -- 1117 - 0x45d  :   63 - 0x3f
    "00011100", -- 1118 - 0x45e  :   28 - 0x1c
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000011", -- 1120 - 0x460  :    3 - 0x3 -- Sprite 0x8c
    "00001100", -- 1121 - 0x461  :   12 - 0xc
    "00011110", -- 1122 - 0x462  :   30 - 0x1e
    "00100110", -- 1123 - 0x463  :   38 - 0x26
    "01000110", -- 1124 - 0x464  :   70 - 0x46
    "01100100", -- 1125 - 0x465  :  100 - 0x64
    "01110000", -- 1126 - 0x466  :  112 - 0x70
    "11110000", -- 1127 - 0x467  :  240 - 0xf0
    "10101010", -- 1128 - 0x468  :  170 - 0xaa -- Sprite 0x8d
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "01111111", -- 1130 - 0x46a  :  127 - 0x7f
    "00111001", -- 1131 - 0x46b  :   57 - 0x39
    "00011001", -- 1132 - 0x46c  :   25 - 0x19
    "00001011", -- 1133 - 0x46d  :   11 - 0xb
    "00001000", -- 1134 - 0x46e  :    8 - 0x8
    "00000111", -- 1135 - 0x46f  :    7 - 0x7
    "11000000", -- 1136 - 0x470  :  192 - 0xc0 -- Sprite 0x8e
    "00110000", -- 1137 - 0x471  :   48 - 0x30
    "00001000", -- 1138 - 0x472  :    8 - 0x8
    "01000100", -- 1139 - 0x473  :   68 - 0x44
    "01100010", -- 1140 - 0x474  :   98 - 0x62
    "01100010", -- 1141 - 0x475  :   98 - 0x62
    "00000001", -- 1142 - 0x476  :    1 - 0x1
    "00111111", -- 1143 - 0x477  :   63 - 0x3f
    "10001011", -- 1144 - 0x478  :  139 - 0x8b -- Sprite 0x8f
    "11000001", -- 1145 - 0x479  :  193 - 0xc1
    "11111110", -- 1146 - 0x47a  :  254 - 0xfe
    "11111100", -- 1147 - 0x47b  :  252 - 0xfc
    "11110000", -- 1148 - 0x47c  :  240 - 0xf0
    "11110000", -- 1149 - 0x47d  :  240 - 0xf0
    "11111000", -- 1150 - 0x47e  :  248 - 0xf8
    "11110000", -- 1151 - 0x47f  :  240 - 0xf0
    "00000011", -- 1152 - 0x480  :    3 - 0x3 -- Sprite 0x90
    "00001110", -- 1153 - 0x481  :   14 - 0xe
    "00010110", -- 1154 - 0x482  :   22 - 0x16
    "00100110", -- 1155 - 0x483  :   38 - 0x26
    "01100011", -- 1156 - 0x484  :   99 - 0x63
    "01110010", -- 1157 - 0x485  :  114 - 0x72
    "01110000", -- 1158 - 0x486  :  112 - 0x70
    "11010000", -- 1159 - 0x487  :  208 - 0xd0
    "10101010", -- 1160 - 0x488  :  170 - 0xaa -- Sprite 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "01111111", -- 1162 - 0x48a  :  127 - 0x7f
    "00111100", -- 1163 - 0x48b  :   60 - 0x3c
    "00011100", -- 1164 - 0x48c  :   28 - 0x1c
    "00000100", -- 1165 - 0x48d  :    4 - 0x4
    "00000010", -- 1166 - 0x48e  :    2 - 0x2
    "00000001", -- 1167 - 0x48f  :    1 - 0x1
    "11000000", -- 1168 - 0x490  :  192 - 0xc0 -- Sprite 0x92
    "00110000", -- 1169 - 0x491  :   48 - 0x30
    "00001000", -- 1170 - 0x492  :    8 - 0x8
    "00100100", -- 1171 - 0x493  :   36 - 0x24
    "00110010", -- 1172 - 0x494  :   50 - 0x32
    "00110010", -- 1173 - 0x495  :   50 - 0x32
    "00000001", -- 1174 - 0x496  :    1 - 0x1
    "00011111", -- 1175 - 0x497  :   31 - 0x1f
    "10001011", -- 1176 - 0x498  :  139 - 0x8b -- Sprite 0x93
    "11000001", -- 1177 - 0x499  :  193 - 0xc1
    "11111110", -- 1178 - 0x49a  :  254 - 0xfe
    "11111100", -- 1179 - 0x49b  :  252 - 0xfc
    "11110000", -- 1180 - 0x49c  :  240 - 0xf0
    "11000000", -- 1181 - 0x49d  :  192 - 0xc0
    "00100000", -- 1182 - 0x49e  :   32 - 0x20
    "11100000", -- 1183 - 0x49f  :  224 - 0xe0
    "00000011", -- 1184 - 0x4a0  :    3 - 0x3 -- Sprite 0x94
    "00001111", -- 1185 - 0x4a1  :   15 - 0xf
    "00010011", -- 1186 - 0x4a2  :   19 - 0x13
    "00110001", -- 1187 - 0x4a3  :   49 - 0x31
    "01111001", -- 1188 - 0x4a4  :  121 - 0x79
    "01011001", -- 1189 - 0x4a5  :   89 - 0x59
    "01001000", -- 1190 - 0x4a6  :   72 - 0x48
    "11001100", -- 1191 - 0x4a7  :  204 - 0xcc
    "10010101", -- 1192 - 0x4a8  :  149 - 0x95 -- Sprite 0x95
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "01111111", -- 1194 - 0x4aa  :  127 - 0x7f
    "00111110", -- 1195 - 0x4ab  :   62 - 0x3e
    "00011111", -- 1196 - 0x4ac  :   31 - 0x1f
    "00001111", -- 1197 - 0x4ad  :   15 - 0xf
    "00001111", -- 1198 - 0x4ae  :   15 - 0xf
    "00000111", -- 1199 - 0x4af  :    7 - 0x7
    "11000000", -- 1200 - 0x4b0  :  192 - 0xc0 -- Sprite 0x96
    "00110000", -- 1201 - 0x4b1  :   48 - 0x30
    "00001000", -- 1202 - 0x4b2  :    8 - 0x8
    "10010100", -- 1203 - 0x4b3  :  148 - 0x94
    "10011010", -- 1204 - 0x4b4  :  154 - 0x9a
    "00011010", -- 1205 - 0x4b5  :   26 - 0x1a
    "00000001", -- 1206 - 0x4b6  :    1 - 0x1
    "00001111", -- 1207 - 0x4b7  :   15 - 0xf
    "01000101", -- 1208 - 0x4b8  :   69 - 0x45 -- Sprite 0x97
    "11100001", -- 1209 - 0x4b9  :  225 - 0xe1
    "11111110", -- 1210 - 0x4ba  :  254 - 0xfe
    "01111100", -- 1211 - 0x4bb  :  124 - 0x7c
    "00110000", -- 1212 - 0x4bc  :   48 - 0x30
    "00110000", -- 1213 - 0x4bd  :   48 - 0x30
    "10001000", -- 1214 - 0x4be  :  136 - 0x88
    "01111000", -- 1215 - 0x4bf  :  120 - 0x78
    "00000001", -- 1216 - 0x4c0  :    1 - 0x1 -- Sprite 0x98
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000001", -- 1220 - 0x4c4  :    1 - 0x1
    "00000001", -- 1221 - 0x4c5  :    1 - 0x1
    "00000010", -- 1222 - 0x4c6  :    2 - 0x2
    "00000110", -- 1223 - 0x4c7  :    6 - 0x6
    "01111000", -- 1224 - 0x4c8  :  120 - 0x78 -- Sprite 0x99
    "00101010", -- 1225 - 0x4c9  :   42 - 0x2a
    "01010100", -- 1226 - 0x4ca  :   84 - 0x54
    "00101001", -- 1227 - 0x4cb  :   41 - 0x29
    "00101111", -- 1228 - 0x4cc  :   47 - 0x2f
    "00110111", -- 1229 - 0x4cd  :   55 - 0x37
    "00000011", -- 1230 - 0x4ce  :    3 - 0x3
    "00000111", -- 1231 - 0x4cf  :    7 - 0x7
    "10110000", -- 1232 - 0x4d0  :  176 - 0xb0 -- Sprite 0x9a
    "11101000", -- 1233 - 0x4d1  :  232 - 0xe8
    "10001100", -- 1234 - 0x4d2  :  140 - 0x8c
    "10011110", -- 1235 - 0x4d3  :  158 - 0x9e
    "00011111", -- 1236 - 0x4d4  :   31 - 0x1f
    "00001111", -- 1237 - 0x4d5  :   15 - 0xf
    "10010110", -- 1238 - 0x4d6  :  150 - 0x96
    "00011100", -- 1239 - 0x4d7  :   28 - 0x1c
    "00001100", -- 1240 - 0x4d8  :   12 - 0xc -- Sprite 0x9b
    "00111000", -- 1241 - 0x4d9  :   56 - 0x38
    "11101000", -- 1242 - 0x4da  :  232 - 0xe8
    "11010000", -- 1243 - 0x4db  :  208 - 0xd0
    "11100000", -- 1244 - 0x4dc  :  224 - 0xe0
    "10000000", -- 1245 - 0x4dd  :  128 - 0x80
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "10000000", -- 1247 - 0x4df  :  128 - 0x80
    "00000001", -- 1248 - 0x4e0  :    1 - 0x1 -- Sprite 0x9c
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000001", -- 1252 - 0x4e4  :    1 - 0x1
    "00000001", -- 1253 - 0x4e5  :    1 - 0x1
    "00000010", -- 1254 - 0x4e6  :    2 - 0x2
    "00000110", -- 1255 - 0x4e7  :    6 - 0x6
    "01111000", -- 1256 - 0x4e8  :  120 - 0x78 -- Sprite 0x9d
    "00101010", -- 1257 - 0x4e9  :   42 - 0x2a
    "01010100", -- 1258 - 0x4ea  :   84 - 0x54
    "00101001", -- 1259 - 0x4eb  :   41 - 0x29
    "00101111", -- 1260 - 0x4ec  :   47 - 0x2f
    "00111100", -- 1261 - 0x4ed  :   60 - 0x3c
    "00011110", -- 1262 - 0x4ee  :   30 - 0x1e
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "10110000", -- 1264 - 0x4f0  :  176 - 0xb0 -- Sprite 0x9e
    "11101000", -- 1265 - 0x4f1  :  232 - 0xe8
    "10001100", -- 1266 - 0x4f2  :  140 - 0x8c
    "10011110", -- 1267 - 0x4f3  :  158 - 0x9e
    "00011111", -- 1268 - 0x4f4  :   31 - 0x1f
    "00001111", -- 1269 - 0x4f5  :   15 - 0xf
    "10010110", -- 1270 - 0x4f6  :  150 - 0x96
    "00011100", -- 1271 - 0x4f7  :   28 - 0x1c
    "00001100", -- 1272 - 0x4f8  :   12 - 0xc -- Sprite 0x9f
    "00111000", -- 1273 - 0x4f9  :   56 - 0x38
    "11101000", -- 1274 - 0x4fa  :  232 - 0xe8
    "11110000", -- 1275 - 0x4fb  :  240 - 0xf0
    "11000000", -- 1276 - 0x4fc  :  192 - 0xc0
    "01110000", -- 1277 - 0x4fd  :  112 - 0x70
    "11000000", -- 1278 - 0x4fe  :  192 - 0xc0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000011", -- 1280 - 0x500  :    3 - 0x3 -- Sprite 0xa0
    "00001111", -- 1281 - 0x501  :   15 - 0xf
    "00011100", -- 1282 - 0x502  :   28 - 0x1c
    "00110000", -- 1283 - 0x503  :   48 - 0x30
    "01100000", -- 1284 - 0x504  :   96 - 0x60
    "01100000", -- 1285 - 0x505  :   96 - 0x60
    "11000000", -- 1286 - 0x506  :  192 - 0xc0
    "11000000", -- 1287 - 0x507  :  192 - 0xc0
    "11000000", -- 1288 - 0x508  :  192 - 0xc0 -- Sprite 0xa1
    "11000000", -- 1289 - 0x509  :  192 - 0xc0
    "01100000", -- 1290 - 0x50a  :   96 - 0x60
    "01100000", -- 1291 - 0x50b  :   96 - 0x60
    "00110000", -- 1292 - 0x50c  :   48 - 0x30
    "00011010", -- 1293 - 0x50d  :   26 - 0x1a
    "00001101", -- 1294 - 0x50e  :   13 - 0xd
    "00000011", -- 1295 - 0x50f  :    3 - 0x3
    "11000000", -- 1296 - 0x510  :  192 - 0xc0 -- Sprite 0xa2
    "11110000", -- 1297 - 0x511  :  240 - 0xf0
    "00111000", -- 1298 - 0x512  :   56 - 0x38
    "00001100", -- 1299 - 0x513  :   12 - 0xc
    "00000110", -- 1300 - 0x514  :    6 - 0x6
    "00000010", -- 1301 - 0x515  :    2 - 0x2
    "00000101", -- 1302 - 0x516  :    5 - 0x5
    "00000011", -- 1303 - 0x517  :    3 - 0x3
    "00000101", -- 1304 - 0x518  :    5 - 0x5 -- Sprite 0xa3
    "00001011", -- 1305 - 0x519  :   11 - 0xb
    "00010110", -- 1306 - 0x51a  :   22 - 0x16
    "00101010", -- 1307 - 0x51b  :   42 - 0x2a
    "01010100", -- 1308 - 0x51c  :   84 - 0x54
    "10101000", -- 1309 - 0x51d  :  168 - 0xa8
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "11000000", -- 1311 - 0x51f  :  192 - 0xc0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0xa4
    "00001111", -- 1313 - 0x521  :   15 - 0xf
    "00011111", -- 1314 - 0x522  :   31 - 0x1f
    "00110001", -- 1315 - 0x523  :   49 - 0x31
    "00111111", -- 1316 - 0x524  :   63 - 0x3f
    "01111111", -- 1317 - 0x525  :  127 - 0x7f
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11011111", -- 1319 - 0x527  :  223 - 0xdf
    "11000000", -- 1320 - 0x528  :  192 - 0xc0 -- Sprite 0xa5
    "11000111", -- 1321 - 0x529  :  199 - 0xc7
    "01101111", -- 1322 - 0x52a  :  111 - 0x6f
    "01100111", -- 1323 - 0x52b  :  103 - 0x67
    "01100011", -- 1324 - 0x52c  :   99 - 0x63
    "00110000", -- 1325 - 0x52d  :   48 - 0x30
    "00011000", -- 1326 - 0x52e  :   24 - 0x18
    "00000111", -- 1327 - 0x52f  :    7 - 0x7
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "11110000", -- 1329 - 0x531  :  240 - 0xf0
    "11111000", -- 1330 - 0x532  :  248 - 0xf8
    "10001100", -- 1331 - 0x533  :  140 - 0x8c
    "11111100", -- 1332 - 0x534  :  252 - 0xfc
    "11111110", -- 1333 - 0x535  :  254 - 0xfe
    "11111101", -- 1334 - 0x536  :  253 - 0xfd
    "11111001", -- 1335 - 0x537  :  249 - 0xf9
    "00000011", -- 1336 - 0x538  :    3 - 0x3 -- Sprite 0xa7
    "11100101", -- 1337 - 0x539  :  229 - 0xe5
    "11110010", -- 1338 - 0x53a  :  242 - 0xf2
    "11100110", -- 1339 - 0x53b  :  230 - 0xe6
    "11001010", -- 1340 - 0x53c  :  202 - 0xca
    "00010100", -- 1341 - 0x53d  :   20 - 0x14
    "00111000", -- 1342 - 0x53e  :   56 - 0x38
    "11100000", -- 1343 - 0x53f  :  224 - 0xe0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0xa8
    "00001111", -- 1345 - 0x541  :   15 - 0xf
    "00011111", -- 1346 - 0x542  :   31 - 0x1f
    "00110001", -- 1347 - 0x543  :   49 - 0x31
    "00111111", -- 1348 - 0x544  :   63 - 0x3f
    "01111111", -- 1349 - 0x545  :  127 - 0x7f
    "11111111", -- 1350 - 0x546  :  255 - 0xff
    "11011111", -- 1351 - 0x547  :  223 - 0xdf
    "11000000", -- 1352 - 0x548  :  192 - 0xc0 -- Sprite 0xa9
    "11000011", -- 1353 - 0x549  :  195 - 0xc3
    "11000111", -- 1354 - 0x54a  :  199 - 0xc7
    "11001111", -- 1355 - 0x54b  :  207 - 0xcf
    "11000111", -- 1356 - 0x54c  :  199 - 0xc7
    "11000000", -- 1357 - 0x54d  :  192 - 0xc0
    "11100000", -- 1358 - 0x54e  :  224 - 0xe0
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "11110000", -- 1361 - 0x551  :  240 - 0xf0
    "11111000", -- 1362 - 0x552  :  248 - 0xf8
    "10001100", -- 1363 - 0x553  :  140 - 0x8c
    "11111100", -- 1364 - 0x554  :  252 - 0xfc
    "11111110", -- 1365 - 0x555  :  254 - 0xfe
    "11111101", -- 1366 - 0x556  :  253 - 0xfd
    "11111001", -- 1367 - 0x557  :  249 - 0xf9
    "00000011", -- 1368 - 0x558  :    3 - 0x3 -- Sprite 0xab
    "11000101", -- 1369 - 0x559  :  197 - 0xc5
    "11100011", -- 1370 - 0x55a  :  227 - 0xe3
    "11110101", -- 1371 - 0x55b  :  245 - 0xf5
    "11100011", -- 1372 - 0x55c  :  227 - 0xe3
    "00000101", -- 1373 - 0x55d  :    5 - 0x5
    "00001011", -- 1374 - 0x55e  :   11 - 0xb
    "11111111", -- 1375 - 0x55f  :  255 - 0xff
    "10000011", -- 1376 - 0x560  :  131 - 0x83 -- Sprite 0xac
    "10001100", -- 1377 - 0x561  :  140 - 0x8c
    "10010000", -- 1378 - 0x562  :  144 - 0x90
    "10010000", -- 1379 - 0x563  :  144 - 0x90
    "11100000", -- 1380 - 0x564  :  224 - 0xe0
    "10100000", -- 1381 - 0x565  :  160 - 0xa0
    "10101111", -- 1382 - 0x566  :  175 - 0xaf
    "01101111", -- 1383 - 0x567  :  111 - 0x6f
    "11111011", -- 1384 - 0x568  :  251 - 0xfb -- Sprite 0xad
    "00000101", -- 1385 - 0x569  :    5 - 0x5
    "00000101", -- 1386 - 0x56a  :    5 - 0x5
    "00000101", -- 1387 - 0x56b  :    5 - 0x5
    "01000101", -- 1388 - 0x56c  :   69 - 0x45
    "01100101", -- 1389 - 0x56d  :  101 - 0x65
    "11110101", -- 1390 - 0x56e  :  245 - 0xf5
    "11111101", -- 1391 - 0x56f  :  253 - 0xfd
    "10000011", -- 1392 - 0x570  :  131 - 0x83 -- Sprite 0xae
    "10001100", -- 1393 - 0x571  :  140 - 0x8c
    "10010000", -- 1394 - 0x572  :  144 - 0x90
    "10010000", -- 1395 - 0x573  :  144 - 0x90
    "11100000", -- 1396 - 0x574  :  224 - 0xe0
    "10100000", -- 1397 - 0x575  :  160 - 0xa0
    "10101111", -- 1398 - 0x576  :  175 - 0xaf
    "01101111", -- 1399 - 0x577  :  111 - 0x6f
    "11111011", -- 1400 - 0x578  :  251 - 0xfb -- Sprite 0xaf
    "00000101", -- 1401 - 0x579  :    5 - 0x5
    "00000101", -- 1402 - 0x57a  :    5 - 0x5
    "00000101", -- 1403 - 0x57b  :    5 - 0x5
    "11000101", -- 1404 - 0x57c  :  197 - 0xc5
    "11100101", -- 1405 - 0x57d  :  229 - 0xe5
    "11110101", -- 1406 - 0x57e  :  245 - 0xf5
    "11111101", -- 1407 - 0x57f  :  253 - 0xfd
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00000011", -- 1409 - 0x581  :    3 - 0x3
    "00001111", -- 1410 - 0x582  :   15 - 0xf
    "00111111", -- 1411 - 0x583  :   63 - 0x3f
    "01111111", -- 1412 - 0x584  :  127 - 0x7f
    "01111111", -- 1413 - 0x585  :  127 - 0x7f
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "11111111", -- 1416 - 0x588  :  255 - 0xff -- Sprite 0xb1
    "10001111", -- 1417 - 0x589  :  143 - 0x8f
    "10000000", -- 1418 - 0x58a  :  128 - 0x80
    "11110000", -- 1419 - 0x58b  :  240 - 0xf0
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11111111", -- 1421 - 0x58d  :  255 - 0xff
    "01111111", -- 1422 - 0x58e  :  127 - 0x7f
    "00001111", -- 1423 - 0x58f  :   15 - 0xf
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0xb2
    "11000000", -- 1425 - 0x591  :  192 - 0xc0
    "11110000", -- 1426 - 0x592  :  240 - 0xf0
    "11111100", -- 1427 - 0x593  :  252 - 0xfc
    "11111110", -- 1428 - 0x594  :  254 - 0xfe
    "11111110", -- 1429 - 0x595  :  254 - 0xfe
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff -- Sprite 0xb3
    "11110001", -- 1433 - 0x599  :  241 - 0xf1
    "00000001", -- 1434 - 0x59a  :    1 - 0x1
    "00001111", -- 1435 - 0x59b  :   15 - 0xf
    "11111111", -- 1436 - 0x59c  :  255 - 0xff
    "11111111", -- 1437 - 0x59d  :  255 - 0xff
    "11111110", -- 1438 - 0x59e  :  254 - 0xfe
    "11110000", -- 1439 - 0x59f  :  240 - 0xf0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0xb4
    "00000011", -- 1441 - 0x5a1  :    3 - 0x3
    "00001110", -- 1442 - 0x5a2  :   14 - 0xe
    "00110101", -- 1443 - 0x5a3  :   53 - 0x35
    "01101110", -- 1444 - 0x5a4  :  110 - 0x6e
    "01010101", -- 1445 - 0x5a5  :   85 - 0x55
    "10111010", -- 1446 - 0x5a6  :  186 - 0xba
    "11010111", -- 1447 - 0x5a7  :  215 - 0xd7
    "11111010", -- 1448 - 0x5a8  :  250 - 0xfa -- Sprite 0xb5
    "10001111", -- 1449 - 0x5a9  :  143 - 0x8f
    "10000000", -- 1450 - 0x5aa  :  128 - 0x80
    "11110000", -- 1451 - 0x5ab  :  240 - 0xf0
    "10101111", -- 1452 - 0x5ac  :  175 - 0xaf
    "11010101", -- 1453 - 0x5ad  :  213 - 0xd5
    "01111010", -- 1454 - 0x5ae  :  122 - 0x7a
    "00001111", -- 1455 - 0x5af  :   15 - 0xf
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "11000000", -- 1457 - 0x5b1  :  192 - 0xc0
    "10110000", -- 1458 - 0x5b2  :  176 - 0xb0
    "01011100", -- 1459 - 0x5b3  :   92 - 0x5c
    "11101010", -- 1460 - 0x5b4  :  234 - 0xea
    "01011110", -- 1461 - 0x5b5  :   94 - 0x5e
    "10101011", -- 1462 - 0x5b6  :  171 - 0xab
    "01110101", -- 1463 - 0x5b7  :  117 - 0x75
    "10101111", -- 1464 - 0x5b8  :  175 - 0xaf -- Sprite 0xb7
    "11110001", -- 1465 - 0x5b9  :  241 - 0xf1
    "00000001", -- 1466 - 0x5ba  :    1 - 0x1
    "00001111", -- 1467 - 0x5bb  :   15 - 0xf
    "11111011", -- 1468 - 0x5bc  :  251 - 0xfb
    "01010101", -- 1469 - 0x5bd  :   85 - 0x55
    "10101110", -- 1470 - 0x5be  :  174 - 0xae
    "11110000", -- 1471 - 0x5bf  :  240 - 0xf0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0xb8
    "00000011", -- 1473 - 0x5c1  :    3 - 0x3
    "00001100", -- 1474 - 0x5c2  :   12 - 0xc
    "00110000", -- 1475 - 0x5c3  :   48 - 0x30
    "01000100", -- 1476 - 0x5c4  :   68 - 0x44
    "01000000", -- 1477 - 0x5c5  :   64 - 0x40
    "10010000", -- 1478 - 0x5c6  :  144 - 0x90
    "10000010", -- 1479 - 0x5c7  :  130 - 0x82
    "11110000", -- 1480 - 0x5c8  :  240 - 0xf0 -- Sprite 0xb9
    "11111111", -- 1481 - 0x5c9  :  255 - 0xff
    "11111111", -- 1482 - 0x5ca  :  255 - 0xff
    "11111111", -- 1483 - 0x5cb  :  255 - 0xff
    "10001111", -- 1484 - 0x5cc  :  143 - 0x8f
    "10000000", -- 1485 - 0x5cd  :  128 - 0x80
    "01110000", -- 1486 - 0x5ce  :  112 - 0x70
    "00001111", -- 1487 - 0x5cf  :   15 - 0xf
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0xba
    "11000000", -- 1489 - 0x5d1  :  192 - 0xc0
    "00110000", -- 1490 - 0x5d2  :   48 - 0x30
    "00001100", -- 1491 - 0x5d3  :   12 - 0xc
    "01000010", -- 1492 - 0x5d4  :   66 - 0x42
    "00001010", -- 1493 - 0x5d5  :   10 - 0xa
    "00000001", -- 1494 - 0x5d6  :    1 - 0x1
    "00100001", -- 1495 - 0x5d7  :   33 - 0x21
    "00001111", -- 1496 - 0x5d8  :   15 - 0xf -- Sprite 0xbb
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111111", -- 1499 - 0x5db  :  255 - 0xff
    "11110001", -- 1500 - 0x5dc  :  241 - 0xf1
    "00000001", -- 1501 - 0x5dd  :    1 - 0x1
    "00001110", -- 1502 - 0x5de  :   14 - 0xe
    "11110000", -- 1503 - 0x5df  :  240 - 0xf0
    "11110011", -- 1504 - 0x5e0  :  243 - 0xf3 -- Sprite 0xbc
    "11111111", -- 1505 - 0x5e1  :  255 - 0xff
    "11000100", -- 1506 - 0x5e2  :  196 - 0xc4
    "11000000", -- 1507 - 0x5e3  :  192 - 0xc0
    "01000000", -- 1508 - 0x5e4  :   64 - 0x40
    "01100011", -- 1509 - 0x5e5  :   99 - 0x63
    "11000111", -- 1510 - 0x5e6  :  199 - 0xc7
    "11000110", -- 1511 - 0x5e7  :  198 - 0xc6
    "11000110", -- 1512 - 0x5e8  :  198 - 0xc6 -- Sprite 0xbd
    "11000110", -- 1513 - 0x5e9  :  198 - 0xc6
    "01100011", -- 1514 - 0x5ea  :   99 - 0x63
    "01000000", -- 1515 - 0x5eb  :   64 - 0x40
    "11000000", -- 1516 - 0x5ec  :  192 - 0xc0
    "11000100", -- 1517 - 0x5ed  :  196 - 0xc4
    "11001100", -- 1518 - 0x5ee  :  204 - 0xcc
    "11110011", -- 1519 - 0x5ef  :  243 - 0xf3
    "11001111", -- 1520 - 0x5f0  :  207 - 0xcf -- Sprite 0xbe
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "00100001", -- 1522 - 0x5f2  :   33 - 0x21
    "00000001", -- 1523 - 0x5f3  :    1 - 0x1
    "00000010", -- 1524 - 0x5f4  :    2 - 0x2
    "11000110", -- 1525 - 0x5f5  :  198 - 0xc6
    "11100001", -- 1526 - 0x5f6  :  225 - 0xe1
    "00100001", -- 1527 - 0x5f7  :   33 - 0x21
    "00100001", -- 1528 - 0x5f8  :   33 - 0x21 -- Sprite 0xbf
    "00100001", -- 1529 - 0x5f9  :   33 - 0x21
    "11000110", -- 1530 - 0x5fa  :  198 - 0xc6
    "00000010", -- 1531 - 0x5fb  :    2 - 0x2
    "00000001", -- 1532 - 0x5fc  :    1 - 0x1
    "00100001", -- 1533 - 0x5fd  :   33 - 0x21
    "00110001", -- 1534 - 0x5fe  :   49 - 0x31
    "11001111", -- 1535 - 0x5ff  :  207 - 0xcf
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "01010000", -- 1537 - 0x601  :   80 - 0x50
    "10110011", -- 1538 - 0x602  :  179 - 0xb3
    "10010111", -- 1539 - 0x603  :  151 - 0x97
    "10011111", -- 1540 - 0x604  :  159 - 0x9f
    "01101111", -- 1541 - 0x605  :  111 - 0x6f
    "00011111", -- 1542 - 0x606  :   31 - 0x1f
    "00011111", -- 1543 - 0x607  :   31 - 0x1f
    "00011111", -- 1544 - 0x608  :   31 - 0x1f -- Sprite 0xc1
    "00011111", -- 1545 - 0x609  :   31 - 0x1f
    "00001111", -- 1546 - 0x60a  :   15 - 0xf
    "00000111", -- 1547 - 0x60b  :    7 - 0x7
    "00011101", -- 1548 - 0x60c  :   29 - 0x1d
    "00101100", -- 1549 - 0x60d  :   44 - 0x2c
    "01010100", -- 1550 - 0x60e  :   84 - 0x54
    "01111100", -- 1551 - 0x60f  :  124 - 0x7c
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00001010", -- 1553 - 0x611  :   10 - 0xa
    "11001101", -- 1554 - 0x612  :  205 - 0xcd
    "11101001", -- 1555 - 0x613  :  233 - 0xe9
    "11111001", -- 1556 - 0x614  :  249 - 0xf9
    "11110110", -- 1557 - 0x615  :  246 - 0xf6
    "11110000", -- 1558 - 0x616  :  240 - 0xf0
    "11111000", -- 1559 - 0x617  :  248 - 0xf8
    "11111000", -- 1560 - 0x618  :  248 - 0xf8 -- Sprite 0xc3
    "11111000", -- 1561 - 0x619  :  248 - 0xf8
    "11110000", -- 1562 - 0x61a  :  240 - 0xf0
    "11000000", -- 1563 - 0x61b  :  192 - 0xc0
    "10111000", -- 1564 - 0x61c  :  184 - 0xb8
    "00110100", -- 1565 - 0x61d  :   52 - 0x34
    "00101010", -- 1566 - 0x61e  :   42 - 0x2a
    "00111110", -- 1567 - 0x61f  :   62 - 0x3e
    "00000101", -- 1568 - 0x620  :    5 - 0x5 -- Sprite 0xc4
    "00001010", -- 1569 - 0x621  :   10 - 0xa
    "00001000", -- 1570 - 0x622  :    8 - 0x8
    "00001111", -- 1571 - 0x623  :   15 - 0xf
    "00000001", -- 1572 - 0x624  :    1 - 0x1
    "00000011", -- 1573 - 0x625  :    3 - 0x3
    "00000111", -- 1574 - 0x626  :    7 - 0x7
    "00001111", -- 1575 - 0x627  :   15 - 0xf
    "00001111", -- 1576 - 0x628  :   15 - 0xf -- Sprite 0xc5
    "11101111", -- 1577 - 0x629  :  239 - 0xef
    "11011111", -- 1578 - 0x62a  :  223 - 0xdf
    "10101111", -- 1579 - 0x62b  :  175 - 0xaf
    "01100111", -- 1580 - 0x62c  :  103 - 0x67
    "00001101", -- 1581 - 0x62d  :   13 - 0xd
    "00001010", -- 1582 - 0x62e  :   10 - 0xa
    "00000111", -- 1583 - 0x62f  :    7 - 0x7
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0xc6
    "10000000", -- 1585 - 0x631  :  128 - 0x80
    "10000000", -- 1586 - 0x632  :  128 - 0x80
    "11110000", -- 1587 - 0x633  :  240 - 0xf0
    "11111000", -- 1588 - 0x634  :  248 - 0xf8
    "11111100", -- 1589 - 0x635  :  252 - 0xfc
    "11111100", -- 1590 - 0x636  :  252 - 0xfc
    "11111100", -- 1591 - 0x637  :  252 - 0xfc
    "11111100", -- 1592 - 0x638  :  252 - 0xfc -- Sprite 0xc7
    "11111110", -- 1593 - 0x639  :  254 - 0xfe
    "11111001", -- 1594 - 0x63a  :  249 - 0xf9
    "11111010", -- 1595 - 0x63b  :  250 - 0xfa
    "11101001", -- 1596 - 0x63c  :  233 - 0xe9
    "00001110", -- 1597 - 0x63d  :   14 - 0xe
    "10000000", -- 1598 - 0x63e  :  128 - 0x80
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "11000000", -- 1601 - 0x641  :  192 - 0xc0
    "10100000", -- 1602 - 0x642  :  160 - 0xa0
    "11010011", -- 1603 - 0x643  :  211 - 0xd3
    "10110111", -- 1604 - 0x644  :  183 - 0xb7
    "11111111", -- 1605 - 0x645  :  255 - 0xff
    "00001111", -- 1606 - 0x646  :   15 - 0xf
    "00011111", -- 1607 - 0x647  :   31 - 0x1f
    "00011111", -- 1608 - 0x648  :   31 - 0x1f -- Sprite 0xc9
    "00001111", -- 1609 - 0x649  :   15 - 0xf
    "11110111", -- 1610 - 0x64a  :  247 - 0xf7
    "10110111", -- 1611 - 0x64b  :  183 - 0xb7
    "11010011", -- 1612 - 0x64c  :  211 - 0xd3
    "10100000", -- 1613 - 0x64d  :  160 - 0xa0
    "11000000", -- 1614 - 0x64e  :  192 - 0xc0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00011100", -- 1616 - 0x650  :   28 - 0x1c -- Sprite 0xca
    "00100010", -- 1617 - 0x651  :   34 - 0x22
    "00100100", -- 1618 - 0x652  :   36 - 0x24
    "11011110", -- 1619 - 0x653  :  222 - 0xde
    "11110000", -- 1620 - 0x654  :  240 - 0xf0
    "11111000", -- 1621 - 0x655  :  248 - 0xf8
    "11111100", -- 1622 - 0x656  :  252 - 0xfc
    "11111100", -- 1623 - 0x657  :  252 - 0xfc
    "11111100", -- 1624 - 0x658  :  252 - 0xfc -- Sprite 0xcb
    "11111100", -- 1625 - 0x659  :  252 - 0xfc
    "11111000", -- 1626 - 0x65a  :  248 - 0xf8
    "11110000", -- 1627 - 0x65b  :  240 - 0xf0
    "10011110", -- 1628 - 0x65c  :  158 - 0x9e
    "00100100", -- 1629 - 0x65d  :   36 - 0x24
    "00100010", -- 1630 - 0x65e  :   34 - 0x22
    "00011100", -- 1631 - 0x65f  :   28 - 0x1c
    "00001110", -- 1632 - 0x660  :   14 - 0xe -- Sprite 0xcc
    "00010110", -- 1633 - 0x661  :   22 - 0x16
    "00011010", -- 1634 - 0x662  :   26 - 0x1a
    "00000100", -- 1635 - 0x663  :    4 - 0x4
    "01101111", -- 1636 - 0x664  :  111 - 0x6f
    "10111111", -- 1637 - 0x665  :  191 - 0xbf
    "11011111", -- 1638 - 0x666  :  223 - 0xdf
    "10111111", -- 1639 - 0x667  :  191 - 0xbf
    "01011111", -- 1640 - 0x668  :   95 - 0x5f -- Sprite 0xcd
    "00011111", -- 1641 - 0x669  :   31 - 0x1f
    "00011111", -- 1642 - 0x66a  :   31 - 0x1f
    "00001111", -- 1643 - 0x66b  :   15 - 0xf
    "00111111", -- 1644 - 0x66c  :   63 - 0x3f
    "00100011", -- 1645 - 0x66d  :   35 - 0x23
    "00101010", -- 1646 - 0x66e  :   42 - 0x2a
    "00010100", -- 1647 - 0x66f  :   20 - 0x14
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "10001110", -- 1652 - 0x674  :  142 - 0x8e
    "11001001", -- 1653 - 0x675  :  201 - 0xc9
    "11101010", -- 1654 - 0x676  :  234 - 0xea
    "11111001", -- 1655 - 0x677  :  249 - 0xf9
    "11111110", -- 1656 - 0x678  :  254 - 0xfe -- Sprite 0xcf
    "11111000", -- 1657 - 0x679  :  248 - 0xf8
    "11111000", -- 1658 - 0x67a  :  248 - 0xf8
    "11111000", -- 1659 - 0x67b  :  248 - 0xf8
    "11110000", -- 1660 - 0x67c  :  240 - 0xf0
    "11100000", -- 1661 - 0x67d  :  224 - 0xe0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000100", -- 1666 - 0x682  :    4 - 0x4
    "00100110", -- 1667 - 0x683  :   38 - 0x26
    "00101011", -- 1668 - 0x684  :   43 - 0x2b
    "01110001", -- 1669 - 0x685  :  113 - 0x71
    "01000000", -- 1670 - 0x686  :   64 - 0x40
    "01000111", -- 1671 - 0x687  :   71 - 0x47
    "10001111", -- 1672 - 0x688  :  143 - 0x8f -- Sprite 0xd1
    "10001111", -- 1673 - 0x689  :  143 - 0x8f
    "01001111", -- 1674 - 0x68a  :   79 - 0x4f
    "01001111", -- 1675 - 0x68b  :   79 - 0x4f
    "00111111", -- 1676 - 0x68c  :   63 - 0x3f
    "00010011", -- 1677 - 0x68d  :   19 - 0x13
    "00010001", -- 1678 - 0x68e  :   17 - 0x11
    "00011111", -- 1679 - 0x68f  :   31 - 0x1f
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0xd2
    "10000000", -- 1681 - 0x691  :  128 - 0x80
    "11001000", -- 1682 - 0x692  :  200 - 0xc8
    "11010100", -- 1683 - 0x693  :  212 - 0xd4
    "00100100", -- 1684 - 0x694  :   36 - 0x24
    "00000010", -- 1685 - 0x695  :    2 - 0x2
    "00000010", -- 1686 - 0x696  :    2 - 0x2
    "11110010", -- 1687 - 0x697  :  242 - 0xf2
    "11110010", -- 1688 - 0x698  :  242 - 0xf2 -- Sprite 0xd3
    "11110010", -- 1689 - 0x699  :  242 - 0xf2
    "11110100", -- 1690 - 0x69a  :  244 - 0xf4
    "11110100", -- 1691 - 0x69b  :  244 - 0xf4
    "11110100", -- 1692 - 0x69c  :  244 - 0xf4
    "11001000", -- 1693 - 0x69d  :  200 - 0xc8
    "01000100", -- 1694 - 0x69e  :   68 - 0x44
    "01111100", -- 1695 - 0x69f  :  124 - 0x7c
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00001001", -- 1699 - 0x6a3  :    9 - 0x9
    "00011010", -- 1700 - 0x6a4  :   26 - 0x1a
    "00010100", -- 1701 - 0x6a5  :   20 - 0x14
    "00100000", -- 1702 - 0x6a6  :   32 - 0x20
    "01000111", -- 1703 - 0x6a7  :   71 - 0x47
    "10001111", -- 1704 - 0x6a8  :  143 - 0x8f -- Sprite 0xd5
    "10001111", -- 1705 - 0x6a9  :  143 - 0x8f
    "01001111", -- 1706 - 0x6aa  :   79 - 0x4f
    "01001111", -- 1707 - 0x6ab  :   79 - 0x4f
    "00111111", -- 1708 - 0x6ac  :   63 - 0x3f
    "01000111", -- 1709 - 0x6ad  :   71 - 0x47
    "00100010", -- 1710 - 0x6ae  :   34 - 0x22
    "00011100", -- 1711 - 0x6af  :   28 - 0x1c
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "01000000", -- 1713 - 0x6b1  :   64 - 0x40
    "11000000", -- 1714 - 0x6b2  :  192 - 0xc0
    "00101100", -- 1715 - 0x6b3  :   44 - 0x2c
    "00110100", -- 1716 - 0x6b4  :   52 - 0x34
    "00000100", -- 1717 - 0x6b5  :    4 - 0x4
    "00000010", -- 1718 - 0x6b6  :    2 - 0x2
    "11110010", -- 1719 - 0x6b7  :  242 - 0xf2
    "11110010", -- 1720 - 0x6b8  :  242 - 0xf2 -- Sprite 0xd7
    "11110010", -- 1721 - 0x6b9  :  242 - 0xf2
    "11110100", -- 1722 - 0x6ba  :  244 - 0xf4
    "11110111", -- 1723 - 0x6bb  :  247 - 0xf7
    "11111101", -- 1724 - 0x6bc  :  253 - 0xfd
    "11100001", -- 1725 - 0x6bd  :  225 - 0xe1
    "00010010", -- 1726 - 0x6be  :   18 - 0x12
    "00001100", -- 1727 - 0x6bf  :   12 - 0xc
    "01111000", -- 1728 - 0x6c0  :  120 - 0x78 -- Sprite 0xd8
    "01001110", -- 1729 - 0x6c1  :   78 - 0x4e
    "11000010", -- 1730 - 0x6c2  :  194 - 0xc2
    "10011010", -- 1731 - 0x6c3  :  154 - 0x9a
    "10011011", -- 1732 - 0x6c4  :  155 - 0x9b
    "11011001", -- 1733 - 0x6c5  :  217 - 0xd9
    "01100011", -- 1734 - 0x6c6  :   99 - 0x63
    "00111110", -- 1735 - 0x6c7  :   62 - 0x3e
    "00011110", -- 1736 - 0x6c8  :   30 - 0x1e -- Sprite 0xd9
    "01110001", -- 1737 - 0x6c9  :  113 - 0x71
    "01001001", -- 1738 - 0x6ca  :   73 - 0x49
    "10111001", -- 1739 - 0x6cb  :  185 - 0xb9
    "10011101", -- 1740 - 0x6cc  :  157 - 0x9d
    "01010010", -- 1741 - 0x6cd  :   82 - 0x52
    "01110010", -- 1742 - 0x6ce  :  114 - 0x72
    "00011110", -- 1743 - 0x6cf  :   30 - 0x1e
    "01100000", -- 1744 - 0x6d0  :   96 - 0x60 -- Sprite 0xda
    "01011110", -- 1745 - 0x6d1  :   94 - 0x5e
    "10001001", -- 1746 - 0x6d2  :  137 - 0x89
    "10111101", -- 1747 - 0x6d3  :  189 - 0xbd
    "10011101", -- 1748 - 0x6d4  :  157 - 0x9d
    "11010011", -- 1749 - 0x6d5  :  211 - 0xd3
    "01000110", -- 1750 - 0x6d6  :   70 - 0x46
    "01111100", -- 1751 - 0x6d7  :  124 - 0x7c
    "00011110", -- 1752 - 0x6d8  :   30 - 0x1e -- Sprite 0xdb
    "00100011", -- 1753 - 0x6d9  :   35 - 0x23
    "01001001", -- 1754 - 0x6da  :   73 - 0x49
    "10111101", -- 1755 - 0x6db  :  189 - 0xbd
    "10011001", -- 1756 - 0x6dc  :  153 - 0x99
    "01000011", -- 1757 - 0x6dd  :   67 - 0x43
    "01101110", -- 1758 - 0x6de  :  110 - 0x6e
    "00011000", -- 1759 - 0x6df  :   24 - 0x18
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000001", -- 1762 - 0x6e2  :    1 - 0x1
    "00000010", -- 1763 - 0x6e3  :    2 - 0x2
    "00000100", -- 1764 - 0x6e4  :    4 - 0x4
    "00000010", -- 1765 - 0x6e5  :    2 - 0x2
    "00011110", -- 1766 - 0x6e6  :   30 - 0x1e
    "00010000", -- 1767 - 0x6e7  :   16 - 0x10
    "00001000", -- 1768 - 0x6e8  :    8 - 0x8 -- Sprite 0xdd
    "00001101", -- 1769 - 0x6e9  :   13 - 0xd
    "00111010", -- 1770 - 0x6ea  :   58 - 0x3a
    "00100101", -- 1771 - 0x6eb  :   37 - 0x25
    "00011011", -- 1772 - 0x6ec  :   27 - 0x1b
    "00001111", -- 1773 - 0x6ed  :   15 - 0xf
    "00000111", -- 1774 - 0x6ee  :    7 - 0x7
    "00000011", -- 1775 - 0x6ef  :    3 - 0x3
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0xde
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "11000000", -- 1779 - 0x6f3  :  192 - 0xc0
    "01000000", -- 1780 - 0x6f4  :   64 - 0x40
    "01011000", -- 1781 - 0x6f5  :   88 - 0x58
    "01101000", -- 1782 - 0x6f6  :  104 - 0x68
    "00001000", -- 1783 - 0x6f7  :    8 - 0x8
    "00010000", -- 1784 - 0x6f8  :   16 - 0x10 -- Sprite 0xdf
    "01011100", -- 1785 - 0x6f9  :   92 - 0x5c
    "10101000", -- 1786 - 0x6fa  :  168 - 0xa8
    "11011000", -- 1787 - 0x6fb  :  216 - 0xd8
    "10111000", -- 1788 - 0x6fc  :  184 - 0xb8
    "11110000", -- 1789 - 0x6fd  :  240 - 0xf0
    "11100000", -- 1790 - 0x6fe  :  224 - 0xe0
    "11000000", -- 1791 - 0x6ff  :  192 - 0xc0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00010011", -- 1795 - 0x703  :   19 - 0x13
    "00010011", -- 1796 - 0x704  :   19 - 0x13
    "00110111", -- 1797 - 0x705  :   55 - 0x37
    "00110111", -- 1798 - 0x706  :   55 - 0x37
    "00000111", -- 1799 - 0x707  :    7 - 0x7
    "00000111", -- 1800 - 0x708  :    7 - 0x7 -- Sprite 0xe1
    "00000100", -- 1801 - 0x709  :    4 - 0x4
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00100000", -- 1805 - 0x70d  :   32 - 0x20
    "01110000", -- 1806 - 0x70e  :  112 - 0x70
    "11111000", -- 1807 - 0x70f  :  248 - 0xf8
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0xe2
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "11111000", -- 1811 - 0x713  :  248 - 0xf8
    "11111100", -- 1812 - 0x714  :  252 - 0xfc
    "11111100", -- 1813 - 0x715  :  252 - 0xfc
    "11111100", -- 1814 - 0x716  :  252 - 0xfc
    "11111101", -- 1815 - 0x717  :  253 - 0xfd
    "11111100", -- 1816 - 0x718  :  252 - 0xfc -- Sprite 0xe3
    "00011100", -- 1817 - 0x719  :   28 - 0x1c
    "11000000", -- 1818 - 0x71a  :  192 - 0xc0
    "11100000", -- 1819 - 0x71b  :  224 - 0xe0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000110", -- 1822 - 0x71e  :    6 - 0x6
    "00001111", -- 1823 - 0x71f  :   15 - 0xf
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00010011", -- 1827 - 0x723  :   19 - 0x13
    "00010011", -- 1828 - 0x724  :   19 - 0x13
    "00110111", -- 1829 - 0x725  :   55 - 0x37
    "00110111", -- 1830 - 0x726  :   55 - 0x37
    "00000111", -- 1831 - 0x727  :    7 - 0x7
    "00000111", -- 1832 - 0x728  :    7 - 0x7 -- Sprite 0xe5
    "00000100", -- 1833 - 0x729  :    4 - 0x4
    "00000001", -- 1834 - 0x72a  :    1 - 0x1
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00100000", -- 1837 - 0x72d  :   32 - 0x20
    "01110000", -- 1838 - 0x72e  :  112 - 0x70
    "11111000", -- 1839 - 0x72f  :  248 - 0xf8
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "11111100", -- 1843 - 0x733  :  252 - 0xfc
    "11111100", -- 1844 - 0x734  :  252 - 0xfc
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11111100", -- 1846 - 0x736  :  252 - 0xfc
    "11111101", -- 1847 - 0x737  :  253 - 0xfd
    "11111100", -- 1848 - 0x738  :  252 - 0xfc -- Sprite 0xe7
    "00001100", -- 1849 - 0x739  :   12 - 0xc
    "11000000", -- 1850 - 0x73a  :  192 - 0xc0
    "11110000", -- 1851 - 0x73b  :  240 - 0xf0
    "11110000", -- 1852 - 0x73c  :  240 - 0xf0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000110", -- 1854 - 0x73e  :    6 - 0x6
    "00001111", -- 1855 - 0x73f  :   15 - 0xf
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "01111111", -- 1858 - 0x742  :  127 - 0x7f
    "01111111", -- 1859 - 0x743  :  127 - 0x7f
    "01111111", -- 1860 - 0x744  :  127 - 0x7f
    "00111111", -- 1861 - 0x745  :   63 - 0x3f
    "00111111", -- 1862 - 0x746  :   63 - 0x3f
    "00111111", -- 1863 - 0x747  :   63 - 0x3f
    "00111100", -- 1864 - 0x748  :   60 - 0x3c -- Sprite 0xe9
    "00111110", -- 1865 - 0x749  :   62 - 0x3e
    "00011111", -- 1866 - 0x74a  :   31 - 0x1f
    "00001111", -- 1867 - 0x74b  :   15 - 0xf
    "00000111", -- 1868 - 0x74c  :    7 - 0x7
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0xea
    "11111110", -- 1873 - 0x751  :  254 - 0xfe
    "11111110", -- 1874 - 0x752  :  254 - 0xfe
    "11111100", -- 1875 - 0x753  :  252 - 0xfc
    "11111000", -- 1876 - 0x754  :  248 - 0xf8
    "11110000", -- 1877 - 0x755  :  240 - 0xf0
    "10110000", -- 1878 - 0x756  :  176 - 0xb0
    "00111001", -- 1879 - 0x757  :   57 - 0x39
    "00011111", -- 1880 - 0x758  :   31 - 0x1f -- Sprite 0xeb
    "11001111", -- 1881 - 0x759  :  207 - 0xcf
    "11000110", -- 1882 - 0x75a  :  198 - 0xc6
    "10000000", -- 1883 - 0x75b  :  128 - 0x80
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00001100", -- 1894 - 0x766  :   12 - 0xc
    "00001100", -- 1895 - 0x767  :   12 - 0xc
    "00110000", -- 1896 - 0x768  :   48 - 0x30 -- Sprite 0xed
    "01000011", -- 1897 - 0x769  :   67 - 0x43
    "01000000", -- 1898 - 0x76a  :   64 - 0x40
    "01100000", -- 1899 - 0x76b  :   96 - 0x60
    "00000011", -- 1900 - 0x76c  :    3 - 0x3
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "01111111", -- 1902 - 0x76e  :  127 - 0x7f
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00110000", -- 1910 - 0x776  :   48 - 0x30
    "00110000", -- 1911 - 0x777  :   48 - 0x30
    "00001110", -- 1912 - 0x778  :   14 - 0xe -- Sprite 0xef
    "11001011", -- 1913 - 0x779  :  203 - 0xcb
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "11000000", -- 1916 - 0x77c  :  192 - 0xc0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "11111110", -- 1918 - 0x77e  :  254 - 0xfe
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00001100", -- 1926 - 0x786  :   12 - 0xc
    "00001100", -- 1927 - 0x787  :   12 - 0xc
    "00110000", -- 1928 - 0x788  :   48 - 0x30 -- Sprite 0xf1
    "00100011", -- 1929 - 0x789  :   35 - 0x23
    "00100000", -- 1930 - 0x78a  :   32 - 0x20
    "01100000", -- 1931 - 0x78b  :   96 - 0x60
    "00000011", -- 1932 - 0x78c  :    3 - 0x3
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "01111111", -- 1934 - 0x78e  :  127 - 0x7f
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00110000", -- 1942 - 0x796  :   48 - 0x30
    "00110000", -- 1943 - 0x797  :   48 - 0x30
    "00001001", -- 1944 - 0x798  :    9 - 0x9 -- Sprite 0xf3
    "11001111", -- 1945 - 0x799  :  207 - 0xcf
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "11000000", -- 1948 - 0x79c  :  192 - 0xc0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "11111110", -- 1950 - 0x79e  :  254 - 0xfe
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00111111", -- 1952 - 0x7a0  :   63 - 0x3f -- Sprite 0xf4
    "00110101", -- 1953 - 0x7a1  :   53 - 0x35
    "00011010", -- 1954 - 0x7a2  :   26 - 0x1a
    "00001101", -- 1955 - 0x7a3  :   13 - 0xd
    "00001010", -- 1956 - 0x7a4  :   10 - 0xa
    "00001101", -- 1957 - 0x7a5  :   13 - 0xd
    "00001000", -- 1958 - 0x7a6  :    8 - 0x8
    "00111000", -- 1959 - 0x7a7  :   56 - 0x38
    "01110011", -- 1960 - 0x7a8  :  115 - 0x73 -- Sprite 0xf5
    "11000100", -- 1961 - 0x7a9  :  196 - 0xc4
    "11000100", -- 1962 - 0x7aa  :  196 - 0xc4
    "11000000", -- 1963 - 0x7ab  :  192 - 0xc0
    "11000001", -- 1964 - 0x7ac  :  193 - 0xc1
    "11000000", -- 1965 - 0x7ad  :  192 - 0xc0
    "01100001", -- 1966 - 0x7ae  :   97 - 0x61
    "00111111", -- 1967 - 0x7af  :   63 - 0x3f
    "11111100", -- 1968 - 0x7b0  :  252 - 0xfc -- Sprite 0xf6
    "01010100", -- 1969 - 0x7b1  :   84 - 0x54
    "10101000", -- 1970 - 0x7b2  :  168 - 0xa8
    "01010000", -- 1971 - 0x7b3  :   80 - 0x50
    "10110000", -- 1972 - 0x7b4  :  176 - 0xb0
    "01010000", -- 1973 - 0x7b5  :   80 - 0x50
    "10010000", -- 1974 - 0x7b6  :  144 - 0x90
    "00011100", -- 1975 - 0x7b7  :   28 - 0x1c
    "10000110", -- 1976 - 0x7b8  :  134 - 0x86 -- Sprite 0xf7
    "01000010", -- 1977 - 0x7b9  :   66 - 0x42
    "01000111", -- 1978 - 0x7ba  :   71 - 0x47
    "01000001", -- 1979 - 0x7bb  :   65 - 0x41
    "10000011", -- 1980 - 0x7bc  :  131 - 0x83
    "00000001", -- 1981 - 0x7bd  :    1 - 0x1
    "10000110", -- 1982 - 0x7be  :  134 - 0x86
    "11111100", -- 1983 - 0x7bf  :  252 - 0xfc
    "11100100", -- 1984 - 0x7c0  :  228 - 0xe4 -- Sprite 0xf8
    "11100100", -- 1985 - 0x7c1  :  228 - 0xe4
    "11101111", -- 1986 - 0x7c2  :  239 - 0xef
    "11101111", -- 1987 - 0x7c3  :  239 - 0xef
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "01111111", -- 1990 - 0x7c6  :  127 - 0x7f
    "01111111", -- 1991 - 0x7c7  :  127 - 0x7f
    "00111111", -- 1992 - 0x7c8  :   63 - 0x3f -- Sprite 0xf9
    "01111111", -- 1993 - 0x7c9  :  127 - 0x7f
    "01111111", -- 1994 - 0x7ca  :  127 - 0x7f
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "00010011", -- 2000 - 0x7d0  :   19 - 0x13 -- Sprite 0xfa
    "00010011", -- 2001 - 0x7d1  :   19 - 0x13
    "11111011", -- 2002 - 0x7d2  :  251 - 0xfb
    "11111011", -- 2003 - 0x7d3  :  251 - 0xfb
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111110", -- 2006 - 0x7d6  :  254 - 0xfe
    "11111110", -- 2007 - 0x7d7  :  254 - 0xfe
    "11111110", -- 2008 - 0x7d8  :  254 - 0xfe -- Sprite 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "01111100", -- 2018 - 0x7e2  :  124 - 0x7c
    "11111110", -- 2019 - 0x7e3  :  254 - 0xfe
    "11111110", -- 2020 - 0x7e4  :  254 - 0xfe
    "01111100", -- 2021 - 0x7e5  :  124 - 0x7c
    "01000100", -- 2022 - 0x7e6  :   68 - 0x44
    "10000010", -- 2023 - 0x7e7  :  130 - 0x82
    "10000010", -- 2024 - 0x7e8  :  130 - 0x82 -- Sprite 0xfd
    "10000010", -- 2025 - 0x7e9  :  130 - 0x82
    "10000010", -- 2026 - 0x7ea  :  130 - 0x82
    "11000110", -- 2027 - 0x7eb  :  198 - 0xc6
    "11111110", -- 2028 - 0x7ec  :  254 - 0xfe
    "11111110", -- 2029 - 0x7ed  :  254 - 0xfe
    "10111010", -- 2030 - 0x7ee  :  186 - 0xba
    "01111100", -- 2031 - 0x7ef  :  124 - 0x7c
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00011001", -- 2033 - 0x7f1  :   25 - 0x19
    "00111110", -- 2034 - 0x7f2  :   62 - 0x3e
    "00111100", -- 2035 - 0x7f3  :   60 - 0x3c
    "00111100", -- 2036 - 0x7f4  :   60 - 0x3c
    "00111100", -- 2037 - 0x7f5  :   60 - 0x3c
    "00111110", -- 2038 - 0x7f6  :   62 - 0x3e
    "00011001", -- 2039 - 0x7f7  :   25 - 0x19
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "11111110", -- 2041 - 0x7f9  :  254 - 0xfe
    "00011101", -- 2042 - 0x7fa  :   29 - 0x1d
    "00001111", -- 2043 - 0x7fb  :   15 - 0xf
    "00001111", -- 2044 - 0x7fc  :   15 - 0xf
    "00001111", -- 2045 - 0x7fd  :   15 - 0xf
    "00011101", -- 2046 - 0x7fe  :   29 - 0x1d
    "11111110", -- 2047 - 0x7ff  :  254 - 0xfe
          -- Background pattern Table
    "11111111", -- 2048 - 0x800  :  255 - 0xff -- Background 0x0
    "11111111", -- 2049 - 0x801  :  255 - 0xff
    "11000000", -- 2050 - 0x802  :  192 - 0xc0
    "11000000", -- 2051 - 0x803  :  192 - 0xc0
    "11000000", -- 2052 - 0x804  :  192 - 0xc0
    "11000000", -- 2053 - 0x805  :  192 - 0xc0
    "11010101", -- 2054 - 0x806  :  213 - 0xd5
    "11111111", -- 2055 - 0x807  :  255 - 0xff
    "11111111", -- 2056 - 0x808  :  255 - 0xff -- Background 0x1
    "11111111", -- 2057 - 0x809  :  255 - 0xff
    "11001110", -- 2058 - 0x80a  :  206 - 0xce
    "11000110", -- 2059 - 0x80b  :  198 - 0xc6
    "11001110", -- 2060 - 0x80c  :  206 - 0xce
    "11000110", -- 2061 - 0x80d  :  198 - 0xc6
    "11101110", -- 2062 - 0x80e  :  238 - 0xee
    "11111111", -- 2063 - 0x80f  :  255 - 0xff
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Background 0x2
    "11111111", -- 2065 - 0x811  :  255 - 0xff
    "01110001", -- 2066 - 0x812  :  113 - 0x71
    "00110011", -- 2067 - 0x813  :   51 - 0x33
    "01110001", -- 2068 - 0x814  :  113 - 0x71
    "00110011", -- 2069 - 0x815  :   51 - 0x33
    "01110101", -- 2070 - 0x816  :  117 - 0x75
    "11111111", -- 2071 - 0x817  :  255 - 0xff
    "11111111", -- 2072 - 0x818  :  255 - 0xff -- Background 0x3
    "11111111", -- 2073 - 0x819  :  255 - 0xff
    "00000011", -- 2074 - 0x81a  :    3 - 0x3
    "00000001", -- 2075 - 0x81b  :    1 - 0x1
    "00000011", -- 2076 - 0x81c  :    3 - 0x3
    "00000001", -- 2077 - 0x81d  :    1 - 0x1
    "10101011", -- 2078 - 0x81e  :  171 - 0xab
    "11111111", -- 2079 - 0x81f  :  255 - 0xff
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Background 0x4
    "11111111", -- 2081 - 0x821  :  255 - 0xff
    "11100000", -- 2082 - 0x822  :  224 - 0xe0
    "11000110", -- 2083 - 0x823  :  198 - 0xc6
    "11000110", -- 2084 - 0x824  :  198 - 0xc6
    "11110110", -- 2085 - 0x825  :  246 - 0xf6
    "11110000", -- 2086 - 0x826  :  240 - 0xf0
    "11110001", -- 2087 - 0x827  :  241 - 0xf1
    "11000111", -- 2088 - 0x828  :  199 - 0xc7 -- Background 0x5
    "11001111", -- 2089 - 0x829  :  207 - 0xcf
    "11011111", -- 2090 - 0x82a  :  223 - 0xdf
    "11011111", -- 2091 - 0x82b  :  223 - 0xdf
    "11001110", -- 2092 - 0x82c  :  206 - 0xce
    "11100000", -- 2093 - 0x82d  :  224 - 0xe0
    "11111111", -- 2094 - 0x82e  :  255 - 0xff
    "11111111", -- 2095 - 0x82f  :  255 - 0xff
    "11111111", -- 2096 - 0x830  :  255 - 0xff -- Background 0x6
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "00000111", -- 2098 - 0x832  :    7 - 0x7
    "01100011", -- 2099 - 0x833  :   99 - 0x63
    "01100011", -- 2100 - 0x834  :   99 - 0x63
    "01101111", -- 2101 - 0x835  :  111 - 0x6f
    "00001111", -- 2102 - 0x836  :   15 - 0xf
    "10001111", -- 2103 - 0x837  :  143 - 0x8f
    "11100011", -- 2104 - 0x838  :  227 - 0xe3 -- Background 0x7
    "11110011", -- 2105 - 0x839  :  243 - 0xf3
    "11111011", -- 2106 - 0x83a  :  251 - 0xfb
    "11111011", -- 2107 - 0x83b  :  251 - 0xfb
    "01110011", -- 2108 - 0x83c  :  115 - 0x73
    "00000111", -- 2109 - 0x83d  :    7 - 0x7
    "11111111", -- 2110 - 0x83e  :  255 - 0xff
    "11111111", -- 2111 - 0x83f  :  255 - 0xff
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Background 0x8
    "11010101", -- 2113 - 0x841  :  213 - 0xd5
    "10101010", -- 2114 - 0x842  :  170 - 0xaa
    "11010101", -- 2115 - 0x843  :  213 - 0xd5
    "10101010", -- 2116 - 0x844  :  170 - 0xaa
    "11010101", -- 2117 - 0x845  :  213 - 0xd5
    "10101010", -- 2118 - 0x846  :  170 - 0xaa
    "11010101", -- 2119 - 0x847  :  213 - 0xd5
    "10101010", -- 2120 - 0x848  :  170 - 0xaa -- Background 0x9
    "11010101", -- 2121 - 0x849  :  213 - 0xd5
    "10101010", -- 2122 - 0x84a  :  170 - 0xaa
    "11010101", -- 2123 - 0x84b  :  213 - 0xd5
    "10101010", -- 2124 - 0x84c  :  170 - 0xaa
    "11110101", -- 2125 - 0x84d  :  245 - 0xf5
    "10101010", -- 2126 - 0x84e  :  170 - 0xaa
    "11111111", -- 2127 - 0x84f  :  255 - 0xff
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Background 0xa
    "01010101", -- 2129 - 0x851  :   85 - 0x55
    "10101111", -- 2130 - 0x852  :  175 - 0xaf
    "01010101", -- 2131 - 0x853  :   85 - 0x55
    "10101011", -- 2132 - 0x854  :  171 - 0xab
    "01010101", -- 2133 - 0x855  :   85 - 0x55
    "10101011", -- 2134 - 0x856  :  171 - 0xab
    "01010101", -- 2135 - 0x857  :   85 - 0x55
    "10101011", -- 2136 - 0x858  :  171 - 0xab -- Background 0xb
    "01010101", -- 2137 - 0x859  :   85 - 0x55
    "10101011", -- 2138 - 0x85a  :  171 - 0xab
    "01010101", -- 2139 - 0x85b  :   85 - 0x55
    "10101011", -- 2140 - 0x85c  :  171 - 0xab
    "01010101", -- 2141 - 0x85d  :   85 - 0x55
    "10101011", -- 2142 - 0x85e  :  171 - 0xab
    "11111111", -- 2143 - 0x85f  :  255 - 0xff
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Background 0xc
    "11010101", -- 2145 - 0x861  :  213 - 0xd5
    "10100000", -- 2146 - 0x862  :  160 - 0xa0
    "11010000", -- 2147 - 0x863  :  208 - 0xd0
    "10001111", -- 2148 - 0x864  :  143 - 0x8f
    "11001000", -- 2149 - 0x865  :  200 - 0xc8
    "10001000", -- 2150 - 0x866  :  136 - 0x88
    "11001000", -- 2151 - 0x867  :  200 - 0xc8
    "10001000", -- 2152 - 0x868  :  136 - 0x88 -- Background 0xd
    "11001000", -- 2153 - 0x869  :  200 - 0xc8
    "10001000", -- 2154 - 0x86a  :  136 - 0x88
    "11001111", -- 2155 - 0x86b  :  207 - 0xcf
    "10010000", -- 2156 - 0x86c  :  144 - 0x90
    "11100000", -- 2157 - 0x86d  :  224 - 0xe0
    "11101010", -- 2158 - 0x86e  :  234 - 0xea
    "11111111", -- 2159 - 0x86f  :  255 - 0xff
    "11111111", -- 2160 - 0x870  :  255 - 0xff -- Background 0xe
    "01011011", -- 2161 - 0x871  :   91 - 0x5b
    "00000111", -- 2162 - 0x872  :    7 - 0x7
    "00001001", -- 2163 - 0x873  :    9 - 0x9
    "11110011", -- 2164 - 0x874  :  243 - 0xf3
    "00010001", -- 2165 - 0x875  :   17 - 0x11
    "00010011", -- 2166 - 0x876  :   19 - 0x13
    "00010001", -- 2167 - 0x877  :   17 - 0x11
    "00010011", -- 2168 - 0x878  :   19 - 0x13 -- Background 0xf
    "00010001", -- 2169 - 0x879  :   17 - 0x11
    "00010011", -- 2170 - 0x87a  :   19 - 0x13
    "11110001", -- 2171 - 0x87b  :  241 - 0xf1
    "00001011", -- 2172 - 0x87c  :   11 - 0xb
    "00000101", -- 2173 - 0x87d  :    5 - 0x5
    "10101011", -- 2174 - 0x87e  :  171 - 0xab
    "11111111", -- 2175 - 0x87f  :  255 - 0xff
    "11010000", -- 2176 - 0x880  :  208 - 0xd0 -- Background 0x10
    "10010000", -- 2177 - 0x881  :  144 - 0x90
    "11011111", -- 2178 - 0x882  :  223 - 0xdf
    "10011010", -- 2179 - 0x883  :  154 - 0x9a
    "11010101", -- 2180 - 0x884  :  213 - 0xd5
    "10011111", -- 2181 - 0x885  :  159 - 0x9f
    "11010000", -- 2182 - 0x886  :  208 - 0xd0
    "10010000", -- 2183 - 0x887  :  144 - 0x90
    "00001001", -- 2184 - 0x888  :    9 - 0x9 -- Background 0x11
    "00001011", -- 2185 - 0x889  :   11 - 0xb
    "11111001", -- 2186 - 0x88a  :  249 - 0xf9
    "10101011", -- 2187 - 0x88b  :  171 - 0xab
    "01011001", -- 2188 - 0x88c  :   89 - 0x59
    "11111011", -- 2189 - 0x88d  :  251 - 0xfb
    "00001001", -- 2190 - 0x88e  :    9 - 0x9
    "00001011", -- 2191 - 0x88f  :   11 - 0xb
    "00011000", -- 2192 - 0x890  :   24 - 0x18 -- Background 0x12
    "00010100", -- 2193 - 0x891  :   20 - 0x14
    "00010100", -- 2194 - 0x892  :   20 - 0x14
    "00111010", -- 2195 - 0x893  :   58 - 0x3a
    "00111010", -- 2196 - 0x894  :   58 - 0x3a
    "01111010", -- 2197 - 0x895  :  122 - 0x7a
    "01111010", -- 2198 - 0x896  :  122 - 0x7a
    "01111010", -- 2199 - 0x897  :  122 - 0x7a
    "11111011", -- 2200 - 0x898  :  251 - 0xfb -- Background 0x13
    "11111101", -- 2201 - 0x899  :  253 - 0xfd
    "11111101", -- 2202 - 0x89a  :  253 - 0xfd
    "11111101", -- 2203 - 0x89b  :  253 - 0xfd
    "11111101", -- 2204 - 0x89c  :  253 - 0xfd
    "11111101", -- 2205 - 0x89d  :  253 - 0xfd
    "10000001", -- 2206 - 0x89e  :  129 - 0x81
    "11111111", -- 2207 - 0x89f  :  255 - 0xff
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x14
    "00000111", -- 2209 - 0x8a1  :    7 - 0x7
    "00000010", -- 2210 - 0x8a2  :    2 - 0x2
    "00000100", -- 2211 - 0x8a3  :    4 - 0x4
    "00000011", -- 2212 - 0x8a4  :    3 - 0x3
    "00000011", -- 2213 - 0x8a5  :    3 - 0x3
    "00001101", -- 2214 - 0x8a6  :   13 - 0xd
    "00010111", -- 2215 - 0x8a7  :   23 - 0x17
    "00101111", -- 2216 - 0x8a8  :   47 - 0x2f -- Background 0x15
    "01001111", -- 2217 - 0x8a9  :   79 - 0x4f
    "01001111", -- 2218 - 0x8aa  :   79 - 0x4f
    "01001111", -- 2219 - 0x8ab  :   79 - 0x4f
    "01001111", -- 2220 - 0x8ac  :   79 - 0x4f
    "00100111", -- 2221 - 0x8ad  :   39 - 0x27
    "00010000", -- 2222 - 0x8ae  :   16 - 0x10
    "00001111", -- 2223 - 0x8af  :   15 - 0xf
    "00000000", -- 2224 - 0x8b0  :    0 - 0x0 -- Background 0x16
    "11100000", -- 2225 - 0x8b1  :  224 - 0xe0
    "10100000", -- 2226 - 0x8b2  :  160 - 0xa0
    "00100000", -- 2227 - 0x8b3  :   32 - 0x20
    "11000000", -- 2228 - 0x8b4  :  192 - 0xc0
    "01000000", -- 2229 - 0x8b5  :   64 - 0x40
    "00110000", -- 2230 - 0x8b6  :   48 - 0x30
    "11101000", -- 2231 - 0x8b7  :  232 - 0xe8
    "11110100", -- 2232 - 0x8b8  :  244 - 0xf4 -- Background 0x17
    "11110010", -- 2233 - 0x8b9  :  242 - 0xf2
    "11110010", -- 2234 - 0x8ba  :  242 - 0xf2
    "11110010", -- 2235 - 0x8bb  :  242 - 0xf2
    "11110010", -- 2236 - 0x8bc  :  242 - 0xf2
    "11100100", -- 2237 - 0x8bd  :  228 - 0xe4
    "00001000", -- 2238 - 0x8be  :    8 - 0x8
    "11110000", -- 2239 - 0x8bf  :  240 - 0xf0
    "00111111", -- 2240 - 0x8c0  :   63 - 0x3f -- Background 0x18
    "01000000", -- 2241 - 0x8c1  :   64 - 0x40
    "01000000", -- 2242 - 0x8c2  :   64 - 0x40
    "10000000", -- 2243 - 0x8c3  :  128 - 0x80
    "10000000", -- 2244 - 0x8c4  :  128 - 0x80
    "01111111", -- 2245 - 0x8c5  :  127 - 0x7f
    "00000001", -- 2246 - 0x8c6  :    1 - 0x1
    "01111111", -- 2247 - 0x8c7  :  127 - 0x7f
    "11111100", -- 2248 - 0x8c8  :  252 - 0xfc -- Background 0x19
    "00000010", -- 2249 - 0x8c9  :    2 - 0x2
    "00000010", -- 2250 - 0x8ca  :    2 - 0x2
    "00000001", -- 2251 - 0x8cb  :    1 - 0x1
    "00000001", -- 2252 - 0x8cc  :    1 - 0x1
    "11111110", -- 2253 - 0x8cd  :  254 - 0xfe
    "10000000", -- 2254 - 0x8ce  :  128 - 0x80
    "11111110", -- 2255 - 0x8cf  :  254 - 0xfe
    "00000000", -- 2256 - 0x8d0  :    0 - 0x0 -- Background 0x1a
    "00000000", -- 2257 - 0x8d1  :    0 - 0x0
    "00111111", -- 2258 - 0x8d2  :   63 - 0x3f
    "01000000", -- 2259 - 0x8d3  :   64 - 0x40
    "01000000", -- 2260 - 0x8d4  :   64 - 0x40
    "10000000", -- 2261 - 0x8d5  :  128 - 0x80
    "10000000", -- 2262 - 0x8d6  :  128 - 0x80
    "01111111", -- 2263 - 0x8d7  :  127 - 0x7f
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- Background 0x1b
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "11111100", -- 2266 - 0x8da  :  252 - 0xfc
    "00000010", -- 2267 - 0x8db  :    2 - 0x2
    "00000010", -- 2268 - 0x8dc  :    2 - 0x2
    "00000001", -- 2269 - 0x8dd  :    1 - 0x1
    "00000001", -- 2270 - 0x8de  :    1 - 0x1
    "11111110", -- 2271 - 0x8df  :  254 - 0xfe
    "01111111", -- 2272 - 0x8e0  :  127 - 0x7f -- Background 0x1c
    "10000000", -- 2273 - 0x8e1  :  128 - 0x80
    "10000000", -- 2274 - 0x8e2  :  128 - 0x80
    "10000000", -- 2275 - 0x8e3  :  128 - 0x80
    "10011011", -- 2276 - 0x8e4  :  155 - 0x9b
    "10100100", -- 2277 - 0x8e5  :  164 - 0xa4
    "10100110", -- 2278 - 0x8e6  :  166 - 0xa6
    "10000000", -- 2279 - 0x8e7  :  128 - 0x80
    "10000000", -- 2280 - 0x8e8  :  128 - 0x80 -- Background 0x1d
    "01111111", -- 2281 - 0x8e9  :  127 - 0x7f
    "00000010", -- 2282 - 0x8ea  :    2 - 0x2
    "00000010", -- 2283 - 0x8eb  :    2 - 0x2
    "00000010", -- 2284 - 0x8ec  :    2 - 0x2
    "00000010", -- 2285 - 0x8ed  :    2 - 0x2
    "00000010", -- 2286 - 0x8ee  :    2 - 0x2
    "00001111", -- 2287 - 0x8ef  :   15 - 0xf
    "11111110", -- 2288 - 0x8f0  :  254 - 0xfe -- Background 0x1e
    "00000001", -- 2289 - 0x8f1  :    1 - 0x1
    "00000001", -- 2290 - 0x8f2  :    1 - 0x1
    "00000001", -- 2291 - 0x8f3  :    1 - 0x1
    "01000001", -- 2292 - 0x8f4  :   65 - 0x41
    "11110101", -- 2293 - 0x8f5  :  245 - 0xf5
    "00011101", -- 2294 - 0x8f6  :   29 - 0x1d
    "00000001", -- 2295 - 0x8f7  :    1 - 0x1
    "00000001", -- 2296 - 0x8f8  :    1 - 0x1 -- Background 0x1f
    "11111110", -- 2297 - 0x8f9  :  254 - 0xfe
    "01000000", -- 2298 - 0x8fa  :   64 - 0x40
    "01000000", -- 2299 - 0x8fb  :   64 - 0x40
    "01000000", -- 2300 - 0x8fc  :   64 - 0x40
    "01000000", -- 2301 - 0x8fd  :   64 - 0x40
    "01000000", -- 2302 - 0x8fe  :   64 - 0x40
    "11110000", -- 2303 - 0x8ff  :  240 - 0xf0
    "00000111", -- 2304 - 0x900  :    7 - 0x7 -- Background 0x20
    "00011111", -- 2305 - 0x901  :   31 - 0x1f
    "00111111", -- 2306 - 0x902  :   63 - 0x3f
    "01111111", -- 2307 - 0x903  :  127 - 0x7f
    "01111111", -- 2308 - 0x904  :  127 - 0x7f
    "11111111", -- 2309 - 0x905  :  255 - 0xff
    "11111111", -- 2310 - 0x906  :  255 - 0xff
    "11111111", -- 2311 - 0x907  :  255 - 0xff
    "11100000", -- 2312 - 0x908  :  224 - 0xe0 -- Background 0x21
    "11111000", -- 2313 - 0x909  :  248 - 0xf8
    "11111100", -- 2314 - 0x90a  :  252 - 0xfc
    "11111110", -- 2315 - 0x90b  :  254 - 0xfe
    "11111110", -- 2316 - 0x90c  :  254 - 0xfe
    "11111111", -- 2317 - 0x90d  :  255 - 0xff
    "11111111", -- 2318 - 0x90e  :  255 - 0xff
    "11111111", -- 2319 - 0x90f  :  255 - 0xff
    "00000111", -- 2320 - 0x910  :    7 - 0x7 -- Background 0x22
    "00011111", -- 2321 - 0x911  :   31 - 0x1f
    "00111111", -- 2322 - 0x912  :   63 - 0x3f
    "01111111", -- 2323 - 0x913  :  127 - 0x7f
    "01111111", -- 2324 - 0x914  :  127 - 0x7f
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "11111111", -- 2326 - 0x916  :  255 - 0xff
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "11100000", -- 2328 - 0x918  :  224 - 0xe0 -- Background 0x23
    "11111000", -- 2329 - 0x919  :  248 - 0xf8
    "11111100", -- 2330 - 0x91a  :  252 - 0xfc
    "11111110", -- 2331 - 0x91b  :  254 - 0xfe
    "11111110", -- 2332 - 0x91c  :  254 - 0xfe
    "11111111", -- 2333 - 0x91d  :  255 - 0xff
    "11111111", -- 2334 - 0x91e  :  255 - 0xff
    "11111111", -- 2335 - 0x91f  :  255 - 0xff
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Background 0x24
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00101111", -- 2344 - 0x928  :   47 - 0x2f -- Background 0x25
    "01001111", -- 2345 - 0x929  :   79 - 0x4f
    "01001111", -- 2346 - 0x92a  :   79 - 0x4f
    "01001111", -- 2347 - 0x92b  :   79 - 0x4f
    "01001111", -- 2348 - 0x92c  :   79 - 0x4f
    "00100111", -- 2349 - 0x92d  :   39 - 0x27
    "00010000", -- 2350 - 0x92e  :   16 - 0x10
    "00001111", -- 2351 - 0x92f  :   15 - 0xf
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "11100000", -- 2353 - 0x931  :  224 - 0xe0
    "10100000", -- 2354 - 0x932  :  160 - 0xa0
    "00100000", -- 2355 - 0x933  :   32 - 0x20
    "11000000", -- 2356 - 0x934  :  192 - 0xc0
    "01000000", -- 2357 - 0x935  :   64 - 0x40
    "00110000", -- 2358 - 0x936  :   48 - 0x30
    "11101000", -- 2359 - 0x937  :  232 - 0xe8
    "11110100", -- 2360 - 0x938  :  244 - 0xf4 -- Background 0x27
    "11110010", -- 2361 - 0x939  :  242 - 0xf2
    "11110010", -- 2362 - 0x93a  :  242 - 0xf2
    "11110010", -- 2363 - 0x93b  :  242 - 0xf2
    "11110010", -- 2364 - 0x93c  :  242 - 0xf2
    "11100100", -- 2365 - 0x93d  :  228 - 0xe4
    "00001000", -- 2366 - 0x93e  :    8 - 0x8
    "11110000", -- 2367 - 0x93f  :  240 - 0xf0
    "11111111", -- 2368 - 0x940  :  255 - 0xff -- Background 0x28
    "11010101", -- 2369 - 0x941  :  213 - 0xd5
    "10100011", -- 2370 - 0x942  :  163 - 0xa3
    "11010111", -- 2371 - 0x943  :  215 - 0xd7
    "10001111", -- 2372 - 0x944  :  143 - 0x8f
    "11001111", -- 2373 - 0x945  :  207 - 0xcf
    "10001011", -- 2374 - 0x946  :  139 - 0x8b
    "11001011", -- 2375 - 0x947  :  203 - 0xcb
    "10001111", -- 2376 - 0x948  :  143 - 0x8f -- Background 0x29
    "11001111", -- 2377 - 0x949  :  207 - 0xcf
    "10001111", -- 2378 - 0x94a  :  143 - 0x8f
    "11001111", -- 2379 - 0x94b  :  207 - 0xcf
    "10010000", -- 2380 - 0x94c  :  144 - 0x90
    "11100000", -- 2381 - 0x94d  :  224 - 0xe0
    "11101010", -- 2382 - 0x94e  :  234 - 0xea
    "11111111", -- 2383 - 0x94f  :  255 - 0xff
    "11111111", -- 2384 - 0x950  :  255 - 0xff -- Background 0x2a
    "11011011", -- 2385 - 0x951  :  219 - 0xdb
    "11000111", -- 2386 - 0x952  :  199 - 0xc7
    "11101001", -- 2387 - 0x953  :  233 - 0xe9
    "11110011", -- 2388 - 0x954  :  243 - 0xf3
    "11110001", -- 2389 - 0x955  :  241 - 0xf1
    "11010011", -- 2390 - 0x956  :  211 - 0xd3
    "11010001", -- 2391 - 0x957  :  209 - 0xd1
    "11110011", -- 2392 - 0x958  :  243 - 0xf3 -- Background 0x2b
    "11110001", -- 2393 - 0x959  :  241 - 0xf1
    "11110011", -- 2394 - 0x95a  :  243 - 0xf3
    "11110001", -- 2395 - 0x95b  :  241 - 0xf1
    "00001011", -- 2396 - 0x95c  :   11 - 0xb
    "00000101", -- 2397 - 0x95d  :    5 - 0x5
    "10101011", -- 2398 - 0x95e  :  171 - 0xab
    "11111111", -- 2399 - 0x95f  :  255 - 0xff
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00101111", -- 2408 - 0x968  :   47 - 0x2f -- Background 0x2d
    "01001111", -- 2409 - 0x969  :   79 - 0x4f
    "01001111", -- 2410 - 0x96a  :   79 - 0x4f
    "01001111", -- 2411 - 0x96b  :   79 - 0x4f
    "01001111", -- 2412 - 0x96c  :   79 - 0x4f
    "00100111", -- 2413 - 0x96d  :   39 - 0x27
    "00010000", -- 2414 - 0x96e  :   16 - 0x10
    "00001111", -- 2415 - 0x96f  :   15 - 0xf
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "11110100", -- 2424 - 0x978  :  244 - 0xf4 -- Background 0x2f
    "11110010", -- 2425 - 0x979  :  242 - 0xf2
    "11110010", -- 2426 - 0x97a  :  242 - 0xf2
    "11110010", -- 2427 - 0x97b  :  242 - 0xf2
    "11110010", -- 2428 - 0x97c  :  242 - 0xf2
    "11100100", -- 2429 - 0x97d  :  228 - 0xe4
    "00001000", -- 2430 - 0x97e  :    8 - 0x8
    "11110000", -- 2431 - 0x97f  :  240 - 0xf0
    "00011000", -- 2432 - 0x980  :   24 - 0x18 -- Background 0x30
    "00100100", -- 2433 - 0x981  :   36 - 0x24
    "01000010", -- 2434 - 0x982  :   66 - 0x42
    "10100101", -- 2435 - 0x983  :  165 - 0xa5
    "11100111", -- 2436 - 0x984  :  231 - 0xe7
    "00100100", -- 2437 - 0x985  :   36 - 0x24
    "00100100", -- 2438 - 0x986  :   36 - 0x24
    "00111100", -- 2439 - 0x987  :   60 - 0x3c
    "00111100", -- 2440 - 0x988  :   60 - 0x3c -- Background 0x31
    "00100100", -- 2441 - 0x989  :   36 - 0x24
    "00100100", -- 2442 - 0x98a  :   36 - 0x24
    "01100110", -- 2443 - 0x98b  :  102 - 0x66
    "10100101", -- 2444 - 0x98c  :  165 - 0xa5
    "01000010", -- 2445 - 0x98d  :   66 - 0x42
    "00100100", -- 2446 - 0x98e  :   36 - 0x24
    "00011000", -- 2447 - 0x98f  :   24 - 0x18
    "00000010", -- 2448 - 0x990  :    2 - 0x2 -- Background 0x32
    "00000010", -- 2449 - 0x991  :    2 - 0x2
    "00000011", -- 2450 - 0x992  :    3 - 0x3
    "00000010", -- 2451 - 0x993  :    2 - 0x2
    "00000010", -- 2452 - 0x994  :    2 - 0x2
    "00000010", -- 2453 - 0x995  :    2 - 0x2
    "00000011", -- 2454 - 0x996  :    3 - 0x3
    "00000010", -- 2455 - 0x997  :    2 - 0x2
    "01000000", -- 2456 - 0x998  :   64 - 0x40 -- Background 0x33
    "11000000", -- 2457 - 0x999  :  192 - 0xc0
    "01000000", -- 2458 - 0x99a  :   64 - 0x40
    "01000000", -- 2459 - 0x99b  :   64 - 0x40
    "01000000", -- 2460 - 0x99c  :   64 - 0x40
    "11000000", -- 2461 - 0x99d  :  192 - 0xc0
    "01000000", -- 2462 - 0x99e  :   64 - 0x40
    "01000000", -- 2463 - 0x99f  :   64 - 0x40
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Background 0x34
    "00011000", -- 2465 - 0x9a1  :   24 - 0x18
    "00111100", -- 2466 - 0x9a2  :   60 - 0x3c
    "01100010", -- 2467 - 0x9a3  :   98 - 0x62
    "01100001", -- 2468 - 0x9a4  :   97 - 0x61
    "11000000", -- 2469 - 0x9a5  :  192 - 0xc0
    "11000000", -- 2470 - 0x9a6  :  192 - 0xc0
    "11000000", -- 2471 - 0x9a7  :  192 - 0xc0
    "01100000", -- 2472 - 0x9a8  :   96 - 0x60 -- Background 0x35
    "01100000", -- 2473 - 0x9a9  :   96 - 0x60
    "00110000", -- 2474 - 0x9aa  :   48 - 0x30
    "00011000", -- 2475 - 0x9ab  :   24 - 0x18
    "00001100", -- 2476 - 0x9ac  :   12 - 0xc
    "00000110", -- 2477 - 0x9ad  :    6 - 0x6
    "00000010", -- 2478 - 0x9ae  :    2 - 0x2
    "00000001", -- 2479 - 0x9af  :    1 - 0x1
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0 -- Background 0x36
    "00011000", -- 2481 - 0x9b1  :   24 - 0x18
    "00100100", -- 2482 - 0x9b2  :   36 - 0x24
    "01000010", -- 2483 - 0x9b3  :   66 - 0x42
    "10000010", -- 2484 - 0x9b4  :  130 - 0x82
    "00000001", -- 2485 - 0x9b5  :    1 - 0x1
    "00000001", -- 2486 - 0x9b6  :    1 - 0x1
    "00000001", -- 2487 - 0x9b7  :    1 - 0x1
    "00000010", -- 2488 - 0x9b8  :    2 - 0x2 -- Background 0x37
    "00000010", -- 2489 - 0x9b9  :    2 - 0x2
    "00000100", -- 2490 - 0x9ba  :    4 - 0x4
    "00001000", -- 2491 - 0x9bb  :    8 - 0x8
    "00010000", -- 2492 - 0x9bc  :   16 - 0x10
    "00100000", -- 2493 - 0x9bd  :   32 - 0x20
    "01000000", -- 2494 - 0x9be  :   64 - 0x40
    "10000000", -- 2495 - 0x9bf  :  128 - 0x80
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000110", -- 2497 - 0x9c1  :    6 - 0x6
    "00001101", -- 2498 - 0x9c2  :   13 - 0xd
    "00001100", -- 2499 - 0x9c3  :   12 - 0xc
    "00001100", -- 2500 - 0x9c4  :   12 - 0xc
    "00000110", -- 2501 - 0x9c5  :    6 - 0x6
    "00000010", -- 2502 - 0x9c6  :    2 - 0x2
    "00000001", -- 2503 - 0x9c7  :    1 - 0x1
    "11111111", -- 2504 - 0x9c8  :  255 - 0xff -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "01100000", -- 2513 - 0x9d1  :   96 - 0x60
    "10010000", -- 2514 - 0x9d2  :  144 - 0x90
    "00010000", -- 2515 - 0x9d3  :   16 - 0x10
    "00010000", -- 2516 - 0x9d4  :   16 - 0x10
    "00100000", -- 2517 - 0x9d5  :   32 - 0x20
    "01000000", -- 2518 - 0x9d6  :   64 - 0x40
    "10000000", -- 2519 - 0x9d7  :  128 - 0x80
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "01010100", -- 2521 - 0x9d9  :   84 - 0x54
    "00000010", -- 2522 - 0x9da  :    2 - 0x2
    "01000000", -- 2523 - 0x9db  :   64 - 0x40
    "00000010", -- 2524 - 0x9dc  :    2 - 0x2
    "01000000", -- 2525 - 0x9dd  :   64 - 0x40
    "00101010", -- 2526 - 0x9de  :   42 - 0x2a
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "11111111", -- 2528 - 0x9e0  :  255 - 0xff -- Background 0x3c
    "11111111", -- 2529 - 0x9e1  :  255 - 0xff
    "11111111", -- 2530 - 0x9e2  :  255 - 0xff
    "11111111", -- 2531 - 0x9e3  :  255 - 0xff
    "11111111", -- 2532 - 0x9e4  :  255 - 0xff
    "11111111", -- 2533 - 0x9e5  :  255 - 0xff
    "11111111", -- 2534 - 0x9e6  :  255 - 0xff
    "11111111", -- 2535 - 0x9e7  :  255 - 0xff
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "11111111", -- 2544 - 0x9f0  :  255 - 0xff -- Background 0x3e
    "11111111", -- 2545 - 0x9f1  :  255 - 0xff
    "11111111", -- 2546 - 0x9f2  :  255 - 0xff
    "11111111", -- 2547 - 0x9f3  :  255 - 0xff
    "11111111", -- 2548 - 0x9f4  :  255 - 0xff
    "11111111", -- 2549 - 0x9f5  :  255 - 0xff
    "11111111", -- 2550 - 0x9f6  :  255 - 0xff
    "11111111", -- 2551 - 0x9f7  :  255 - 0xff
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00111100", -- 2560 - 0xa00  :   60 - 0x3c -- Background 0x40
    "01000010", -- 2561 - 0xa01  :   66 - 0x42
    "10011001", -- 2562 - 0xa02  :  153 - 0x99
    "10100101", -- 2563 - 0xa03  :  165 - 0xa5
    "10100101", -- 2564 - 0xa04  :  165 - 0xa5
    "10011010", -- 2565 - 0xa05  :  154 - 0x9a
    "01000000", -- 2566 - 0xa06  :   64 - 0x40
    "00111100", -- 2567 - 0xa07  :   60 - 0x3c
    "00001100", -- 2568 - 0xa08  :   12 - 0xc -- Background 0x41
    "00010010", -- 2569 - 0xa09  :   18 - 0x12
    "00100010", -- 2570 - 0xa0a  :   34 - 0x22
    "00100010", -- 2571 - 0xa0b  :   34 - 0x22
    "01111110", -- 2572 - 0xa0c  :  126 - 0x7e
    "00100010", -- 2573 - 0xa0d  :   34 - 0x22
    "00100100", -- 2574 - 0xa0e  :   36 - 0x24
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00111100", -- 2576 - 0xa10  :   60 - 0x3c -- Background 0x42
    "01000010", -- 2577 - 0xa11  :   66 - 0x42
    "01010010", -- 2578 - 0xa12  :   82 - 0x52
    "00011100", -- 2579 - 0xa13  :   28 - 0x1c
    "00010010", -- 2580 - 0xa14  :   18 - 0x12
    "00110010", -- 2581 - 0xa15  :   50 - 0x32
    "00011100", -- 2582 - 0xa16  :   28 - 0x1c
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00011000", -- 2584 - 0xa18  :   24 - 0x18 -- Background 0x43
    "00100100", -- 2585 - 0xa19  :   36 - 0x24
    "01010100", -- 2586 - 0xa1a  :   84 - 0x54
    "01001000", -- 2587 - 0xa1b  :   72 - 0x48
    "01000010", -- 2588 - 0xa1c  :   66 - 0x42
    "00100100", -- 2589 - 0xa1d  :   36 - 0x24
    "00011000", -- 2590 - 0xa1e  :   24 - 0x18
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "01011000", -- 2592 - 0xa20  :   88 - 0x58 -- Background 0x44
    "11100100", -- 2593 - 0xa21  :  228 - 0xe4
    "01000010", -- 2594 - 0xa22  :   66 - 0x42
    "01000010", -- 2595 - 0xa23  :   66 - 0x42
    "00100010", -- 2596 - 0xa24  :   34 - 0x22
    "01100100", -- 2597 - 0xa25  :  100 - 0x64
    "00111000", -- 2598 - 0xa26  :   56 - 0x38
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00011100", -- 2600 - 0xa28  :   28 - 0x1c -- Background 0x45
    "00100000", -- 2601 - 0xa29  :   32 - 0x20
    "00100000", -- 2602 - 0xa2a  :   32 - 0x20
    "00101100", -- 2603 - 0xa2b  :   44 - 0x2c
    "01110000", -- 2604 - 0xa2c  :  112 - 0x70
    "00100010", -- 2605 - 0xa2d  :   34 - 0x22
    "00011100", -- 2606 - 0xa2e  :   28 - 0x1c
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00011100", -- 2608 - 0xa30  :   28 - 0x1c -- Background 0x46
    "00100000", -- 2609 - 0xa31  :   32 - 0x20
    "00100000", -- 2610 - 0xa32  :   32 - 0x20
    "00101100", -- 2611 - 0xa33  :   44 - 0x2c
    "01110000", -- 2612 - 0xa34  :  112 - 0x70
    "00010000", -- 2613 - 0xa35  :   16 - 0x10
    "00010000", -- 2614 - 0xa36  :   16 - 0x10
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00011000", -- 2616 - 0xa38  :   24 - 0x18 -- Background 0x47
    "00100100", -- 2617 - 0xa39  :   36 - 0x24
    "01000000", -- 2618 - 0xa3a  :   64 - 0x40
    "01001110", -- 2619 - 0xa3b  :   78 - 0x4e
    "01000010", -- 2620 - 0xa3c  :   66 - 0x42
    "00100100", -- 2621 - 0xa3d  :   36 - 0x24
    "00011000", -- 2622 - 0xa3e  :   24 - 0x18
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00100000", -- 2624 - 0xa40  :   32 - 0x20 -- Background 0x48
    "01000100", -- 2625 - 0xa41  :   68 - 0x44
    "01000100", -- 2626 - 0xa42  :   68 - 0x44
    "01000100", -- 2627 - 0xa43  :   68 - 0x44
    "11111100", -- 2628 - 0xa44  :  252 - 0xfc
    "01000100", -- 2629 - 0xa45  :   68 - 0x44
    "01001000", -- 2630 - 0xa46  :   72 - 0x48
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00010000", -- 2632 - 0xa48  :   16 - 0x10 -- Background 0x49
    "00010000", -- 2633 - 0xa49  :   16 - 0x10
    "00010000", -- 2634 - 0xa4a  :   16 - 0x10
    "00010000", -- 2635 - 0xa4b  :   16 - 0x10
    "00010000", -- 2636 - 0xa4c  :   16 - 0x10
    "00001000", -- 2637 - 0xa4d  :    8 - 0x8
    "00001000", -- 2638 - 0xa4e  :    8 - 0x8
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00001000", -- 2640 - 0xa50  :    8 - 0x8 -- Background 0x4a
    "00001000", -- 2641 - 0xa51  :    8 - 0x8
    "00000100", -- 2642 - 0xa52  :    4 - 0x4
    "00000100", -- 2643 - 0xa53  :    4 - 0x4
    "01000100", -- 2644 - 0xa54  :   68 - 0x44
    "01001000", -- 2645 - 0xa55  :   72 - 0x48
    "00110000", -- 2646 - 0xa56  :   48 - 0x30
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "01000100", -- 2648 - 0xa58  :   68 - 0x44 -- Background 0x4b
    "01000100", -- 2649 - 0xa59  :   68 - 0x44
    "01001000", -- 2650 - 0xa5a  :   72 - 0x48
    "01110000", -- 2651 - 0xa5b  :  112 - 0x70
    "01001000", -- 2652 - 0xa5c  :   72 - 0x48
    "00100100", -- 2653 - 0xa5d  :   36 - 0x24
    "00100010", -- 2654 - 0xa5e  :   34 - 0x22
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00010000", -- 2656 - 0xa60  :   16 - 0x10 -- Background 0x4c
    "00100000", -- 2657 - 0xa61  :   32 - 0x20
    "00100000", -- 2658 - 0xa62  :   32 - 0x20
    "00100000", -- 2659 - 0xa63  :   32 - 0x20
    "01000000", -- 2660 - 0xa64  :   64 - 0x40
    "01000000", -- 2661 - 0xa65  :   64 - 0x40
    "01000110", -- 2662 - 0xa66  :   70 - 0x46
    "00111000", -- 2663 - 0xa67  :   56 - 0x38
    "00100100", -- 2664 - 0xa68  :   36 - 0x24 -- Background 0x4d
    "01011010", -- 2665 - 0xa69  :   90 - 0x5a
    "01011010", -- 2666 - 0xa6a  :   90 - 0x5a
    "01011010", -- 2667 - 0xa6b  :   90 - 0x5a
    "01000010", -- 2668 - 0xa6c  :   66 - 0x42
    "01000010", -- 2669 - 0xa6d  :   66 - 0x42
    "00100010", -- 2670 - 0xa6e  :   34 - 0x22
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00100100", -- 2672 - 0xa70  :   36 - 0x24 -- Background 0x4e
    "01010010", -- 2673 - 0xa71  :   82 - 0x52
    "01010010", -- 2674 - 0xa72  :   82 - 0x52
    "01010010", -- 2675 - 0xa73  :   82 - 0x52
    "01010010", -- 2676 - 0xa74  :   82 - 0x52
    "01010010", -- 2677 - 0xa75  :   82 - 0x52
    "01001100", -- 2678 - 0xa76  :   76 - 0x4c
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00111000", -- 2680 - 0xa78  :   56 - 0x38 -- Background 0x4f
    "01000100", -- 2681 - 0xa79  :   68 - 0x44
    "10000010", -- 2682 - 0xa7a  :  130 - 0x82
    "10000010", -- 2683 - 0xa7b  :  130 - 0x82
    "10000010", -- 2684 - 0xa7c  :  130 - 0x82
    "01000100", -- 2685 - 0xa7d  :   68 - 0x44
    "00111000", -- 2686 - 0xa7e  :   56 - 0x38
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "01111111", -- 2688 - 0xa80  :  127 - 0x7f -- Background 0x50
    "11000000", -- 2689 - 0xa81  :  192 - 0xc0
    "10000000", -- 2690 - 0xa82  :  128 - 0x80
    "10000000", -- 2691 - 0xa83  :  128 - 0x80
    "10000000", -- 2692 - 0xa84  :  128 - 0x80
    "11000011", -- 2693 - 0xa85  :  195 - 0xc3
    "11111111", -- 2694 - 0xa86  :  255 - 0xff
    "11111111", -- 2695 - 0xa87  :  255 - 0xff
    "11111110", -- 2696 - 0xa88  :  254 - 0xfe -- Background 0x51
    "00000011", -- 2697 - 0xa89  :    3 - 0x3
    "00000001", -- 2698 - 0xa8a  :    1 - 0x1
    "00000001", -- 2699 - 0xa8b  :    1 - 0x1
    "00000001", -- 2700 - 0xa8c  :    1 - 0x1
    "11000011", -- 2701 - 0xa8d  :  195 - 0xc3
    "11111111", -- 2702 - 0xa8e  :  255 - 0xff
    "11111111", -- 2703 - 0xa8f  :  255 - 0xff
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00000111", -- 2705 - 0xa91  :    7 - 0x7
    "00001100", -- 2706 - 0xa92  :   12 - 0xc
    "00011000", -- 2707 - 0xa93  :   24 - 0x18
    "00110000", -- 2708 - 0xa94  :   48 - 0x30
    "01100000", -- 2709 - 0xa95  :   96 - 0x60
    "01000000", -- 2710 - 0xa96  :   64 - 0x40
    "01001111", -- 2711 - 0xa97  :   79 - 0x4f
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- Background 0x53
    "11110000", -- 2713 - 0xa99  :  240 - 0xf0
    "01010000", -- 2714 - 0xa9a  :   80 - 0x50
    "01001000", -- 2715 - 0xa9b  :   72 - 0x48
    "01001100", -- 2716 - 0xa9c  :   76 - 0x4c
    "01000100", -- 2717 - 0xa9d  :   68 - 0x44
    "10000010", -- 2718 - 0xa9e  :  130 - 0x82
    "10000011", -- 2719 - 0xa9f  :  131 - 0x83
    "01111111", -- 2720 - 0xaa0  :  127 - 0x7f -- Background 0x54
    "11011110", -- 2721 - 0xaa1  :  222 - 0xde
    "10001110", -- 2722 - 0xaa2  :  142 - 0x8e
    "11000101", -- 2723 - 0xaa3  :  197 - 0xc5
    "10010010", -- 2724 - 0xaa4  :  146 - 0x92
    "11000111", -- 2725 - 0xaa5  :  199 - 0xc7
    "11100010", -- 2726 - 0xaa6  :  226 - 0xe2
    "11010000", -- 2727 - 0xaa7  :  208 - 0xd0
    "11111111", -- 2728 - 0xaa8  :  255 - 0xff -- Background 0x55
    "11011110", -- 2729 - 0xaa9  :  222 - 0xde
    "10001110", -- 2730 - 0xaaa  :  142 - 0x8e
    "11000101", -- 2731 - 0xaab  :  197 - 0xc5
    "10010010", -- 2732 - 0xaac  :  146 - 0x92
    "01000111", -- 2733 - 0xaad  :   71 - 0x47
    "11100010", -- 2734 - 0xaae  :  226 - 0xe2
    "01010000", -- 2735 - 0xaaf  :   80 - 0x50
    "11111110", -- 2736 - 0xab0  :  254 - 0xfe -- Background 0x56
    "11011111", -- 2737 - 0xab1  :  223 - 0xdf
    "10001111", -- 2738 - 0xab2  :  143 - 0x8f
    "11000101", -- 2739 - 0xab3  :  197 - 0xc5
    "10010011", -- 2740 - 0xab4  :  147 - 0x93
    "01000111", -- 2741 - 0xab5  :   71 - 0x47
    "11100011", -- 2742 - 0xab6  :  227 - 0xe3
    "01010001", -- 2743 - 0xab7  :   81 - 0x51
    "01111111", -- 2744 - 0xab8  :  127 - 0x7f -- Background 0x57
    "10000000", -- 2745 - 0xab9  :  128 - 0x80
    "10110011", -- 2746 - 0xaba  :  179 - 0xb3
    "01001100", -- 2747 - 0xabb  :   76 - 0x4c
    "00111111", -- 2748 - 0xabc  :   63 - 0x3f
    "00000011", -- 2749 - 0xabd  :    3 - 0x3
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "11111111", -- 2752 - 0xac0  :  255 - 0xff -- Background 0x58
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00110011", -- 2754 - 0xac2  :   51 - 0x33
    "11001100", -- 2755 - 0xac3  :  204 - 0xcc
    "00110011", -- 2756 - 0xac4  :   51 - 0x33
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "11111110", -- 2760 - 0xac8  :  254 - 0xfe -- Background 0x59
    "00000001", -- 2761 - 0xac9  :    1 - 0x1
    "00110011", -- 2762 - 0xaca  :   51 - 0x33
    "11001110", -- 2763 - 0xacb  :  206 - 0xce
    "00111100", -- 2764 - 0xacc  :   60 - 0x3c
    "11000000", -- 2765 - 0xacd  :  192 - 0xc0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "00000000", -- 2771 - 0xad3  :    0 - 0x0
    "00000000", -- 2772 - 0xad4  :    0 - 0x0
    "00000000", -- 2773 - 0xad5  :    0 - 0x0
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000001", -- 2779 - 0xadb  :    1 - 0x1
    "00000011", -- 2780 - 0xadc  :    3 - 0x3
    "00000011", -- 2781 - 0xadd  :    3 - 0x3
    "00000111", -- 2782 - 0xade  :    7 - 0x7
    "00111111", -- 2783 - 0xadf  :   63 - 0x3f
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Background 0x5c
    "00000001", -- 2785 - 0xae1  :    1 - 0x1
    "01111111", -- 2786 - 0xae2  :  127 - 0x7f
    "11111111", -- 2787 - 0xae3  :  255 - 0xff
    "11111111", -- 2788 - 0xae4  :  255 - 0xff
    "11111111", -- 2789 - 0xae5  :  255 - 0xff
    "11111111", -- 2790 - 0xae6  :  255 - 0xff
    "11111111", -- 2791 - 0xae7  :  255 - 0xff
    "11111111", -- 2792 - 0xae8  :  255 - 0xff -- Background 0x5d
    "11111111", -- 2793 - 0xae9  :  255 - 0xff
    "11111111", -- 2794 - 0xaea  :  255 - 0xff
    "11111111", -- 2795 - 0xaeb  :  255 - 0xff
    "11111111", -- 2796 - 0xaec  :  255 - 0xff
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "11111111", -- 2798 - 0xaee  :  255 - 0xff
    "11111111", -- 2799 - 0xaef  :  255 - 0xff
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0x5e
    "10000000", -- 2801 - 0xaf1  :  128 - 0x80
    "11111110", -- 2802 - 0xaf2  :  254 - 0xfe
    "11111111", -- 2803 - 0xaf3  :  255 - 0xff
    "11111111", -- 2804 - 0xaf4  :  255 - 0xff
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111111", -- 2806 - 0xaf6  :  255 - 0xff
    "11111111", -- 2807 - 0xaf7  :  255 - 0xff
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "10000000", -- 2811 - 0xafb  :  128 - 0x80
    "11000000", -- 2812 - 0xafc  :  192 - 0xc0
    "11000000", -- 2813 - 0xafd  :  192 - 0xc0
    "11100000", -- 2814 - 0xafe  :  224 - 0xe0
    "11111000", -- 2815 - 0xaff  :  248 - 0xf8
    "11111111", -- 2816 - 0xb00  :  255 - 0xff -- Background 0x60
    "11111111", -- 2817 - 0xb01  :  255 - 0xff
    "11111111", -- 2818 - 0xb02  :  255 - 0xff
    "11111111", -- 2819 - 0xb03  :  255 - 0xff
    "11111111", -- 2820 - 0xb04  :  255 - 0xff
    "11111111", -- 2821 - 0xb05  :  255 - 0xff
    "11111111", -- 2822 - 0xb06  :  255 - 0xff
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "11111111", -- 2824 - 0xb08  :  255 - 0xff -- Background 0x61
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11111111", -- 2826 - 0xb0a  :  255 - 0xff
    "11111111", -- 2827 - 0xb0b  :  255 - 0xff
    "11111111", -- 2828 - 0xb0c  :  255 - 0xff
    "11111111", -- 2829 - 0xb0d  :  255 - 0xff
    "11111111", -- 2830 - 0xb0e  :  255 - 0xff
    "11111111", -- 2831 - 0xb0f  :  255 - 0xff
    "01111000", -- 2832 - 0xb10  :  120 - 0x78 -- Background 0x62
    "01100000", -- 2833 - 0xb11  :   96 - 0x60
    "01000000", -- 2834 - 0xb12  :   64 - 0x40
    "01000000", -- 2835 - 0xb13  :   64 - 0x40
    "01000000", -- 2836 - 0xb14  :   64 - 0x40
    "01100000", -- 2837 - 0xb15  :   96 - 0x60
    "00110000", -- 2838 - 0xb16  :   48 - 0x30
    "00011111", -- 2839 - 0xb17  :   31 - 0x1f
    "10000001", -- 2840 - 0xb18  :  129 - 0x81 -- Background 0x63
    "10000011", -- 2841 - 0xb19  :  131 - 0x83
    "11000001", -- 2842 - 0xb1a  :  193 - 0xc1
    "01000011", -- 2843 - 0xb1b  :   67 - 0x43
    "01000001", -- 2844 - 0xb1c  :   65 - 0x41
    "01100011", -- 2845 - 0xb1d  :   99 - 0x63
    "00100110", -- 2846 - 0xb1e  :   38 - 0x26
    "11111000", -- 2847 - 0xb1f  :  248 - 0xf8
    "10111001", -- 2848 - 0xb20  :  185 - 0xb9 -- Background 0x64
    "10010100", -- 2849 - 0xb21  :  148 - 0x94
    "10001110", -- 2850 - 0xb22  :  142 - 0x8e
    "11000101", -- 2851 - 0xb23  :  197 - 0xc5
    "10010010", -- 2852 - 0xb24  :  146 - 0x92
    "11000111", -- 2853 - 0xb25  :  199 - 0xc7
    "11100010", -- 2854 - 0xb26  :  226 - 0xe2
    "11010000", -- 2855 - 0xb27  :  208 - 0xd0
    "10111001", -- 2856 - 0xb28  :  185 - 0xb9 -- Background 0x65
    "00010100", -- 2857 - 0xb29  :   20 - 0x14
    "10001110", -- 2858 - 0xb2a  :  142 - 0x8e
    "11000101", -- 2859 - 0xb2b  :  197 - 0xc5
    "10010010", -- 2860 - 0xb2c  :  146 - 0x92
    "01000111", -- 2861 - 0xb2d  :   71 - 0x47
    "11100010", -- 2862 - 0xb2e  :  226 - 0xe2
    "01010000", -- 2863 - 0xb2f  :   80 - 0x50
    "10111001", -- 2864 - 0xb30  :  185 - 0xb9 -- Background 0x66
    "00010101", -- 2865 - 0xb31  :   21 - 0x15
    "10001111", -- 2866 - 0xb32  :  143 - 0x8f
    "11000101", -- 2867 - 0xb33  :  197 - 0xc5
    "10010011", -- 2868 - 0xb34  :  147 - 0x93
    "01000111", -- 2869 - 0xb35  :   71 - 0x47
    "11100011", -- 2870 - 0xb36  :  227 - 0xe3
    "01010001", -- 2871 - 0xb37  :   81 - 0x51
    "01111111", -- 2872 - 0xb38  :  127 - 0x7f -- Background 0x67
    "10000000", -- 2873 - 0xb39  :  128 - 0x80
    "11001100", -- 2874 - 0xb3a  :  204 - 0xcc
    "01111111", -- 2875 - 0xb3b  :  127 - 0x7f
    "00111111", -- 2876 - 0xb3c  :   63 - 0x3f
    "00000011", -- 2877 - 0xb3d  :    3 - 0x3
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "11111111", -- 2880 - 0xb40  :  255 - 0xff -- Background 0x68
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "11001100", -- 2882 - 0xb42  :  204 - 0xcc
    "00110011", -- 2883 - 0xb43  :   51 - 0x33
    "11111111", -- 2884 - 0xb44  :  255 - 0xff
    "11111111", -- 2885 - 0xb45  :  255 - 0xff
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "11111110", -- 2888 - 0xb48  :  254 - 0xfe -- Background 0x69
    "00000001", -- 2889 - 0xb49  :    1 - 0x1
    "11001101", -- 2890 - 0xb4a  :  205 - 0xcd
    "00111110", -- 2891 - 0xb4b  :   62 - 0x3e
    "11111100", -- 2892 - 0xb4c  :  252 - 0xfc
    "11000000", -- 2893 - 0xb4d  :  192 - 0xc0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "01111111", -- 2904 - 0xb58  :  127 - 0x7f -- Background 0x6b
    "11111111", -- 2905 - 0xb59  :  255 - 0xff
    "11111111", -- 2906 - 0xb5a  :  255 - 0xff
    "11111111", -- 2907 - 0xb5b  :  255 - 0xff
    "01111111", -- 2908 - 0xb5c  :  127 - 0x7f
    "00110000", -- 2909 - 0xb5d  :   48 - 0x30
    "00001111", -- 2910 - 0xb5e  :   15 - 0xf
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Background 0x6c
    "11111111", -- 2913 - 0xb61  :  255 - 0xff
    "11111111", -- 2914 - 0xb62  :  255 - 0xff
    "11111111", -- 2915 - 0xb63  :  255 - 0xff
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11111110", -- 2917 - 0xb65  :  254 - 0xfe
    "00000001", -- 2918 - 0xb66  :    1 - 0x1
    "11111110", -- 2919 - 0xb67  :  254 - 0xfe
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "11111100", -- 2936 - 0xb78  :  252 - 0xfc -- Background 0x6f
    "11111110", -- 2937 - 0xb79  :  254 - 0xfe
    "11111111", -- 2938 - 0xb7a  :  255 - 0xff
    "11111111", -- 2939 - 0xb7b  :  255 - 0xff
    "11110010", -- 2940 - 0xb7c  :  242 - 0xf2
    "00001100", -- 2941 - 0xb7d  :   12 - 0xc
    "11110000", -- 2942 - 0xb7e  :  240 - 0xf0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "01111111", -- 2944 - 0xb80  :  127 - 0x7f -- Background 0x70
    "11000000", -- 2945 - 0xb81  :  192 - 0xc0
    "10000000", -- 2946 - 0xb82  :  128 - 0x80
    "10000000", -- 2947 - 0xb83  :  128 - 0x80
    "11100011", -- 2948 - 0xb84  :  227 - 0xe3
    "11111111", -- 2949 - 0xb85  :  255 - 0xff
    "11111111", -- 2950 - 0xb86  :  255 - 0xff
    "11111111", -- 2951 - 0xb87  :  255 - 0xff
    "11111111", -- 2952 - 0xb88  :  255 - 0xff -- Background 0x71
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "11000011", -- 2957 - 0xb8d  :  195 - 0xc3
    "11111111", -- 2958 - 0xb8e  :  255 - 0xff
    "11111111", -- 2959 - 0xb8f  :  255 - 0xff
    "11111110", -- 2960 - 0xb90  :  254 - 0xfe -- Background 0x72
    "00000011", -- 2961 - 0xb91  :    3 - 0x3
    "00000001", -- 2962 - 0xb92  :    1 - 0x1
    "00000001", -- 2963 - 0xb93  :    1 - 0x1
    "11000111", -- 2964 - 0xb94  :  199 - 0xc7
    "11111111", -- 2965 - 0xb95  :  255 - 0xff
    "11111111", -- 2966 - 0xb96  :  255 - 0xff
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "11111111", -- 2968 - 0xb98  :  255 - 0xff -- Background 0x73
    "11111111", -- 2969 - 0xb99  :  255 - 0xff
    "11111111", -- 2970 - 0xb9a  :  255 - 0xff
    "11111111", -- 2971 - 0xb9b  :  255 - 0xff
    "11111111", -- 2972 - 0xb9c  :  255 - 0xff
    "11111111", -- 2973 - 0xb9d  :  255 - 0xff
    "11111111", -- 2974 - 0xb9e  :  255 - 0xff
    "11111111", -- 2975 - 0xb9f  :  255 - 0xff
    "10111001", -- 2976 - 0xba0  :  185 - 0xb9 -- Background 0x74
    "10010100", -- 2977 - 0xba1  :  148 - 0x94
    "10001110", -- 2978 - 0xba2  :  142 - 0x8e
    "11000101", -- 2979 - 0xba3  :  197 - 0xc5
    "10010010", -- 2980 - 0xba4  :  146 - 0x92
    "11000111", -- 2981 - 0xba5  :  199 - 0xc7
    "11100010", -- 2982 - 0xba6  :  226 - 0xe2
    "01111111", -- 2983 - 0xba7  :  127 - 0x7f
    "10111001", -- 2984 - 0xba8  :  185 - 0xb9 -- Background 0x75
    "00010100", -- 2985 - 0xba9  :   20 - 0x14
    "10001110", -- 2986 - 0xbaa  :  142 - 0x8e
    "11000101", -- 2987 - 0xbab  :  197 - 0xc5
    "10010010", -- 2988 - 0xbac  :  146 - 0x92
    "01000111", -- 2989 - 0xbad  :   71 - 0x47
    "11100010", -- 2990 - 0xbae  :  226 - 0xe2
    "11111111", -- 2991 - 0xbaf  :  255 - 0xff
    "10111001", -- 2992 - 0xbb0  :  185 - 0xb9 -- Background 0x76
    "00010101", -- 2993 - 0xbb1  :   21 - 0x15
    "10001111", -- 2994 - 0xbb2  :  143 - 0x8f
    "11000101", -- 2995 - 0xbb3  :  197 - 0xc5
    "10010011", -- 2996 - 0xbb4  :  147 - 0x93
    "01000111", -- 2997 - 0xbb5  :   71 - 0x47
    "11100011", -- 2998 - 0xbb6  :  227 - 0xe3
    "11111110", -- 2999 - 0xbb7  :  254 - 0xfe
    "11111111", -- 3000 - 0xbb8  :  255 - 0xff -- Background 0x77
    "11111111", -- 3001 - 0xbb9  :  255 - 0xff
    "11111111", -- 3002 - 0xbba  :  255 - 0xff
    "11111111", -- 3003 - 0xbbb  :  255 - 0xff
    "11111111", -- 3004 - 0xbbc  :  255 - 0xff
    "11111111", -- 3005 - 0xbbd  :  255 - 0xff
    "11111111", -- 3006 - 0xbbe  :  255 - 0xff
    "11111111", -- 3007 - 0xbbf  :  255 - 0xff
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- Background 0x79
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00100010", -- 3040 - 0xbe0  :   34 - 0x22 -- Background 0x7c
    "01010101", -- 3041 - 0xbe1  :   85 - 0x55
    "10101010", -- 3042 - 0xbe2  :  170 - 0xaa
    "00000101", -- 3043 - 0xbe3  :    5 - 0x5
    "00000100", -- 3044 - 0xbe4  :    4 - 0x4
    "00001010", -- 3045 - 0xbe5  :   10 - 0xa
    "01010000", -- 3046 - 0xbe6  :   80 - 0x50
    "00000010", -- 3047 - 0xbe7  :    2 - 0x2
    "01110011", -- 3048 - 0xbe8  :  115 - 0x73 -- Background 0x7d
    "11111111", -- 3049 - 0xbe9  :  255 - 0xff
    "11111111", -- 3050 - 0xbea  :  255 - 0xff
    "10111101", -- 3051 - 0xbeb  :  189 - 0xbd
    "01101110", -- 3052 - 0xbec  :  110 - 0x6e
    "00001010", -- 3053 - 0xbed  :   10 - 0xa
    "01010000", -- 3054 - 0xbee  :   80 - 0x50
    "00000010", -- 3055 - 0xbef  :    2 - 0x2
    "00100000", -- 3056 - 0xbf0  :   32 - 0x20 -- Background 0x7e
    "01010000", -- 3057 - 0xbf1  :   80 - 0x50
    "10000100", -- 3058 - 0xbf2  :  132 - 0x84
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00100100", -- 3060 - 0xbf4  :   36 - 0x24
    "01011010", -- 3061 - 0xbf5  :   90 - 0x5a
    "00010000", -- 3062 - 0xbf6  :   16 - 0x10
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "11111111", -- 3064 - 0xbf8  :  255 - 0xff -- Background 0x7f
    "01010000", -- 3065 - 0xbf9  :   80 - 0x50
    "10000100", -- 3066 - 0xbfa  :  132 - 0x84
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00100100", -- 3068 - 0xbfc  :   36 - 0x24
    "01011010", -- 3069 - 0xbfd  :   90 - 0x5a
    "00010000", -- 3070 - 0xbfe  :   16 - 0x10
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "11111111", -- 3072 - 0xc00  :  255 - 0xff -- Background 0x80
    "10000000", -- 3073 - 0xc01  :  128 - 0x80
    "11001111", -- 3074 - 0xc02  :  207 - 0xcf
    "01001000", -- 3075 - 0xc03  :   72 - 0x48
    "11001111", -- 3076 - 0xc04  :  207 - 0xcf
    "10000000", -- 3077 - 0xc05  :  128 - 0x80
    "11001111", -- 3078 - 0xc06  :  207 - 0xcf
    "01001000", -- 3079 - 0xc07  :   72 - 0x48
    "11111111", -- 3080 - 0xc08  :  255 - 0xff -- Background 0x81
    "10000000", -- 3081 - 0xc09  :  128 - 0x80
    "11111111", -- 3082 - 0xc0a  :  255 - 0xff
    "10000000", -- 3083 - 0xc0b  :  128 - 0x80
    "10000000", -- 3084 - 0xc0c  :  128 - 0x80
    "11011111", -- 3085 - 0xc0d  :  223 - 0xdf
    "10110000", -- 3086 - 0xc0e  :  176 - 0xb0
    "11000000", -- 3087 - 0xc0f  :  192 - 0xc0
    "11111111", -- 3088 - 0xc10  :  255 - 0xff -- Background 0x82
    "00000001", -- 3089 - 0xc11  :    1 - 0x1
    "11110011", -- 3090 - 0xc12  :  243 - 0xf3
    "00010010", -- 3091 - 0xc13  :   18 - 0x12
    "11110011", -- 3092 - 0xc14  :  243 - 0xf3
    "00000001", -- 3093 - 0xc15  :    1 - 0x1
    "11110011", -- 3094 - 0xc16  :  243 - 0xf3
    "00010010", -- 3095 - 0xc17  :   18 - 0x12
    "11111111", -- 3096 - 0xc18  :  255 - 0xff -- Background 0x83
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "11111111", -- 3098 - 0xc1a  :  255 - 0xff
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "11111111", -- 3101 - 0xc1d  :  255 - 0xff
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "11111111", -- 3104 - 0xc20  :  255 - 0xff -- Background 0x84
    "10000010", -- 3105 - 0xc21  :  130 - 0x82
    "00010000", -- 3106 - 0xc22  :   16 - 0x10
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00010000", -- 3109 - 0xc25  :   16 - 0x10
    "01000100", -- 3110 - 0xc26  :   68 - 0x44
    "11111111", -- 3111 - 0xc27  :  255 - 0xff
    "11111111", -- 3112 - 0xc28  :  255 - 0xff -- Background 0x85
    "00000001", -- 3113 - 0xc29  :    1 - 0x1
    "11111111", -- 3114 - 0xc2a  :  255 - 0xff
    "00000001", -- 3115 - 0xc2b  :    1 - 0x1
    "00000001", -- 3116 - 0xc2c  :    1 - 0x1
    "11110011", -- 3117 - 0xc2d  :  243 - 0xf3
    "00001101", -- 3118 - 0xc2e  :   13 - 0xd
    "00000011", -- 3119 - 0xc2f  :    3 - 0x3
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0x86
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "00000000", -- 3126 - 0xc36  :    0 - 0x0
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- Background 0x87
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000111", -- 3136 - 0xc40  :    7 - 0x7 -- Background 0x88
    "00011110", -- 3137 - 0xc41  :   30 - 0x1e
    "00101111", -- 3138 - 0xc42  :   47 - 0x2f
    "01010011", -- 3139 - 0xc43  :   83 - 0x53
    "01101110", -- 3140 - 0xc44  :  110 - 0x6e
    "11011011", -- 3141 - 0xc45  :  219 - 0xdb
    "11111010", -- 3142 - 0xc46  :  250 - 0xfa
    "11010101", -- 3143 - 0xc47  :  213 - 0xd5
    "10111011", -- 3144 - 0xc48  :  187 - 0xbb -- Background 0x89
    "11110010", -- 3145 - 0xc49  :  242 - 0xf2
    "11011101", -- 3146 - 0xc4a  :  221 - 0xdd
    "01001111", -- 3147 - 0xc4b  :   79 - 0x4f
    "01111011", -- 3148 - 0xc4c  :  123 - 0x7b
    "00110010", -- 3149 - 0xc4d  :   50 - 0x32
    "00011111", -- 3150 - 0xc4e  :   31 - 0x1f
    "00000111", -- 3151 - 0xc4f  :    7 - 0x7
    "11100000", -- 3152 - 0xc50  :  224 - 0xe0 -- Background 0x8a
    "11011000", -- 3153 - 0xc51  :  216 - 0xd8
    "01010100", -- 3154 - 0xc52  :   84 - 0x54
    "11101010", -- 3155 - 0xc53  :  234 - 0xea
    "10111010", -- 3156 - 0xc54  :  186 - 0xba
    "10010011", -- 3157 - 0xc55  :  147 - 0x93
    "11011111", -- 3158 - 0xc56  :  223 - 0xdf
    "10111101", -- 3159 - 0xc57  :  189 - 0xbd
    "01101011", -- 3160 - 0xc58  :  107 - 0x6b -- Background 0x8b
    "10011111", -- 3161 - 0xc59  :  159 - 0x9f
    "01011101", -- 3162 - 0xc5a  :   93 - 0x5d
    "10110110", -- 3163 - 0xc5b  :  182 - 0xb6
    "11101010", -- 3164 - 0xc5c  :  234 - 0xea
    "11001100", -- 3165 - 0xc5d  :  204 - 0xcc
    "01111000", -- 3166 - 0xc5e  :  120 - 0x78
    "11100000", -- 3167 - 0xc5f  :  224 - 0xe0
    "00000111", -- 3168 - 0xc60  :    7 - 0x7 -- Background 0x8c
    "00011000", -- 3169 - 0xc61  :   24 - 0x18
    "00100011", -- 3170 - 0xc62  :   35 - 0x23
    "01001100", -- 3171 - 0xc63  :   76 - 0x4c
    "01110000", -- 3172 - 0xc64  :  112 - 0x70
    "10100001", -- 3173 - 0xc65  :  161 - 0xa1
    "10100110", -- 3174 - 0xc66  :  166 - 0xa6
    "10101000", -- 3175 - 0xc67  :  168 - 0xa8
    "10100101", -- 3176 - 0xc68  :  165 - 0xa5 -- Background 0x8d
    "10100010", -- 3177 - 0xc69  :  162 - 0xa2
    "10010000", -- 3178 - 0xc6a  :  144 - 0x90
    "01001000", -- 3179 - 0xc6b  :   72 - 0x48
    "01000111", -- 3180 - 0xc6c  :   71 - 0x47
    "00100000", -- 3181 - 0xc6d  :   32 - 0x20
    "00011001", -- 3182 - 0xc6e  :   25 - 0x19
    "00000111", -- 3183 - 0xc6f  :    7 - 0x7
    "11100000", -- 3184 - 0xc70  :  224 - 0xe0 -- Background 0x8e
    "00011000", -- 3185 - 0xc71  :   24 - 0x18
    "00000100", -- 3186 - 0xc72  :    4 - 0x4
    "11000010", -- 3187 - 0xc73  :  194 - 0xc2
    "00110010", -- 3188 - 0xc74  :   50 - 0x32
    "00001001", -- 3189 - 0xc75  :    9 - 0x9
    "11000101", -- 3190 - 0xc76  :  197 - 0xc5
    "00100101", -- 3191 - 0xc77  :   37 - 0x25
    "10100101", -- 3192 - 0xc78  :  165 - 0xa5 -- Background 0x8f
    "01100101", -- 3193 - 0xc79  :  101 - 0x65
    "01000101", -- 3194 - 0xc7a  :   69 - 0x45
    "10001010", -- 3195 - 0xc7b  :  138 - 0x8a
    "10010010", -- 3196 - 0xc7c  :  146 - 0x92
    "00100100", -- 3197 - 0xc7d  :   36 - 0x24
    "11011000", -- 3198 - 0xc7e  :  216 - 0xd8
    "11100000", -- 3199 - 0xc7f  :  224 - 0xe0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00100000", -- 3202 - 0xc82  :   32 - 0x20
    "00110000", -- 3203 - 0xc83  :   48 - 0x30
    "00101100", -- 3204 - 0xc84  :   44 - 0x2c
    "00100010", -- 3205 - 0xc85  :   34 - 0x22
    "00010001", -- 3206 - 0xc86  :   17 - 0x11
    "00001000", -- 3207 - 0xc87  :    8 - 0x8
    "00000100", -- 3208 - 0xc88  :    4 - 0x4 -- Background 0x91
    "11110010", -- 3209 - 0xc89  :  242 - 0xf2
    "11001111", -- 3210 - 0xc8a  :  207 - 0xcf
    "00110000", -- 3211 - 0xc8b  :   48 - 0x30
    "00001100", -- 3212 - 0xc8c  :   12 - 0xc
    "11111111", -- 3213 - 0xc8d  :  255 - 0xff
    "10000000", -- 3214 - 0xc8e  :  128 - 0x80
    "11111111", -- 3215 - 0xc8f  :  255 - 0xff
    "01000010", -- 3216 - 0xc90  :   66 - 0x42 -- Background 0x92
    "10100101", -- 3217 - 0xc91  :  165 - 0xa5
    "10100101", -- 3218 - 0xc92  :  165 - 0xa5
    "10011001", -- 3219 - 0xc93  :  153 - 0x99
    "10011001", -- 3220 - 0xc94  :  153 - 0x99
    "10011001", -- 3221 - 0xc95  :  153 - 0x99
    "00000001", -- 3222 - 0xc96  :    1 - 0x1
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "11111111", -- 3224 - 0xc98  :  255 - 0xff -- Background 0x93
    "11111111", -- 3225 - 0xc99  :  255 - 0xff
    "11111111", -- 3226 - 0xc9a  :  255 - 0xff
    "10000001", -- 3227 - 0xc9b  :  129 - 0x81
    "11111111", -- 3228 - 0xc9c  :  255 - 0xff
    "11111111", -- 3229 - 0xc9d  :  255 - 0xff
    "11111111", -- 3230 - 0xc9e  :  255 - 0xff
    "10000001", -- 3231 - 0xc9f  :  129 - 0x81
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000100", -- 3234 - 0xca2  :    4 - 0x4
    "00001100", -- 3235 - 0xca3  :   12 - 0xc
    "00110100", -- 3236 - 0xca4  :   52 - 0x34
    "01000100", -- 3237 - 0xca5  :   68 - 0x44
    "10001000", -- 3238 - 0xca6  :  136 - 0x88
    "00010000", -- 3239 - 0xca7  :   16 - 0x10
    "00100000", -- 3240 - 0xca8  :   32 - 0x20 -- Background 0x95
    "01001111", -- 3241 - 0xca9  :   79 - 0x4f
    "11110011", -- 3242 - 0xcaa  :  243 - 0xf3
    "00001100", -- 3243 - 0xcab  :   12 - 0xc
    "00110000", -- 3244 - 0xcac  :   48 - 0x30
    "11111111", -- 3245 - 0xcad  :  255 - 0xff
    "00000001", -- 3246 - 0xcae  :    1 - 0x1
    "11111111", -- 3247 - 0xcaf  :  255 - 0xff
    "01111111", -- 3248 - 0xcb0  :  127 - 0x7f -- Background 0x96
    "11111111", -- 3249 - 0xcb1  :  255 - 0xff
    "11111111", -- 3250 - 0xcb2  :  255 - 0xff
    "11111111", -- 3251 - 0xcb3  :  255 - 0xff
    "11111011", -- 3252 - 0xcb4  :  251 - 0xfb
    "11111111", -- 3253 - 0xcb5  :  255 - 0xff
    "11111111", -- 3254 - 0xcb6  :  255 - 0xff
    "11111111", -- 3255 - 0xcb7  :  255 - 0xff
    "11111111", -- 3256 - 0xcb8  :  255 - 0xff -- Background 0x97
    "11111111", -- 3257 - 0xcb9  :  255 - 0xff
    "11111111", -- 3258 - 0xcba  :  255 - 0xff
    "11111111", -- 3259 - 0xcbb  :  255 - 0xff
    "11111111", -- 3260 - 0xcbc  :  255 - 0xff
    "11111111", -- 3261 - 0xcbd  :  255 - 0xff
    "11111110", -- 3262 - 0xcbe  :  254 - 0xfe
    "11111111", -- 3263 - 0xcbf  :  255 - 0xff
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff -- Background 0x98
    "10111111", -- 3265 - 0xcc1  :  191 - 0xbf
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111111", -- 3267 - 0xcc3  :  255 - 0xff
    "11111011", -- 3268 - 0xcc4  :  251 - 0xfb
    "11111111", -- 3269 - 0xcc5  :  255 - 0xff
    "11111111", -- 3270 - 0xcc6  :  255 - 0xff
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "11111111", -- 3272 - 0xcc8  :  255 - 0xff -- Background 0x99
    "11111111", -- 3273 - 0xcc9  :  255 - 0xff
    "11111111", -- 3274 - 0xcca  :  255 - 0xff
    "11111111", -- 3275 - 0xccb  :  255 - 0xff
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "11111111", -- 3277 - 0xccd  :  255 - 0xff
    "11111110", -- 3278 - 0xcce  :  254 - 0xfe
    "11111111", -- 3279 - 0xccf  :  255 - 0xff
    "11111110", -- 3280 - 0xcd0  :  254 - 0xfe -- Background 0x9a
    "11111111", -- 3281 - 0xcd1  :  255 - 0xff
    "11111111", -- 3282 - 0xcd2  :  255 - 0xff
    "11111111", -- 3283 - 0xcd3  :  255 - 0xff
    "11111011", -- 3284 - 0xcd4  :  251 - 0xfb
    "11111111", -- 3285 - 0xcd5  :  255 - 0xff
    "11111111", -- 3286 - 0xcd6  :  255 - 0xff
    "11111111", -- 3287 - 0xcd7  :  255 - 0xff
    "11111111", -- 3288 - 0xcd8  :  255 - 0xff -- Background 0x9b
    "11111111", -- 3289 - 0xcd9  :  255 - 0xff
    "11111111", -- 3290 - 0xcda  :  255 - 0xff
    "11111111", -- 3291 - 0xcdb  :  255 - 0xff
    "11111111", -- 3292 - 0xcdc  :  255 - 0xff
    "11111111", -- 3293 - 0xcdd  :  255 - 0xff
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "11111111", -- 3296 - 0xce0  :  255 - 0xff -- Background 0x9c
    "11111111", -- 3297 - 0xce1  :  255 - 0xff
    "10100000", -- 3298 - 0xce2  :  160 - 0xa0
    "10010000", -- 3299 - 0xce3  :  144 - 0x90
    "10001000", -- 3300 - 0xce4  :  136 - 0x88
    "10000100", -- 3301 - 0xce5  :  132 - 0x84
    "01101010", -- 3302 - 0xce6  :  106 - 0x6a
    "00111111", -- 3303 - 0xce7  :   63 - 0x3f
    "11111111", -- 3304 - 0xce8  :  255 - 0xff -- Background 0x9d
    "11111111", -- 3305 - 0xce9  :  255 - 0xff
    "00100001", -- 3306 - 0xcea  :   33 - 0x21
    "00010001", -- 3307 - 0xceb  :   17 - 0x11
    "00001001", -- 3308 - 0xcec  :    9 - 0x9
    "00000101", -- 3309 - 0xced  :    5 - 0x5
    "10101010", -- 3310 - 0xcee  :  170 - 0xaa
    "11111100", -- 3311 - 0xcef  :  252 - 0xfc
    "11111111", -- 3312 - 0xcf0  :  255 - 0xff -- Background 0x9e
    "11111111", -- 3313 - 0xcf1  :  255 - 0xff
    "00100000", -- 3314 - 0xcf2  :   32 - 0x20
    "00010000", -- 3315 - 0xcf3  :   16 - 0x10
    "00001000", -- 3316 - 0xcf4  :    8 - 0x8
    "00000100", -- 3317 - 0xcf5  :    4 - 0x4
    "10101010", -- 3318 - 0xcf6  :  170 - 0xaa
    "11111111", -- 3319 - 0xcf7  :  255 - 0xff
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "11111111", -- 3328 - 0xd00  :  255 - 0xff -- Background 0xa0
    "11010101", -- 3329 - 0xd01  :  213 - 0xd5
    "11111111", -- 3330 - 0xd02  :  255 - 0xff
    "00000010", -- 3331 - 0xd03  :    2 - 0x2
    "00000010", -- 3332 - 0xd04  :    2 - 0x2
    "00000010", -- 3333 - 0xd05  :    2 - 0x2
    "00000010", -- 3334 - 0xd06  :    2 - 0x2
    "00000010", -- 3335 - 0xd07  :    2 - 0x2
    "00000010", -- 3336 - 0xd08  :    2 - 0x2 -- Background 0xa1
    "00000010", -- 3337 - 0xd09  :    2 - 0x2
    "00000010", -- 3338 - 0xd0a  :    2 - 0x2
    "00000010", -- 3339 - 0xd0b  :    2 - 0x2
    "00000010", -- 3340 - 0xd0c  :    2 - 0x2
    "00000010", -- 3341 - 0xd0d  :    2 - 0x2
    "00000010", -- 3342 - 0xd0e  :    2 - 0x2
    "00000010", -- 3343 - 0xd0f  :    2 - 0x2
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Background 0xa2
    "01010101", -- 3345 - 0xd11  :   85 - 0x55
    "11111111", -- 3346 - 0xd12  :  255 - 0xff
    "01000000", -- 3347 - 0xd13  :   64 - 0x40
    "01000000", -- 3348 - 0xd14  :   64 - 0x40
    "01000000", -- 3349 - 0xd15  :   64 - 0x40
    "01000000", -- 3350 - 0xd16  :   64 - 0x40
    "01000000", -- 3351 - 0xd17  :   64 - 0x40
    "01000000", -- 3352 - 0xd18  :   64 - 0x40 -- Background 0xa3
    "01000000", -- 3353 - 0xd19  :   64 - 0x40
    "01000000", -- 3354 - 0xd1a  :   64 - 0x40
    "01000000", -- 3355 - 0xd1b  :   64 - 0x40
    "01000000", -- 3356 - 0xd1c  :   64 - 0x40
    "01000000", -- 3357 - 0xd1d  :   64 - 0x40
    "01000000", -- 3358 - 0xd1e  :   64 - 0x40
    "01000000", -- 3359 - 0xd1f  :   64 - 0x40
    "00110001", -- 3360 - 0xd20  :   49 - 0x31 -- Background 0xa4
    "01001000", -- 3361 - 0xd21  :   72 - 0x48
    "01000101", -- 3362 - 0xd22  :   69 - 0x45
    "10000101", -- 3363 - 0xd23  :  133 - 0x85
    "10000011", -- 3364 - 0xd24  :  131 - 0x83
    "10000010", -- 3365 - 0xd25  :  130 - 0x82
    "01100010", -- 3366 - 0xd26  :   98 - 0x62
    "00010010", -- 3367 - 0xd27  :   18 - 0x12
    "00110010", -- 3368 - 0xd28  :   50 - 0x32 -- Background 0xa5
    "00100010", -- 3369 - 0xd29  :   34 - 0x22
    "01000010", -- 3370 - 0xd2a  :   66 - 0x42
    "01000000", -- 3371 - 0xd2b  :   64 - 0x40
    "01000000", -- 3372 - 0xd2c  :   64 - 0x40
    "00100000", -- 3373 - 0xd2d  :   32 - 0x20
    "00011110", -- 3374 - 0xd2e  :   30 - 0x1e
    "00000111", -- 3375 - 0xd2f  :    7 - 0x7
    "10000000", -- 3376 - 0xd30  :  128 - 0x80 -- Background 0xa6
    "11100000", -- 3377 - 0xd31  :  224 - 0xe0
    "00111000", -- 3378 - 0xd32  :   56 - 0x38
    "00100100", -- 3379 - 0xd33  :   36 - 0x24
    "00000100", -- 3380 - 0xd34  :    4 - 0x4
    "00001000", -- 3381 - 0xd35  :    8 - 0x8
    "00110000", -- 3382 - 0xd36  :   48 - 0x30
    "00100000", -- 3383 - 0xd37  :   32 - 0x20
    "00110000", -- 3384 - 0xd38  :   48 - 0x30 -- Background 0xa7
    "00001000", -- 3385 - 0xd39  :    8 - 0x8
    "00001000", -- 3386 - 0xd3a  :    8 - 0x8
    "00110000", -- 3387 - 0xd3b  :   48 - 0x30
    "00100000", -- 3388 - 0xd3c  :   32 - 0x20
    "00100000", -- 3389 - 0xd3d  :   32 - 0x20
    "00110000", -- 3390 - 0xd3e  :   48 - 0x30
    "11110000", -- 3391 - 0xd3f  :  240 - 0xf0
    "11111111", -- 3392 - 0xd40  :  255 - 0xff -- Background 0xa8
    "11010010", -- 3393 - 0xd41  :  210 - 0xd2
    "11110100", -- 3394 - 0xd42  :  244 - 0xf4
    "11011000", -- 3395 - 0xd43  :  216 - 0xd8
    "11111000", -- 3396 - 0xd44  :  248 - 0xf8
    "11010100", -- 3397 - 0xd45  :  212 - 0xd4
    "11110010", -- 3398 - 0xd46  :  242 - 0xf2
    "11010001", -- 3399 - 0xd47  :  209 - 0xd1
    "11110001", -- 3400 - 0xd48  :  241 - 0xf1 -- Background 0xa9
    "11010010", -- 3401 - 0xd49  :  210 - 0xd2
    "11110100", -- 3402 - 0xd4a  :  244 - 0xf4
    "11011000", -- 3403 - 0xd4b  :  216 - 0xd8
    "11111000", -- 3404 - 0xd4c  :  248 - 0xf8
    "11010100", -- 3405 - 0xd4d  :  212 - 0xd4
    "11110010", -- 3406 - 0xd4e  :  242 - 0xf2
    "11111111", -- 3407 - 0xd4f  :  255 - 0xff
    "11111111", -- 3408 - 0xd50  :  255 - 0xff -- Background 0xaa
    "01000010", -- 3409 - 0xd51  :   66 - 0x42
    "00100100", -- 3410 - 0xd52  :   36 - 0x24
    "00011000", -- 3411 - 0xd53  :   24 - 0x18
    "00011000", -- 3412 - 0xd54  :   24 - 0x18
    "00100100", -- 3413 - 0xd55  :   36 - 0x24
    "01000010", -- 3414 - 0xd56  :   66 - 0x42
    "10000001", -- 3415 - 0xd57  :  129 - 0x81
    "10000001", -- 3416 - 0xd58  :  129 - 0x81 -- Background 0xab
    "01000010", -- 3417 - 0xd59  :   66 - 0x42
    "00100100", -- 3418 - 0xd5a  :   36 - 0x24
    "00011000", -- 3419 - 0xd5b  :   24 - 0x18
    "00011000", -- 3420 - 0xd5c  :   24 - 0x18
    "00100100", -- 3421 - 0xd5d  :   36 - 0x24
    "01000010", -- 3422 - 0xd5e  :   66 - 0x42
    "11111111", -- 3423 - 0xd5f  :  255 - 0xff
    "11111111", -- 3424 - 0xd60  :  255 - 0xff -- Background 0xac
    "01001101", -- 3425 - 0xd61  :   77 - 0x4d
    "00101111", -- 3426 - 0xd62  :   47 - 0x2f
    "00011101", -- 3427 - 0xd63  :   29 - 0x1d
    "00011111", -- 3428 - 0xd64  :   31 - 0x1f
    "00101101", -- 3429 - 0xd65  :   45 - 0x2d
    "01001111", -- 3430 - 0xd66  :   79 - 0x4f
    "10001101", -- 3431 - 0xd67  :  141 - 0x8d
    "10001111", -- 3432 - 0xd68  :  143 - 0x8f -- Background 0xad
    "01001101", -- 3433 - 0xd69  :   77 - 0x4d
    "00101111", -- 3434 - 0xd6a  :   47 - 0x2f
    "00011101", -- 3435 - 0xd6b  :   29 - 0x1d
    "00011111", -- 3436 - 0xd6c  :   31 - 0x1f
    "00101101", -- 3437 - 0xd6d  :   45 - 0x2d
    "01001111", -- 3438 - 0xd6e  :   79 - 0x4f
    "11111111", -- 3439 - 0xd6f  :  255 - 0xff
    "00000001", -- 3440 - 0xd70  :    1 - 0x1 -- Background 0xae
    "00000011", -- 3441 - 0xd71  :    3 - 0x3
    "00000110", -- 3442 - 0xd72  :    6 - 0x6
    "00000111", -- 3443 - 0xd73  :    7 - 0x7
    "00000111", -- 3444 - 0xd74  :    7 - 0x7
    "00000111", -- 3445 - 0xd75  :    7 - 0x7
    "00000110", -- 3446 - 0xd76  :    6 - 0x6
    "00000111", -- 3447 - 0xd77  :    7 - 0x7
    "00000110", -- 3448 - 0xd78  :    6 - 0x6 -- Background 0xaf
    "00000110", -- 3449 - 0xd79  :    6 - 0x6
    "00001110", -- 3450 - 0xd7a  :   14 - 0xe
    "00001111", -- 3451 - 0xd7b  :   15 - 0xf
    "00001110", -- 3452 - 0xd7c  :   14 - 0xe
    "00011010", -- 3453 - 0xd7d  :   26 - 0x1a
    "00011011", -- 3454 - 0xd7e  :   27 - 0x1b
    "00001111", -- 3455 - 0xd7f  :   15 - 0xf
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xb0
    "11000000", -- 3457 - 0xd81  :  192 - 0xc0
    "11110000", -- 3458 - 0xd82  :  240 - 0xf0
    "10001000", -- 3459 - 0xd83  :  136 - 0x88
    "00010100", -- 3460 - 0xd84  :   20 - 0x14
    "01101000", -- 3461 - 0xd85  :  104 - 0x68
    "10101000", -- 3462 - 0xd86  :  168 - 0xa8
    "00101100", -- 3463 - 0xd87  :   44 - 0x2c
    "00000100", -- 3464 - 0xd88  :    4 - 0x4 -- Background 0xb1
    "00111000", -- 3465 - 0xd89  :   56 - 0x38
    "00010000", -- 3466 - 0xd8a  :   16 - 0x10
    "10100000", -- 3467 - 0xd8b  :  160 - 0xa0
    "01100000", -- 3468 - 0xd8c  :   96 - 0x60
    "00100000", -- 3469 - 0xd8d  :   32 - 0x20
    "00010000", -- 3470 - 0xd8e  :   16 - 0x10
    "10001000", -- 3471 - 0xd8f  :  136 - 0x88
    "00001111", -- 3472 - 0xd90  :   15 - 0xf -- Background 0xb2
    "00011011", -- 3473 - 0xd91  :   27 - 0x1b
    "00011011", -- 3474 - 0xd92  :   27 - 0x1b
    "00001110", -- 3475 - 0xd93  :   14 - 0xe
    "00000110", -- 3476 - 0xd94  :    6 - 0x6
    "00001100", -- 3477 - 0xd95  :   12 - 0xc
    "00001100", -- 3478 - 0xd96  :   12 - 0xc
    "00111111", -- 3479 - 0xd97  :   63 - 0x3f
    "01111111", -- 3480 - 0xd98  :  127 - 0x7f -- Background 0xb3
    "01100000", -- 3481 - 0xd99  :   96 - 0x60
    "01100000", -- 3482 - 0xd9a  :   96 - 0x60
    "01100000", -- 3483 - 0xd9b  :   96 - 0x60
    "01100000", -- 3484 - 0xd9c  :   96 - 0x60
    "01100000", -- 3485 - 0xd9d  :   96 - 0x60
    "01101010", -- 3486 - 0xd9e  :  106 - 0x6a
    "01111111", -- 3487 - 0xd9f  :  127 - 0x7f
    "01001000", -- 3488 - 0xda0  :   72 - 0x48 -- Background 0xb4
    "00110000", -- 3489 - 0xda1  :   48 - 0x30
    "00010000", -- 3490 - 0xda2  :   16 - 0x10
    "00010000", -- 3491 - 0xda3  :   16 - 0x10
    "00001000", -- 3492 - 0xda4  :    8 - 0x8
    "00001000", -- 3493 - 0xda5  :    8 - 0x8
    "00001000", -- 3494 - 0xda6  :    8 - 0x8
    "11111100", -- 3495 - 0xda7  :  252 - 0xfc
    "11111110", -- 3496 - 0xda8  :  254 - 0xfe -- Background 0xb5
    "00000110", -- 3497 - 0xda9  :    6 - 0x6
    "00000010", -- 3498 - 0xdaa  :    2 - 0x2
    "00000110", -- 3499 - 0xdab  :    6 - 0x6
    "00000010", -- 3500 - 0xdac  :    2 - 0x2
    "00000110", -- 3501 - 0xdad  :    6 - 0x6
    "10101010", -- 3502 - 0xdae  :  170 - 0xaa
    "11111110", -- 3503 - 0xdaf  :  254 - 0xfe
    "11111111", -- 3504 - 0xdb0  :  255 - 0xff -- Background 0xb6
    "10000000", -- 3505 - 0xdb1  :  128 - 0x80
    "10000000", -- 3506 - 0xdb2  :  128 - 0x80
    "10000000", -- 3507 - 0xdb3  :  128 - 0x80
    "10000000", -- 3508 - 0xdb4  :  128 - 0x80
    "10000000", -- 3509 - 0xdb5  :  128 - 0x80
    "10010101", -- 3510 - 0xdb6  :  149 - 0x95
    "11111111", -- 3511 - 0xdb7  :  255 - 0xff
    "11111111", -- 3512 - 0xdb8  :  255 - 0xff -- Background 0xb7
    "10000100", -- 3513 - 0xdb9  :  132 - 0x84
    "10001100", -- 3514 - 0xdba  :  140 - 0x8c
    "10000100", -- 3515 - 0xdbb  :  132 - 0x84
    "10001100", -- 3516 - 0xdbc  :  140 - 0x8c
    "10000100", -- 3517 - 0xdbd  :  132 - 0x84
    "10101100", -- 3518 - 0xdbe  :  172 - 0xac
    "11111111", -- 3519 - 0xdbf  :  255 - 0xff
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Background 0xb8
    "00100001", -- 3521 - 0xdc1  :   33 - 0x21
    "01100001", -- 3522 - 0xdc2  :   97 - 0x61
    "00100011", -- 3523 - 0xdc3  :   35 - 0x23
    "01100001", -- 3524 - 0xdc4  :   97 - 0x61
    "00100011", -- 3525 - 0xdc5  :   35 - 0x23
    "01100101", -- 3526 - 0xdc6  :  101 - 0x65
    "11111111", -- 3527 - 0xdc7  :  255 - 0xff
    "11111111", -- 3528 - 0xdc8  :  255 - 0xff -- Background 0xb9
    "00000001", -- 3529 - 0xdc9  :    1 - 0x1
    "00000011", -- 3530 - 0xdca  :    3 - 0x3
    "00000001", -- 3531 - 0xdcb  :    1 - 0x1
    "00000011", -- 3532 - 0xdcc  :    3 - 0x3
    "00000001", -- 3533 - 0xdcd  :    1 - 0x1
    "10101011", -- 3534 - 0xdce  :  171 - 0xab
    "11111111", -- 3535 - 0xdcf  :  255 - 0xff
    "11111111", -- 3536 - 0xdd0  :  255 - 0xff -- Background 0xba
    "11010101", -- 3537 - 0xdd1  :  213 - 0xd5
    "10101010", -- 3538 - 0xdd2  :  170 - 0xaa
    "11111111", -- 3539 - 0xdd3  :  255 - 0xff
    "10000000", -- 3540 - 0xdd4  :  128 - 0x80
    "10000000", -- 3541 - 0xdd5  :  128 - 0x80
    "10010101", -- 3542 - 0xdd6  :  149 - 0x95
    "11111111", -- 3543 - 0xdd7  :  255 - 0xff
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0 -- Background 0xbb
    "00000000", -- 3545 - 0xdd9  :    0 - 0x0
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "11111111", -- 3552 - 0xde0  :  255 - 0xff -- Background 0xbc
    "01010101", -- 3553 - 0xde1  :   85 - 0x55
    "10101011", -- 3554 - 0xde2  :  171 - 0xab
    "11111111", -- 3555 - 0xde3  :  255 - 0xff
    "01100001", -- 3556 - 0xde4  :   97 - 0x61
    "00100011", -- 3557 - 0xde5  :   35 - 0x23
    "01100101", -- 3558 - 0xde6  :  101 - 0x65
    "11111111", -- 3559 - 0xde7  :  255 - 0xff
    "00000000", -- 3560 - 0xde8  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 3569 - 0xdf1  :    0 - 0x0
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "00000000", -- 3573 - 0xdf5  :    0 - 0x0
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00000000", -- 3592 - 0xe08  :    0 - 0x0 -- Background 0xc1
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00000000", -- 3594 - 0xe0a  :    0 - 0x0
    "00000000", -- 3595 - 0xe0b  :    0 - 0x0
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00000000", -- 3608 - 0xe18  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00000000", -- 3611 - 0xe1b  :    0 - 0x0
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "00000000", -- 3624 - 0xe28  :    0 - 0x0 -- Background 0xc5
    "00000000", -- 3625 - 0xe29  :    0 - 0x0
    "00000001", -- 3626 - 0xe2a  :    1 - 0x1
    "00000110", -- 3627 - 0xe2b  :    6 - 0x6
    "00001010", -- 3628 - 0xe2c  :   10 - 0xa
    "00010100", -- 3629 - 0xe2d  :   20 - 0x14
    "00010000", -- 3630 - 0xe2e  :   16 - 0x10
    "00101000", -- 3631 - 0xe2f  :   40 - 0x28
    "00011111", -- 3632 - 0xe30  :   31 - 0x1f -- Background 0xc6
    "01100000", -- 3633 - 0xe31  :   96 - 0x60
    "10100000", -- 3634 - 0xe32  :  160 - 0xa0
    "01000000", -- 3635 - 0xe33  :   64 - 0x40
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "00000000", -- 3637 - 0xe35  :    0 - 0x0
    "00000000", -- 3638 - 0xe36  :    0 - 0x0
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "00110000", -- 3640 - 0xe38  :   48 - 0x30 -- Background 0xc7
    "01000000", -- 3641 - 0xe39  :   64 - 0x40
    "01100000", -- 3642 - 0xe3a  :   96 - 0x60
    "11000000", -- 3643 - 0xe3b  :  192 - 0xc0
    "10000000", -- 3644 - 0xe3c  :  128 - 0x80
    "10100000", -- 3645 - 0xe3d  :  160 - 0xa0
    "11000000", -- 3646 - 0xe3e  :  192 - 0xc0
    "10000000", -- 3647 - 0xe3f  :  128 - 0x80
    "11111111", -- 3648 - 0xe40  :  255 - 0xff -- Background 0xc8
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00010100", -- 3656 - 0xe48  :   20 - 0x14 -- Background 0xc9
    "00101010", -- 3657 - 0xe49  :   42 - 0x2a
    "00010110", -- 3658 - 0xe4a  :   22 - 0x16
    "00101011", -- 3659 - 0xe4b  :   43 - 0x2b
    "00010101", -- 3660 - 0xe4c  :   21 - 0x15
    "00101011", -- 3661 - 0xe4d  :   43 - 0x2b
    "00010101", -- 3662 - 0xe4e  :   21 - 0x15
    "00101011", -- 3663 - 0xe4f  :   43 - 0x2b
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Background 0xca
    "00000100", -- 3665 - 0xe51  :    4 - 0x4
    "00000100", -- 3666 - 0xe52  :    4 - 0x4
    "00000101", -- 3667 - 0xe53  :    5 - 0x5
    "00010101", -- 3668 - 0xe54  :   21 - 0x15
    "00010101", -- 3669 - 0xe55  :   21 - 0x15
    "01010101", -- 3670 - 0xe56  :   85 - 0x55
    "01010101", -- 3671 - 0xe57  :   85 - 0x55
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00010000", -- 3674 - 0xe5a  :   16 - 0x10
    "00010000", -- 3675 - 0xe5b  :   16 - 0x10
    "01010001", -- 3676 - 0xe5c  :   81 - 0x51
    "01010101", -- 3677 - 0xe5d  :   85 - 0x55
    "01010101", -- 3678 - 0xe5e  :   85 - 0x55
    "01010101", -- 3679 - 0xe5f  :   85 - 0x55
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000101", -- 3683 - 0xe63  :    5 - 0x5
    "00001111", -- 3684 - 0xe64  :   15 - 0xf
    "00000111", -- 3685 - 0xe65  :    7 - 0x7
    "00000011", -- 3686 - 0xe66  :    3 - 0x3
    "00000001", -- 3687 - 0xe67  :    1 - 0x1
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "10000000", -- 3690 - 0xe6a  :  128 - 0x80
    "11010000", -- 3691 - 0xe6b  :  208 - 0xd0
    "11111000", -- 3692 - 0xe6c  :  248 - 0xf8
    "11110000", -- 3693 - 0xe6d  :  240 - 0xf0
    "11100000", -- 3694 - 0xe6e  :  224 - 0xe0
    "11000000", -- 3695 - 0xe6f  :  192 - 0xc0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "01111000", -- 3699 - 0xe73  :  120 - 0x78
    "11001111", -- 3700 - 0xe74  :  207 - 0xcf
    "10000000", -- 3701 - 0xe75  :  128 - 0x80
    "11001111", -- 3702 - 0xe76  :  207 - 0xcf
    "01001000", -- 3703 - 0xe77  :   72 - 0x48
    "00000000", -- 3704 - 0xe78  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00011110", -- 3707 - 0xe7b  :   30 - 0x1e
    "11110011", -- 3708 - 0xe7c  :  243 - 0xf3
    "00000001", -- 3709 - 0xe7d  :    1 - 0x1
    "11110011", -- 3710 - 0xe7e  :  243 - 0xf3
    "00010010", -- 3711 - 0xe7f  :   18 - 0x12
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00001000", -- 3728 - 0xe90  :    8 - 0x8 -- Background 0xd2
    "00001100", -- 3729 - 0xe91  :   12 - 0xc
    "00001000", -- 3730 - 0xe92  :    8 - 0x8
    "00001000", -- 3731 - 0xe93  :    8 - 0x8
    "00001010", -- 3732 - 0xe94  :   10 - 0xa
    "00001000", -- 3733 - 0xe95  :    8 - 0x8
    "00001000", -- 3734 - 0xe96  :    8 - 0x8
    "00001100", -- 3735 - 0xe97  :   12 - 0xc
    "00010000", -- 3736 - 0xe98  :   16 - 0x10 -- Background 0xd3
    "00010000", -- 3737 - 0xe99  :   16 - 0x10
    "00110000", -- 3738 - 0xe9a  :   48 - 0x30
    "00010000", -- 3739 - 0xe9b  :   16 - 0x10
    "01010000", -- 3740 - 0xe9c  :   80 - 0x50
    "00010000", -- 3741 - 0xe9d  :   16 - 0x10
    "00110000", -- 3742 - 0xe9e  :   48 - 0x30
    "00010000", -- 3743 - 0xe9f  :   16 - 0x10
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "11111000", -- 3752 - 0xea8  :  248 - 0xf8 -- Background 0xd5
    "00000110", -- 3753 - 0xea9  :    6 - 0x6
    "00000001", -- 3754 - 0xeaa  :    1 - 0x1
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "10000000", -- 3762 - 0xeb2  :  128 - 0x80
    "01100000", -- 3763 - 0xeb3  :   96 - 0x60
    "01010000", -- 3764 - 0xeb4  :   80 - 0x50
    "10101000", -- 3765 - 0xeb5  :  168 - 0xa8
    "01011000", -- 3766 - 0xeb6  :   88 - 0x58
    "00101100", -- 3767 - 0xeb7  :   44 - 0x2c
    "10100000", -- 3768 - 0xeb8  :  160 - 0xa0 -- Background 0xd7
    "11000000", -- 3769 - 0xeb9  :  192 - 0xc0
    "10000000", -- 3770 - 0xeba  :  128 - 0x80
    "01010000", -- 3771 - 0xebb  :   80 - 0x50
    "01100000", -- 3772 - 0xebc  :   96 - 0x60
    "00111000", -- 3773 - 0xebd  :   56 - 0x38
    "00001000", -- 3774 - 0xebe  :    8 - 0x8
    "00000111", -- 3775 - 0xebf  :    7 - 0x7
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "11111111", -- 3783 - 0xec7  :  255 - 0xff
    "00010101", -- 3784 - 0xec8  :   21 - 0x15 -- Background 0xd9
    "00101011", -- 3785 - 0xec9  :   43 - 0x2b
    "00010101", -- 3786 - 0xeca  :   21 - 0x15
    "00101010", -- 3787 - 0xecb  :   42 - 0x2a
    "01010110", -- 3788 - 0xecc  :   86 - 0x56
    "10101100", -- 3789 - 0xecd  :  172 - 0xac
    "01010000", -- 3790 - 0xece  :   80 - 0x50
    "11100000", -- 3791 - 0xecf  :  224 - 0xe0
    "00000001", -- 3792 - 0xed0  :    1 - 0x1 -- Background 0xda
    "00001101", -- 3793 - 0xed1  :   13 - 0xd
    "00010011", -- 3794 - 0xed2  :   19 - 0x13
    "00001101", -- 3795 - 0xed3  :   13 - 0xd
    "00000001", -- 3796 - 0xed4  :    1 - 0x1
    "00000001", -- 3797 - 0xed5  :    1 - 0x1
    "00000001", -- 3798 - 0xed6  :    1 - 0x1
    "00000001", -- 3799 - 0xed7  :    1 - 0x1
    "11000000", -- 3800 - 0xed8  :  192 - 0xc0 -- Background 0xdb
    "01000000", -- 3801 - 0xed9  :   64 - 0x40
    "01000000", -- 3802 - 0xeda  :   64 - 0x40
    "01011000", -- 3803 - 0xedb  :   88 - 0x58
    "01100100", -- 3804 - 0xedc  :  100 - 0x64
    "01011000", -- 3805 - 0xedd  :   88 - 0x58
    "01000000", -- 3806 - 0xede  :   64 - 0x40
    "01000000", -- 3807 - 0xedf  :   64 - 0x40
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000110", -- 3811 - 0xee3  :    6 - 0x6
    "00000111", -- 3812 - 0xee4  :    7 - 0x7
    "00000111", -- 3813 - 0xee5  :    7 - 0x7
    "00000111", -- 3814 - 0xee6  :    7 - 0x7
    "00000011", -- 3815 - 0xee7  :    3 - 0x3
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "10110000", -- 3819 - 0xeeb  :  176 - 0xb0
    "11110000", -- 3820 - 0xeec  :  240 - 0xf0
    "11110000", -- 3821 - 0xeed  :  240 - 0xf0
    "11110000", -- 3822 - 0xeee  :  240 - 0xf0
    "11100000", -- 3823 - 0xeef  :  224 - 0xe0
    "11001111", -- 3824 - 0xef0  :  207 - 0xcf -- Background 0xde
    "10000000", -- 3825 - 0xef1  :  128 - 0x80
    "11001111", -- 3826 - 0xef2  :  207 - 0xcf
    "01001000", -- 3827 - 0xef3  :   72 - 0x48
    "01001000", -- 3828 - 0xef4  :   72 - 0x48
    "01001000", -- 3829 - 0xef5  :   72 - 0x48
    "01001000", -- 3830 - 0xef6  :   72 - 0x48
    "01001000", -- 3831 - 0xef7  :   72 - 0x48
    "11110011", -- 3832 - 0xef8  :  243 - 0xf3 -- Background 0xdf
    "00000001", -- 3833 - 0xef9  :    1 - 0x1
    "11110011", -- 3834 - 0xefa  :  243 - 0xf3
    "00010010", -- 3835 - 0xefb  :   18 - 0x12
    "00010010", -- 3836 - 0xefc  :   18 - 0x12
    "00010010", -- 3837 - 0xefd  :   18 - 0x12
    "00010010", -- 3838 - 0xefe  :   18 - 0x12
    "00010010", -- 3839 - 0xeff  :   18 - 0x12
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- Background 0xe1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0 -- Background 0xe3
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000000", -- 3866 - 0xf1a  :    0 - 0x0
    "00000000", -- 3867 - 0xf1b  :    0 - 0x0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "00000000", -- 3880 - 0xf28  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000000", -- 3896 - 0xf38  :    0 - 0x0 -- Background 0xe7
    "00000000", -- 3897 - 0xf39  :    0 - 0x0
    "00000000", -- 3898 - 0xf3a  :    0 - 0x0
    "00000000", -- 3899 - 0xf3b  :    0 - 0x0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "00000000", -- 3915 - 0xf4b  :    0 - 0x0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Background 0xea
    "00000000", -- 3921 - 0xf51  :    0 - 0x0
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 3929 - 0xf59  :    0 - 0x0
    "00000000", -- 3930 - 0xf5a  :    0 - 0x0
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- Background 0xed
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0 -- Background 0xef
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00000000", -- 3976 - 0xf88  :    0 - 0x0 -- Background 0xf1
    "00000000", -- 3977 - 0xf89  :    0 - 0x0
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000000", -- 3979 - 0xf8b  :    0 - 0x0
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Background 0xf4
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- Background 0xf5
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- Background 0xf7
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "00000000", -- 4028 - 0xfbc  :    0 - 0x0
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00000000", -- 4030 - 0xfbe  :    0 - 0x0
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Background 0xf8
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "00000000", -- 4034 - 0xfc2  :    0 - 0x0
    "00000000", -- 4035 - 0xfc3  :    0 - 0x0
    "00000000", -- 4036 - 0xfc4  :    0 - 0x0
    "00000000", -- 4037 - 0xfc5  :    0 - 0x0
    "00000000", -- 4038 - 0xfc6  :    0 - 0x0
    "00000000", -- 4039 - 0xfc7  :    0 - 0x0
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0 -- Background 0xf9
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0 -- Background 0xfb
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "00000000", -- 4059 - 0xfdb  :    0 - 0x0
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "10001110", -- 4066 - 0xfe2  :  142 - 0x8e
    "10001010", -- 4067 - 0xfe3  :  138 - 0x8a
    "10001010", -- 4068 - 0xfe4  :  138 - 0x8a
    "10001010", -- 4069 - 0xfe5  :  138 - 0x8a
    "10001010", -- 4070 - 0xfe6  :  138 - 0x8a
    "11101110", -- 4071 - 0xfe7  :  238 - 0xee
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "01001100", -- 4074 - 0xfea  :   76 - 0x4c
    "10101010", -- 4075 - 0xfeb  :  170 - 0xaa
    "10101010", -- 4076 - 0xfec  :  170 - 0xaa
    "11101010", -- 4077 - 0xfed  :  234 - 0xea
    "10101010", -- 4078 - 0xfee  :  170 - 0xaa
    "10101100", -- 4079 - 0xfef  :  172 - 0xac
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "11101100", -- 4082 - 0xff2  :  236 - 0xec
    "01001010", -- 4083 - 0xff3  :   74 - 0x4a
    "01001010", -- 4084 - 0xff4  :   74 - 0x4a
    "01001010", -- 4085 - 0xff5  :   74 - 0x4a
    "01001010", -- 4086 - 0xff6  :   74 - 0x4a
    "11101010", -- 4087 - 0xff7  :  234 - 0xea
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "01100000", -- 4090 - 0xffa  :   96 - 0x60
    "10001000", -- 4091 - 0xffb  :  136 - 0x88
    "10100000", -- 4092 - 0xffc  :  160 - 0xa0
    "10100000", -- 4093 - 0xffd  :  160 - 0xa0
    "10101000", -- 4094 - 0xffe  :  168 - 0xa8
    "01000000"  -- 4095 - 0xfff  :   64 - 0x40
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
