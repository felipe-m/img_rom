//-   Sprites Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_DONKEYKONG_SPR_PLN1
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 1
      11'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      11'h2: dout <= 8'b00000111; //    2 :   7 - 0x7
      11'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout <= 8'b00000110; //    4 :   6 - 0x6
      11'h5: dout <= 8'b00000110; //    5 :   6 - 0x6
      11'h6: dout <= 8'b00000011; //    6 :   3 - 0x3
      11'h7: dout <= 8'b00000011; //    7 :   3 - 0x3
      11'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      11'h9: dout <= 8'b00010000; //    9 :  16 - 0x10
      11'hA: dout <= 8'b00111100; //   10 :  60 - 0x3c
      11'hB: dout <= 8'b00111111; //   11 :  63 - 0x3f
      11'hC: dout <= 8'b00111111; //   12 :  63 - 0x3f
      11'hD: dout <= 8'b00111100; //   13 :  60 - 0x3c
      11'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      11'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      11'h11: dout <= 8'b11000000; //   17 : 192 - 0xc0
      11'h12: dout <= 8'b11111000; //   18 : 248 - 0xf8
      11'h13: dout <= 8'b01100000; //   19 :  96 - 0x60
      11'h14: dout <= 8'b11011100; //   20 : 220 - 0xdc
      11'h15: dout <= 8'b01101110; //   21 : 110 - 0x6e
      11'h16: dout <= 8'b11000000; //   22 : 192 - 0xc0
      11'h17: dout <= 8'b11111000; //   23 : 248 - 0xf8
      11'h18: dout <= 8'b01010000; //   24 :  80 - 0x50 -- Sprite 0x3
      11'h19: dout <= 8'b00111000; //   25 :  56 - 0x38
      11'h1A: dout <= 8'b00110000; //   26 :  48 - 0x30
      11'h1B: dout <= 8'b11110000; //   27 : 240 - 0xf0
      11'h1C: dout <= 8'b11110000; //   28 : 240 - 0xf0
      11'h1D: dout <= 8'b11100000; //   29 : 224 - 0xe0
      11'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      11'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout <= 8'b00000111; //   32 :   7 - 0x7 -- Sprite 0x4
      11'h21: dout <= 8'b00001111; //   33 :  15 - 0xf
      11'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      11'h23: dout <= 8'b00001101; //   35 :  13 - 0xd
      11'h24: dout <= 8'b00001100; //   36 :  12 - 0xc
      11'h25: dout <= 8'b00000111; //   37 :   7 - 0x7
      11'h26: dout <= 8'b00000111; //   38 :   7 - 0x7
      11'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout <= 8'b00000001; //   40 :   1 - 0x1 -- Sprite 0x5
      11'h29: dout <= 8'b00000011; //   41 :   3 - 0x3
      11'h2A: dout <= 8'b00000001; //   42 :   1 - 0x1
      11'h2B: dout <= 8'b00010111; //   43 :  23 - 0x17
      11'h2C: dout <= 8'b00011111; //   44 :  31 - 0x1f
      11'h2D: dout <= 8'b00011110; //   45 :  30 - 0x1e
      11'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      11'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout <= 8'b10000000; //   48 : 128 - 0x80 -- Sprite 0x6
      11'h31: dout <= 8'b11110000; //   49 : 240 - 0xf0
      11'h32: dout <= 8'b11000000; //   50 : 192 - 0xc0
      11'h33: dout <= 8'b10111000; //   51 : 184 - 0xb8
      11'h34: dout <= 8'b11011100; //   52 : 220 - 0xdc
      11'h35: dout <= 8'b10000000; //   53 : 128 - 0x80
      11'h36: dout <= 8'b11110000; //   54 : 240 - 0xf0
      11'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout <= 8'b10000000; //   56 : 128 - 0x80 -- Sprite 0x7
      11'h39: dout <= 8'b11100000; //   57 : 224 - 0xe0
      11'h3A: dout <= 8'b11110000; //   58 : 240 - 0xf0
      11'h3B: dout <= 8'b11110000; //   59 : 240 - 0xf0
      11'h3C: dout <= 8'b11110000; //   60 : 240 - 0xf0
      11'h3D: dout <= 8'b11100000; //   61 : 224 - 0xe0
      11'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout <= 8'b00000111; //   64 :   7 - 0x7 -- Sprite 0x8
      11'h41: dout <= 8'b00001111; //   65 :  15 - 0xf
      11'h42: dout <= 8'b00000000; //   66 :   0 - 0x0
      11'h43: dout <= 8'b00001101; //   67 :  13 - 0xd
      11'h44: dout <= 8'b00001100; //   68 :  12 - 0xc
      11'h45: dout <= 8'b00000111; //   69 :   7 - 0x7
      11'h46: dout <= 8'b00000111; //   70 :   7 - 0x7
      11'h47: dout <= 8'b00000011; //   71 :   3 - 0x3
      11'h48: dout <= 8'b11000011; //   72 : 195 - 0xc3 -- Sprite 0x9
      11'h49: dout <= 8'b11100011; //   73 : 227 - 0xe3
      11'h4A: dout <= 8'b11001111; //   74 : 207 - 0xcf
      11'h4B: dout <= 8'b00011111; //   75 :  31 - 0x1f
      11'h4C: dout <= 8'b00111111; //   76 :  63 - 0x3f
      11'h4D: dout <= 8'b00001100; //   77 :  12 - 0xc
      11'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      11'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout <= 8'b10000000; //   80 : 128 - 0x80 -- Sprite 0xa
      11'h51: dout <= 8'b11110000; //   81 : 240 - 0xf0
      11'h52: dout <= 8'b11000000; //   82 : 192 - 0xc0
      11'h53: dout <= 8'b10111000; //   83 : 184 - 0xb8
      11'h54: dout <= 8'b11011100; //   84 : 220 - 0xdc
      11'h55: dout <= 8'b10000000; //   85 : 128 - 0x80
      11'h56: dout <= 8'b11110000; //   86 : 240 - 0xf0
      11'h57: dout <= 8'b00000110; //   87 :   6 - 0x6
      11'h58: dout <= 8'b10001110; //   88 : 142 - 0x8e -- Sprite 0xb
      11'h59: dout <= 8'b11100110; //   89 : 230 - 0xe6
      11'h5A: dout <= 8'b11100000; //   90 : 224 - 0xe0
      11'h5B: dout <= 8'b11110000; //   91 : 240 - 0xf0
      11'h5C: dout <= 8'b11110000; //   92 : 240 - 0xf0
      11'h5D: dout <= 8'b01110000; //   93 : 112 - 0x70
      11'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout <= 8'b00000001; //   96 :   1 - 0x1 -- Sprite 0xc
      11'h61: dout <= 8'b00000011; //   97 :   3 - 0x3
      11'h62: dout <= 8'b00000111; //   98 :   7 - 0x7
      11'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      11'h64: dout <= 8'b00000110; //  100 :   6 - 0x6
      11'h65: dout <= 8'b00000110; //  101 :   6 - 0x6
      11'h66: dout <= 8'b00000010; //  102 :   2 - 0x2
      11'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- Sprite 0xd
      11'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      11'h6A: dout <= 8'b00001100; //  106 :  12 - 0xc
      11'h6B: dout <= 8'b00111111; //  107 :  63 - 0x3f
      11'h6C: dout <= 8'b00111111; //  108 :  63 - 0x3f
      11'h6D: dout <= 8'b00111100; //  109 :  60 - 0x3c
      11'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout <= 8'b11000000; //  112 : 192 - 0xc0 -- Sprite 0xe
      11'h71: dout <= 8'b11000000; //  113 : 192 - 0xc0
      11'h72: dout <= 8'b11111000; //  114 : 248 - 0xf8
      11'h73: dout <= 8'b00100000; //  115 :  32 - 0x20
      11'h74: dout <= 8'b00011100; //  116 :  28 - 0x1c
      11'h75: dout <= 8'b00101110; //  117 :  46 - 0x2e
      11'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      11'h77: dout <= 8'b00111000; //  119 :  56 - 0x38
      11'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      11'h79: dout <= 8'b01100000; //  121 :  96 - 0x60
      11'h7A: dout <= 8'b11110000; //  122 : 240 - 0xf0
      11'h7B: dout <= 8'b11110000; //  123 : 240 - 0xf0
      11'h7C: dout <= 8'b11110000; //  124 : 240 - 0xf0
      11'h7D: dout <= 8'b11100000; //  125 : 224 - 0xe0
      11'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      11'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout <= 8'b00000011; //  129 :   3 - 0x3
      11'h82: dout <= 8'b00000111; //  130 :   7 - 0x7
      11'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      11'h84: dout <= 8'b00000110; //  132 :   6 - 0x6
      11'h85: dout <= 8'b00000110; //  133 :   6 - 0x6
      11'h86: dout <= 8'b00000011; //  134 :   3 - 0x3
      11'h87: dout <= 8'b00000011; //  135 :   3 - 0x3
      11'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      11'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      11'h8A: dout <= 8'b00001100; //  138 :  12 - 0xc
      11'h8B: dout <= 8'b00111111; //  139 :  63 - 0x3f
      11'h8C: dout <= 8'b00111111; //  140 :  63 - 0x3f
      11'h8D: dout <= 8'b00111100; //  141 :  60 - 0x3c
      11'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      11'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      11'h91: dout <= 8'b11000000; //  145 : 192 - 0xc0
      11'h92: dout <= 8'b11111000; //  146 : 248 - 0xf8
      11'h93: dout <= 8'b01100000; //  147 :  96 - 0x60
      11'h94: dout <= 8'b11011100; //  148 : 220 - 0xdc
      11'h95: dout <= 8'b01101110; //  149 : 110 - 0x6e
      11'h96: dout <= 8'b11000000; //  150 : 192 - 0xc0
      11'h97: dout <= 8'b11111000; //  151 : 248 - 0xf8
      11'h98: dout <= 8'b01000111; //  152 :  71 - 0x47 -- Sprite 0x13
      11'h99: dout <= 8'b00001111; //  153 :  15 - 0xf
      11'h9A: dout <= 8'b00001110; //  154 :  14 - 0xe
      11'h9B: dout <= 8'b11110000; //  155 : 240 - 0xf0
      11'h9C: dout <= 8'b11110000; //  156 : 240 - 0xf0
      11'h9D: dout <= 8'b11100000; //  157 : 224 - 0xe0
      11'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      11'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout <= 8'b00000111; //  160 :   7 - 0x7 -- Sprite 0x14
      11'hA1: dout <= 8'b00001111; //  161 :  15 - 0xf
      11'hA2: dout <= 8'b00000011; //  162 :   3 - 0x3
      11'hA3: dout <= 8'b00001100; //  163 :  12 - 0xc
      11'hA4: dout <= 8'b00001100; //  164 :  12 - 0xc
      11'hA5: dout <= 8'b00000100; //  165 :   4 - 0x4
      11'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      11'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- Sprite 0x15
      11'hA9: dout <= 8'b00000001; //  169 :   1 - 0x1
      11'hAA: dout <= 8'b00001111; //  170 :  15 - 0xf
      11'hAB: dout <= 8'b00011111; //  171 :  31 - 0x1f
      11'hAC: dout <= 8'b00011111; //  172 :  31 - 0x1f
      11'hAD: dout <= 8'b00011110; //  173 :  30 - 0x1e
      11'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      11'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout <= 8'b10000000; //  176 : 128 - 0x80 -- Sprite 0x16
      11'hB1: dout <= 8'b11110000; //  177 : 240 - 0xf0
      11'hB2: dout <= 8'b11000000; //  178 : 192 - 0xc0
      11'hB3: dout <= 8'b00111000; //  179 :  56 - 0x38
      11'hB4: dout <= 8'b01011100; //  180 :  92 - 0x5c
      11'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      11'hB6: dout <= 8'b01110000; //  182 : 112 - 0x70
      11'hB7: dout <= 8'b01000000; //  183 :  64 - 0x40
      11'hB8: dout <= 8'b11000000; //  184 : 192 - 0xc0 -- Sprite 0x17
      11'hB9: dout <= 8'b11100000; //  185 : 224 - 0xe0
      11'hBA: dout <= 8'b11110000; //  186 : 240 - 0xf0
      11'hBB: dout <= 8'b11110000; //  187 : 240 - 0xf0
      11'hBC: dout <= 8'b11110000; //  188 : 240 - 0xf0
      11'hBD: dout <= 8'b11100000; //  189 : 224 - 0xe0
      11'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      11'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout <= 8'b00000111; //  192 :   7 - 0x7 -- Sprite 0x18
      11'hC1: dout <= 8'b00001111; //  193 :  15 - 0xf
      11'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      11'hC3: dout <= 8'b00001101; //  195 :  13 - 0xd
      11'hC4: dout <= 8'b00001100; //  196 :  12 - 0xc
      11'hC5: dout <= 8'b00000111; //  197 :   7 - 0x7
      11'hC6: dout <= 8'b00000111; //  198 :   7 - 0x7
      11'hC7: dout <= 8'b00000001; //  199 :   1 - 0x1
      11'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x19
      11'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      11'hCA: dout <= 8'b00010011; //  202 :  19 - 0x13
      11'hCB: dout <= 8'b00011111; //  203 :  31 - 0x1f
      11'hCC: dout <= 8'b00011111; //  204 :  31 - 0x1f
      11'hCD: dout <= 8'b00011110; //  205 :  30 - 0x1e
      11'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout <= 8'b10000000; //  208 : 128 - 0x80 -- Sprite 0x1a
      11'hD1: dout <= 8'b11110000; //  209 : 240 - 0xf0
      11'hD2: dout <= 8'b11000000; //  210 : 192 - 0xc0
      11'hD3: dout <= 8'b10111000; //  211 : 184 - 0xb8
      11'hD4: dout <= 8'b11011100; //  212 : 220 - 0xdc
      11'hD5: dout <= 8'b10000000; //  213 : 128 - 0x80
      11'hD6: dout <= 8'b11110000; //  214 : 240 - 0xf0
      11'hD7: dout <= 8'b10000000; //  215 : 128 - 0x80
      11'hD8: dout <= 8'b00000111; //  216 :   7 - 0x7 -- Sprite 0x1b
      11'hD9: dout <= 8'b00000111; //  217 :   7 - 0x7
      11'hDA: dout <= 8'b11111110; //  218 : 254 - 0xfe
      11'hDB: dout <= 8'b11110000; //  219 : 240 - 0xf0
      11'hDC: dout <= 8'b11110000; //  220 : 240 - 0xf0
      11'hDD: dout <= 8'b11100000; //  221 : 224 - 0xe0
      11'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      11'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout <= 8'b00000111; //  224 :   7 - 0x7 -- Sprite 0x1c
      11'hE1: dout <= 8'b00001111; //  225 :  15 - 0xf
      11'hE2: dout <= 8'b00000011; //  226 :   3 - 0x3
      11'hE3: dout <= 8'b00001100; //  227 :  12 - 0xc
      11'hE4: dout <= 8'b00001100; //  228 :  12 - 0xc
      11'hE5: dout <= 8'b00000000; //  229 :   0 - 0x0
      11'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      11'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout <= 8'b00000001; //  232 :   1 - 0x1 -- Sprite 0x1d
      11'hE9: dout <= 8'b00000001; //  233 :   1 - 0x1
      11'hEA: dout <= 8'b00001111; //  234 :  15 - 0xf
      11'hEB: dout <= 8'b00011111; //  235 :  31 - 0x1f
      11'hEC: dout <= 8'b00111111; //  236 :  63 - 0x3f
      11'hED: dout <= 8'b00011100; //  237 :  28 - 0x1c
      11'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout <= 8'b10000000; //  240 : 128 - 0x80 -- Sprite 0x1e
      11'hF1: dout <= 8'b11110000; //  241 : 240 - 0xf0
      11'hF2: dout <= 8'b11000000; //  242 : 192 - 0xc0
      11'hF3: dout <= 8'b00111000; //  243 :  56 - 0x38
      11'hF4: dout <= 8'b01011100; //  244 :  92 - 0x5c
      11'hF5: dout <= 8'b00000000; //  245 :   0 - 0x0
      11'hF6: dout <= 8'b01110000; //  246 : 112 - 0x70
      11'hF7: dout <= 8'b01000000; //  247 :  64 - 0x40
      11'hF8: dout <= 8'b11000000; //  248 : 192 - 0xc0 -- Sprite 0x1f
      11'hF9: dout <= 8'b11100000; //  249 : 224 - 0xe0
      11'hFA: dout <= 8'b11100000; //  250 : 224 - 0xe0
      11'hFB: dout <= 8'b11110000; //  251 : 240 - 0xf0
      11'hFC: dout <= 8'b11110000; //  252 : 240 - 0xf0
      11'hFD: dout <= 8'b01110000; //  253 : 112 - 0x70
      11'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout <= 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x20
      11'h101: dout <= 8'b00001111; //  257 :  15 - 0xf
      11'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout <= 8'b00001101; //  259 :  13 - 0xd
      11'h104: dout <= 8'b00001100; //  260 :  12 - 0xc
      11'h105: dout <= 8'b00000111; //  261 :   7 - 0x7
      11'h106: dout <= 8'b00000111; //  262 :   7 - 0x7
      11'h107: dout <= 8'b00000001; //  263 :   1 - 0x1
      11'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      11'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout <= 8'b00001001; //  266 :   9 - 0x9
      11'h10B: dout <= 8'b00011111; //  267 :  31 - 0x1f
      11'h10C: dout <= 8'b00111111; //  268 :  63 - 0x3f
      11'h10D: dout <= 8'b00011100; //  269 :  28 - 0x1c
      11'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout <= 8'b10000000; //  272 : 128 - 0x80 -- Sprite 0x22
      11'h111: dout <= 8'b11110000; //  273 : 240 - 0xf0
      11'h112: dout <= 8'b11000000; //  274 : 192 - 0xc0
      11'h113: dout <= 8'b10111000; //  275 : 184 - 0xb8
      11'h114: dout <= 8'b11011100; //  276 : 220 - 0xdc
      11'h115: dout <= 8'b10000000; //  277 : 128 - 0x80
      11'h116: dout <= 8'b11110000; //  278 : 240 - 0xf0
      11'h117: dout <= 8'b10000000; //  279 : 128 - 0x80
      11'h118: dout <= 8'b00000111; //  280 :   7 - 0x7 -- Sprite 0x23
      11'h119: dout <= 8'b00000111; //  281 :   7 - 0x7
      11'h11A: dout <= 8'b11101110; //  282 : 238 - 0xee
      11'h11B: dout <= 8'b11110000; //  283 : 240 - 0xf0
      11'h11C: dout <= 8'b11110000; //  284 : 240 - 0xf0
      11'h11D: dout <= 8'b01110000; //  285 : 112 - 0x70
      11'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      11'h121: dout <= 8'b00000111; //  289 :   7 - 0x7
      11'h122: dout <= 8'b00000011; //  290 :   3 - 0x3
      11'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout <= 8'b00000111; //  293 :   7 - 0x7
      11'h126: dout <= 8'b00000100; //  294 :   4 - 0x4
      11'h127: dout <= 8'b00000100; //  295 :   4 - 0x4
      11'h128: dout <= 8'b00011110; //  296 :  30 - 0x1e -- Sprite 0x25
      11'h129: dout <= 8'b00011111; //  297 :  31 - 0x1f
      11'h12A: dout <= 8'b00011111; //  298 :  31 - 0x1f
      11'h12B: dout <= 8'b00011111; //  299 :  31 - 0x1f
      11'h12C: dout <= 8'b00001111; //  300 :  15 - 0xf
      11'h12D: dout <= 8'b00001000; //  301 :   8 - 0x8
      11'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      11'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout <= 8'b00111000; //  304 :  56 - 0x38 -- Sprite 0x26
      11'h131: dout <= 8'b11111000; //  305 : 248 - 0xf8
      11'h132: dout <= 8'b11000000; //  306 : 192 - 0xc0
      11'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout <= 8'b11100000; //  309 : 224 - 0xe0
      11'h136: dout <= 8'b00100000; //  310 :  32 - 0x20
      11'h137: dout <= 8'b00100000; //  311 :  32 - 0x20
      11'h138: dout <= 8'b01111000; //  312 : 120 - 0x78 -- Sprite 0x27
      11'h139: dout <= 8'b11111100; //  313 : 252 - 0xfc
      11'h13A: dout <= 8'b11111100; //  314 : 252 - 0xfc
      11'h13B: dout <= 8'b11111000; //  315 : 248 - 0xf8
      11'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout <= 8'b10000000; //  317 : 128 - 0x80
      11'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      11'h141: dout <= 8'b00000011; //  321 :   3 - 0x3
      11'h142: dout <= 8'b00000111; //  322 :   7 - 0x7
      11'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout <= 8'b00000110; //  324 :   6 - 0x6
      11'h145: dout <= 8'b00000110; //  325 :   6 - 0x6
      11'h146: dout <= 8'b00000011; //  326 :   3 - 0x3
      11'h147: dout <= 8'b01100011; //  327 :  99 - 0x63
      11'h148: dout <= 8'b11100000; //  328 : 224 - 0xe0 -- Sprite 0x29
      11'h149: dout <= 8'b00100001; //  329 :  33 - 0x21
      11'h14A: dout <= 8'b00000001; //  330 :   1 - 0x1
      11'h14B: dout <= 8'b00000111; //  331 :   7 - 0x7
      11'h14C: dout <= 8'b00000111; //  332 :   7 - 0x7
      11'h14D: dout <= 8'b00011111; //  333 :  31 - 0x1f
      11'h14E: dout <= 8'b00001111; //  334 :  15 - 0xf
      11'h14F: dout <= 8'b00000110; //  335 :   6 - 0x6
      11'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x2a
      11'h151: dout <= 8'b11000000; //  337 : 192 - 0xc0
      11'h152: dout <= 8'b11111000; //  338 : 248 - 0xf8
      11'h153: dout <= 8'b01100000; //  339 :  96 - 0x60
      11'h154: dout <= 8'b11011100; //  340 : 220 - 0xdc
      11'h155: dout <= 8'b01101110; //  341 : 110 - 0x6e
      11'h156: dout <= 8'b11000000; //  342 : 192 - 0xc0
      11'h157: dout <= 8'b11111011; //  343 : 251 - 0xfb
      11'h158: dout <= 8'b10000011; //  344 : 131 - 0x83 -- Sprite 0x2b
      11'h159: dout <= 8'b11000000; //  345 : 192 - 0xc0
      11'h15A: dout <= 8'b11110000; //  346 : 240 - 0xf0
      11'h15B: dout <= 8'b11110000; //  347 : 240 - 0xf0
      11'h15C: dout <= 8'b11111100; //  348 : 252 - 0xfc
      11'h15D: dout <= 8'b11111100; //  349 : 252 - 0xfc
      11'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout <= 8'b00000111; //  352 :   7 - 0x7 -- Sprite 0x2c
      11'h161: dout <= 8'b00001111; //  353 :  15 - 0xf
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b00001101; //  355 :  13 - 0xd
      11'h164: dout <= 8'b00001100; //  356 :  12 - 0xc
      11'h165: dout <= 8'b00000111; //  357 :   7 - 0x7
      11'h166: dout <= 8'b00001111; //  358 :  15 - 0xf
      11'h167: dout <= 8'b00000010; //  359 :   2 - 0x2
      11'h168: dout <= 8'b00000001; //  360 :   1 - 0x1 -- Sprite 0x2d
      11'h169: dout <= 8'b11110011; //  361 : 243 - 0xf3
      11'h16A: dout <= 8'b01011111; //  362 :  95 - 0x5f
      11'h16B: dout <= 8'b00011111; //  363 :  31 - 0x1f
      11'h16C: dout <= 8'b00011111; //  364 :  31 - 0x1f
      11'h16D: dout <= 8'b01001111; //  365 :  79 - 0x4f
      11'h16E: dout <= 8'b00110111; //  366 :  55 - 0x37
      11'h16F: dout <= 8'b11000000; //  367 : 192 - 0xc0
      11'h170: dout <= 8'b10000000; //  368 : 128 - 0x80 -- Sprite 0x2e
      11'h171: dout <= 8'b11110000; //  369 : 240 - 0xf0
      11'h172: dout <= 8'b11000000; //  370 : 192 - 0xc0
      11'h173: dout <= 8'b10111000; //  371 : 184 - 0xb8
      11'h174: dout <= 8'b11011100; //  372 : 220 - 0xdc
      11'h175: dout <= 8'b10000000; //  373 : 128 - 0x80
      11'h176: dout <= 8'b11110000; //  374 : 240 - 0xf0
      11'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout <= 8'b10001111; //  376 : 143 - 0x8f -- Sprite 0x2f
      11'h179: dout <= 8'b11100111; //  377 : 231 - 0xe7
      11'h17A: dout <= 8'b11100000; //  378 : 224 - 0xe0
      11'h17B: dout <= 8'b11110000; //  379 : 240 - 0xf0
      11'h17C: dout <= 8'b11001000; //  380 : 200 - 0xc8
      11'h17D: dout <= 8'b10001000; //  381 : 136 - 0x88
      11'h17E: dout <= 8'b00010000; //  382 :  16 - 0x10
      11'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x30
      11'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      11'h182: dout <= 8'b00000000; //  386 :   0 - 0x0
      11'h183: dout <= 8'b00000111; //  387 :   7 - 0x7
      11'h184: dout <= 8'b00001000; //  388 :   8 - 0x8
      11'h185: dout <= 8'b00010000; //  389 :  16 - 0x10
      11'h186: dout <= 8'b00100000; //  390 :  32 - 0x20
      11'h187: dout <= 8'b00100000; //  391 :  32 - 0x20
      11'h188: dout <= 8'b00100000; //  392 :  32 - 0x20 -- Sprite 0x31
      11'h189: dout <= 8'b00100000; //  393 :  32 - 0x20
      11'h18A: dout <= 8'b00010000; //  394 :  16 - 0x10
      11'h18B: dout <= 8'b00001000; //  395 :   8 - 0x8
      11'h18C: dout <= 8'b00000111; //  396 :   7 - 0x7
      11'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      11'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      11'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout <= 8'b11100000; //  403 : 224 - 0xe0
      11'h194: dout <= 8'b00010000; //  404 :  16 - 0x10
      11'h195: dout <= 8'b00001000; //  405 :   8 - 0x8
      11'h196: dout <= 8'b00000100; //  406 :   4 - 0x4
      11'h197: dout <= 8'b00000100; //  407 :   4 - 0x4
      11'h198: dout <= 8'b00000100; //  408 :   4 - 0x4 -- Sprite 0x33
      11'h199: dout <= 8'b00000100; //  409 :   4 - 0x4
      11'h19A: dout <= 8'b00001000; //  410 :   8 - 0x8
      11'h19B: dout <= 8'b00010000; //  411 :  16 - 0x10
      11'h19C: dout <= 8'b11100000; //  412 : 224 - 0xe0
      11'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      11'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      11'h1A2: dout <= 8'b00000000; //  418 :   0 - 0x0
      11'h1A3: dout <= 8'b00000000; //  419 :   0 - 0x0
      11'h1A4: dout <= 8'b00000000; //  420 :   0 - 0x0
      11'h1A5: dout <= 8'b00000011; //  421 :   3 - 0x3
      11'h1A6: dout <= 8'b00000100; //  422 :   4 - 0x4
      11'h1A7: dout <= 8'b00001000; //  423 :   8 - 0x8
      11'h1A8: dout <= 8'b00001000; //  424 :   8 - 0x8 -- Sprite 0x35
      11'h1A9: dout <= 8'b00000100; //  425 :   4 - 0x4
      11'h1AA: dout <= 8'b00000011; //  426 :   3 - 0x3
      11'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      11'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      11'h1B3: dout <= 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout <= 8'b11000000; //  437 : 192 - 0xc0
      11'h1B6: dout <= 8'b00100000; //  438 :  32 - 0x20
      11'h1B7: dout <= 8'b00010000; //  439 :  16 - 0x10
      11'h1B8: dout <= 8'b00010000; //  440 :  16 - 0x10 -- Sprite 0x37
      11'h1B9: dout <= 8'b00100000; //  441 :  32 - 0x20
      11'h1BA: dout <= 8'b11000000; //  442 : 192 - 0xc0
      11'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      11'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      11'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      11'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      11'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout <= 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout <= 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout <= 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout <= 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout <= 8'b00000001; //  456 :   1 - 0x1 -- Sprite 0x39
      11'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout <= 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      11'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout <= 8'b00000001; //  481 :   1 - 0x1
      11'h1E2: dout <= 8'b00000001; //  482 :   1 - 0x1
      11'h1E3: dout <= 8'b01000000; //  483 :  64 - 0x40
      11'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b10000000; //  488 : 128 - 0x80 -- Sprite 0x3d
      11'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b01000000; //  493 :  64 - 0x40
      11'h1EE: dout <= 8'b00000001; //  494 :   1 - 0x1
      11'h1EF: dout <= 8'b00000001; //  495 :   1 - 0x1
      11'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      11'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout <= 8'b00000100; //  499 :   4 - 0x4
      11'h1F4: dout <= 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout <= 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout <= 8'b00000010; //  504 :   2 - 0x2 -- Sprite 0x3f
      11'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout <= 8'b00000100; //  509 :   4 - 0x4
      11'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout <= 8'b00001111; //  512 :  15 - 0xf -- Sprite 0x40
      11'h201: dout <= 8'b00000111; //  513 :   7 - 0x7
      11'h202: dout <= 8'b00000011; //  514 :   3 - 0x3
      11'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout <= 8'b00000001; //  517 :   1 - 0x1
      11'h206: dout <= 8'b00000001; //  518 :   1 - 0x1
      11'h207: dout <= 8'b00000001; //  519 :   1 - 0x1
      11'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      11'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      11'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      11'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      11'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      11'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      11'h20E: dout <= 8'b00000001; //  526 :   1 - 0x1
      11'h20F: dout <= 8'b00000011; //  527 :   3 - 0x3
      11'h210: dout <= 8'b00000111; //  528 :   7 - 0x7 -- Sprite 0x42
      11'h211: dout <= 8'b00000111; //  529 :   7 - 0x7
      11'h212: dout <= 8'b00000111; //  530 :   7 - 0x7
      11'h213: dout <= 8'b00000111; //  531 :   7 - 0x7
      11'h214: dout <= 8'b00000011; //  532 :   3 - 0x3
      11'h215: dout <= 8'b00000001; //  533 :   1 - 0x1
      11'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      11'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      11'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      11'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      11'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      11'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      11'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      11'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout <= 8'b11111111; //  544 : 255 - 0xff -- Sprite 0x44
      11'h221: dout <= 8'b11111111; //  545 : 255 - 0xff
      11'h222: dout <= 8'b11111111; //  546 : 255 - 0xff
      11'h223: dout <= 8'b11111111; //  547 : 255 - 0xff
      11'h224: dout <= 8'b11111111; //  548 : 255 - 0xff
      11'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      11'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      11'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      11'h228: dout <= 8'b11111111; //  552 : 255 - 0xff -- Sprite 0x45
      11'h229: dout <= 8'b01111111; //  553 : 127 - 0x7f
      11'h22A: dout <= 8'b00111111; //  554 :  63 - 0x3f
      11'h22B: dout <= 8'b00011111; //  555 :  31 - 0x1f
      11'h22C: dout <= 8'b00011111; //  556 :  31 - 0x1f
      11'h22D: dout <= 8'b11111111; //  557 : 255 - 0xff
      11'h22E: dout <= 8'b11111111; //  558 : 255 - 0xff
      11'h22F: dout <= 8'b11111111; //  559 : 255 - 0xff
      11'h230: dout <= 8'b11111111; //  560 : 255 - 0xff -- Sprite 0x46
      11'h231: dout <= 8'b11111111; //  561 : 255 - 0xff
      11'h232: dout <= 8'b11111111; //  562 : 255 - 0xff
      11'h233: dout <= 8'b11111111; //  563 : 255 - 0xff
      11'h234: dout <= 8'b11111111; //  564 : 255 - 0xff
      11'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      11'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      11'h237: dout <= 8'b01111111; //  567 : 127 - 0x7f
      11'h238: dout <= 8'b00000111; //  568 :   7 - 0x7 -- Sprite 0x47
      11'h239: dout <= 8'b00000011; //  569 :   3 - 0x3
      11'h23A: dout <= 8'b00000011; //  570 :   3 - 0x3
      11'h23B: dout <= 8'b00000001; //  571 :   1 - 0x1
      11'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      11'h241: dout <= 8'b10000000; //  577 : 128 - 0x80
      11'h242: dout <= 8'b10000000; //  578 : 128 - 0x80
      11'h243: dout <= 8'b11000000; //  579 : 192 - 0xc0
      11'h244: dout <= 8'b11100000; //  580 : 224 - 0xe0
      11'h245: dout <= 8'b11110000; //  581 : 240 - 0xf0
      11'h246: dout <= 8'b11111111; //  582 : 255 - 0xff
      11'h247: dout <= 8'b11111111; //  583 : 255 - 0xff
      11'h248: dout <= 8'b11111111; //  584 : 255 - 0xff -- Sprite 0x49
      11'h249: dout <= 8'b11111111; //  585 : 255 - 0xff
      11'h24A: dout <= 8'b11111111; //  586 : 255 - 0xff
      11'h24B: dout <= 8'b11111111; //  587 : 255 - 0xff
      11'h24C: dout <= 8'b11111111; //  588 : 255 - 0xff
      11'h24D: dout <= 8'b11111111; //  589 : 255 - 0xff
      11'h24E: dout <= 8'b11111111; //  590 : 255 - 0xff
      11'h24F: dout <= 8'b11111111; //  591 : 255 - 0xff
      11'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x4a
      11'h251: dout <= 8'b11111111; //  593 : 255 - 0xff
      11'h252: dout <= 8'b11111111; //  594 : 255 - 0xff
      11'h253: dout <= 8'b11110000; //  595 : 240 - 0xf0
      11'h254: dout <= 8'b10000000; //  596 : 128 - 0x80
      11'h255: dout <= 8'b00000000; //  597 :   0 - 0x0
      11'h256: dout <= 8'b00000000; //  598 :   0 - 0x0
      11'h257: dout <= 8'b10011111; //  599 : 159 - 0x9f
      11'h258: dout <= 8'b11111111; //  600 : 255 - 0xff -- Sprite 0x4b
      11'h259: dout <= 8'b11111111; //  601 : 255 - 0xff
      11'h25A: dout <= 8'b11111001; //  602 : 249 - 0xf9
      11'h25B: dout <= 8'b11111001; //  603 : 249 - 0xf9
      11'h25C: dout <= 8'b01111111; //  604 : 127 - 0x7f
      11'h25D: dout <= 8'b00111111; //  605 :  63 - 0x3f
      11'h25E: dout <= 8'b00011111; //  606 :  31 - 0x1f
      11'h25F: dout <= 8'b00001111; //  607 :  15 - 0xf
      11'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      11'h261: dout <= 8'b00000001; //  609 :   1 - 0x1
      11'h262: dout <= 8'b00000001; //  610 :   1 - 0x1
      11'h263: dout <= 8'b00000011; //  611 :   3 - 0x3
      11'h264: dout <= 8'b00000111; //  612 :   7 - 0x7
      11'h265: dout <= 8'b00001111; //  613 :  15 - 0xf
      11'h266: dout <= 8'b11111111; //  614 : 255 - 0xff
      11'h267: dout <= 8'b11111111; //  615 : 255 - 0xff
      11'h268: dout <= 8'b11111111; //  616 : 255 - 0xff -- Sprite 0x4d
      11'h269: dout <= 8'b11111111; //  617 : 255 - 0xff
      11'h26A: dout <= 8'b11111111; //  618 : 255 - 0xff
      11'h26B: dout <= 8'b11111111; //  619 : 255 - 0xff
      11'h26C: dout <= 8'b11111111; //  620 : 255 - 0xff
      11'h26D: dout <= 8'b11111111; //  621 : 255 - 0xff
      11'h26E: dout <= 8'b11111111; //  622 : 255 - 0xff
      11'h26F: dout <= 8'b11111111; //  623 : 255 - 0xff
      11'h270: dout <= 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x4e
      11'h271: dout <= 8'b11111111; //  625 : 255 - 0xff
      11'h272: dout <= 8'b11111111; //  626 : 255 - 0xff
      11'h273: dout <= 8'b00011111; //  627 :  31 - 0x1f
      11'h274: dout <= 8'b00000011; //  628 :   3 - 0x3
      11'h275: dout <= 8'b00000001; //  629 :   1 - 0x1
      11'h276: dout <= 8'b00000001; //  630 :   1 - 0x1
      11'h277: dout <= 8'b11110011; //  631 : 243 - 0xf3
      11'h278: dout <= 8'b11111111; //  632 : 255 - 0xff -- Sprite 0x4f
      11'h279: dout <= 8'b11111111; //  633 : 255 - 0xff
      11'h27A: dout <= 8'b00111111; //  634 :  63 - 0x3f
      11'h27B: dout <= 8'b00111111; //  635 :  63 - 0x3f
      11'h27C: dout <= 8'b11111100; //  636 : 252 - 0xfc
      11'h27D: dout <= 8'b11111000; //  637 : 248 - 0xf8
      11'h27E: dout <= 8'b11110000; //  638 : 240 - 0xf0
      11'h27F: dout <= 8'b11100000; //  639 : 224 - 0xe0
      11'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x50
      11'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      11'h282: dout <= 8'b11111111; //  642 : 255 - 0xff
      11'h283: dout <= 8'b11111111; //  643 : 255 - 0xff
      11'h284: dout <= 8'b11111111; //  644 : 255 - 0xff
      11'h285: dout <= 8'b11111111; //  645 : 255 - 0xff
      11'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      11'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      11'h288: dout <= 8'b11111111; //  648 : 255 - 0xff -- Sprite 0x51
      11'h289: dout <= 8'b11111110; //  649 : 254 - 0xfe
      11'h28A: dout <= 8'b11111100; //  650 : 252 - 0xfc
      11'h28B: dout <= 8'b11111000; //  651 : 248 - 0xf8
      11'h28C: dout <= 8'b11111000; //  652 : 248 - 0xf8
      11'h28D: dout <= 8'b11111111; //  653 : 255 - 0xff
      11'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      11'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      11'h290: dout <= 8'b11111111; //  656 : 255 - 0xff -- Sprite 0x52
      11'h291: dout <= 8'b11111111; //  657 : 255 - 0xff
      11'h292: dout <= 8'b11111111; //  658 : 255 - 0xff
      11'h293: dout <= 8'b11111111; //  659 : 255 - 0xff
      11'h294: dout <= 8'b11111111; //  660 : 255 - 0xff
      11'h295: dout <= 8'b11111111; //  661 : 255 - 0xff
      11'h296: dout <= 8'b11111110; //  662 : 254 - 0xfe
      11'h297: dout <= 8'b11111100; //  663 : 252 - 0xfc
      11'h298: dout <= 8'b11100000; //  664 : 224 - 0xe0 -- Sprite 0x53
      11'h299: dout <= 8'b10000000; //  665 : 128 - 0x80
      11'h29A: dout <= 8'b10000000; //  666 : 128 - 0x80
      11'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      11'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      11'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      11'h29E: dout <= 8'b00000000; //  670 :   0 - 0x0
      11'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout <= 8'b11110000; //  672 : 240 - 0xf0 -- Sprite 0x54
      11'h2A1: dout <= 8'b11100000; //  673 : 224 - 0xe0
      11'h2A2: dout <= 8'b11000000; //  674 : 192 - 0xc0
      11'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      11'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      11'h2A5: dout <= 8'b10000000; //  677 : 128 - 0x80
      11'h2A6: dout <= 8'b10000000; //  678 : 128 - 0x80
      11'h2A7: dout <= 8'b10000000; //  679 : 128 - 0x80
      11'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      11'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      11'h2AB: dout <= 8'b00000000; //  683 :   0 - 0x0
      11'h2AC: dout <= 8'b00000000; //  684 :   0 - 0x0
      11'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      11'h2AE: dout <= 8'b10000000; //  686 : 128 - 0x80
      11'h2AF: dout <= 8'b11000000; //  687 : 192 - 0xc0
      11'h2B0: dout <= 8'b11100000; //  688 : 224 - 0xe0 -- Sprite 0x56
      11'h2B1: dout <= 8'b11100000; //  689 : 224 - 0xe0
      11'h2B2: dout <= 8'b11100000; //  690 : 224 - 0xe0
      11'h2B3: dout <= 8'b11100000; //  691 : 224 - 0xe0
      11'h2B4: dout <= 8'b11000000; //  692 : 192 - 0xc0
      11'h2B5: dout <= 8'b10000000; //  693 : 128 - 0x80
      11'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      11'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      11'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      11'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      11'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      11'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      11'h2C1: dout <= 8'b11111111; //  705 : 255 - 0xff
      11'h2C2: dout <= 8'b11111111; //  706 : 255 - 0xff
      11'h2C3: dout <= 8'b11111111; //  707 : 255 - 0xff
      11'h2C4: dout <= 8'b11111111; //  708 : 255 - 0xff
      11'h2C5: dout <= 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout <= 8'b11111111; //  710 : 255 - 0xff
      11'h2C7: dout <= 8'b11111111; //  711 : 255 - 0xff
      11'h2C8: dout <= 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      11'h2C9: dout <= 8'b11111111; //  713 : 255 - 0xff
      11'h2CA: dout <= 8'b11111111; //  714 : 255 - 0xff
      11'h2CB: dout <= 8'b11111111; //  715 : 255 - 0xff
      11'h2CC: dout <= 8'b11111111; //  716 : 255 - 0xff
      11'h2CD: dout <= 8'b11111111; //  717 : 255 - 0xff
      11'h2CE: dout <= 8'b11111111; //  718 : 255 - 0xff
      11'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      11'h2D0: dout <= 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      11'h2D1: dout <= 8'b11111111; //  721 : 255 - 0xff
      11'h2D2: dout <= 8'b11111111; //  722 : 255 - 0xff
      11'h2D3: dout <= 8'b11111111; //  723 : 255 - 0xff
      11'h2D4: dout <= 8'b11111111; //  724 : 255 - 0xff
      11'h2D5: dout <= 8'b11111111; //  725 : 255 - 0xff
      11'h2D6: dout <= 8'b11111111; //  726 : 255 - 0xff
      11'h2D7: dout <= 8'b11111111; //  727 : 255 - 0xff
      11'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      11'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      11'h2DA: dout <= 8'b11111111; //  730 : 255 - 0xff
      11'h2DB: dout <= 8'b11111111; //  731 : 255 - 0xff
      11'h2DC: dout <= 8'b11111111; //  732 : 255 - 0xff
      11'h2DD: dout <= 8'b11111111; //  733 : 255 - 0xff
      11'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      11'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      11'h2E0: dout <= 8'b11111111; //  736 : 255 - 0xff -- Sprite 0x5c
      11'h2E1: dout <= 8'b11111111; //  737 : 255 - 0xff
      11'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      11'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      11'h2E7: dout <= 8'b11111111; //  743 : 255 - 0xff
      11'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      11'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      11'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout <= 8'b11111111; //  747 : 255 - 0xff
      11'h2EC: dout <= 8'b11111111; //  748 : 255 - 0xff
      11'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      11'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      11'h2EF: dout <= 8'b11111111; //  751 : 255 - 0xff
      11'h2F0: dout <= 8'b11111111; //  752 : 255 - 0xff -- Sprite 0x5e
      11'h2F1: dout <= 8'b11111111; //  753 : 255 - 0xff
      11'h2F2: dout <= 8'b11111111; //  754 : 255 - 0xff
      11'h2F3: dout <= 8'b11111111; //  755 : 255 - 0xff
      11'h2F4: dout <= 8'b11111111; //  756 : 255 - 0xff
      11'h2F5: dout <= 8'b11111111; //  757 : 255 - 0xff
      11'h2F6: dout <= 8'b11111111; //  758 : 255 - 0xff
      11'h2F7: dout <= 8'b11111111; //  759 : 255 - 0xff
      11'h2F8: dout <= 8'b11111111; //  760 : 255 - 0xff -- Sprite 0x5f
      11'h2F9: dout <= 8'b11111111; //  761 : 255 - 0xff
      11'h2FA: dout <= 8'b11111111; //  762 : 255 - 0xff
      11'h2FB: dout <= 8'b11111111; //  763 : 255 - 0xff
      11'h2FC: dout <= 8'b11111111; //  764 : 255 - 0xff
      11'h2FD: dout <= 8'b11111111; //  765 : 255 - 0xff
      11'h2FE: dout <= 8'b11111111; //  766 : 255 - 0xff
      11'h2FF: dout <= 8'b11111111; //  767 : 255 - 0xff
      11'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout <= 8'b00001111; //  769 :  15 - 0xf
      11'h302: dout <= 8'b00101000; //  770 :  40 - 0x28
      11'h303: dout <= 8'b01011100; //  771 :  92 - 0x5c
      11'h304: dout <= 8'b00111111; //  772 :  63 - 0x3f
      11'h305: dout <= 8'b01111111; //  773 : 127 - 0x7f
      11'h306: dout <= 8'b01111111; //  774 : 127 - 0x7f
      11'h307: dout <= 8'b01111111; //  775 : 127 - 0x7f
      11'h308: dout <= 8'b01111111; //  776 : 127 - 0x7f -- Sprite 0x61
      11'h309: dout <= 8'b00111110; //  777 :  62 - 0x3e
      11'h30A: dout <= 8'b00011111; //  778 :  31 - 0x1f
      11'h30B: dout <= 8'b00011111; //  779 :  31 - 0x1f
      11'h30C: dout <= 8'b00001000; //  780 :   8 - 0x8
      11'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      11'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      11'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      11'h310: dout <= 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      11'h311: dout <= 8'b10000000; //  785 : 128 - 0x80
      11'h312: dout <= 8'b01000000; //  786 :  64 - 0x40
      11'h313: dout <= 8'b11000100; //  787 : 196 - 0xc4
      11'h314: dout <= 8'b11110110; //  788 : 246 - 0xf6
      11'h315: dout <= 8'b11111110; //  789 : 254 - 0xfe
      11'h316: dout <= 8'b11111100; //  790 : 252 - 0xfc
      11'h317: dout <= 8'b11111100; //  791 : 252 - 0xfc
      11'h318: dout <= 8'b11111000; //  792 : 248 - 0xf8 -- Sprite 0x63
      11'h319: dout <= 8'b11110000; //  793 : 240 - 0xf0
      11'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      11'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      11'h31C: dout <= 8'b10000000; //  796 : 128 - 0x80
      11'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      11'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      11'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      11'h321: dout <= 8'b00011100; //  801 :  28 - 0x1c
      11'h322: dout <= 8'b00111111; //  802 :  63 - 0x3f
      11'h323: dout <= 8'b01111111; //  803 : 127 - 0x7f
      11'h324: dout <= 8'b11111111; //  804 : 255 - 0xff
      11'h325: dout <= 8'b11111111; //  805 : 255 - 0xff
      11'h326: dout <= 8'b00111110; //  806 :  62 - 0x3e
      11'h327: dout <= 8'b01110000; //  807 : 112 - 0x70
      11'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      11'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      11'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      11'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      11'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      11'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      11'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      11'h331: dout <= 8'b01100000; //  817 :  96 - 0x60
      11'h332: dout <= 8'b11110000; //  818 : 240 - 0xf0
      11'h333: dout <= 8'b11111000; //  819 : 248 - 0xf8
      11'h334: dout <= 8'b11111100; //  820 : 252 - 0xfc
      11'h335: dout <= 8'b11111100; //  821 : 252 - 0xfc
      11'h336: dout <= 8'b11111100; //  822 : 252 - 0xfc
      11'h337: dout <= 8'b11111111; //  823 : 255 - 0xff
      11'h338: dout <= 8'b01111100; //  824 : 124 - 0x7c -- Sprite 0x67
      11'h339: dout <= 8'b11111100; //  825 : 252 - 0xfc
      11'h33A: dout <= 8'b10001000; //  826 : 136 - 0x88
      11'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      11'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      11'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      11'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      11'h341: dout <= 8'b00000111; //  833 :   7 - 0x7
      11'h342: dout <= 8'b00000011; //  834 :   3 - 0x3
      11'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout <= 8'b00000111; //  837 :   7 - 0x7
      11'h346: dout <= 8'b00000100; //  838 :   4 - 0x4
      11'h347: dout <= 8'b00000100; //  839 :   4 - 0x4
      11'h348: dout <= 8'b00001100; //  840 :  12 - 0xc -- Sprite 0x69
      11'h349: dout <= 8'b10011110; //  841 : 158 - 0x9e
      11'h34A: dout <= 8'b11111111; //  842 : 255 - 0xff
      11'h34B: dout <= 8'b00011111; //  843 :  31 - 0x1f
      11'h34C: dout <= 8'b00011111; //  844 :  31 - 0x1f
      11'h34D: dout <= 8'b00011110; //  845 :  30 - 0x1e
      11'h34E: dout <= 8'b00001111; //  846 :  15 - 0xf
      11'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      11'h351: dout <= 8'b11100000; //  849 : 224 - 0xe0
      11'h352: dout <= 8'b11000000; //  850 : 192 - 0xc0
      11'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout <= 8'b11100000; //  853 : 224 - 0xe0
      11'h356: dout <= 8'b00100000; //  854 :  32 - 0x20
      11'h357: dout <= 8'b00100000; //  855 :  32 - 0x20
      11'h358: dout <= 8'b00110000; //  856 :  48 - 0x30 -- Sprite 0x6b
      11'h359: dout <= 8'b01111001; //  857 : 121 - 0x79
      11'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      11'h35B: dout <= 8'b11111000; //  859 : 248 - 0xf8
      11'h35C: dout <= 8'b11111000; //  860 : 248 - 0xf8
      11'h35D: dout <= 8'b01111000; //  861 : 120 - 0x78
      11'h35E: dout <= 8'b11110000; //  862 : 240 - 0xf0
      11'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout <= 8'b00000011; //  864 :   3 - 0x3 -- Sprite 0x6c
      11'h361: dout <= 8'b00000111; //  865 :   7 - 0x7
      11'h362: dout <= 8'b00000010; //  866 :   2 - 0x2
      11'h363: dout <= 8'b00000111; //  867 :   7 - 0x7
      11'h364: dout <= 8'b00000100; //  868 :   4 - 0x4
      11'h365: dout <= 8'b01000110; //  869 :  70 - 0x46
      11'h366: dout <= 8'b11100011; //  870 : 227 - 0xe3
      11'h367: dout <= 8'b11000010; //  871 : 194 - 0xc2
      11'h368: dout <= 8'b01000010; //  872 :  66 - 0x42 -- Sprite 0x6d
      11'h369: dout <= 8'b00000111; //  873 :   7 - 0x7
      11'h36A: dout <= 8'b00000111; //  874 :   7 - 0x7
      11'h36B: dout <= 8'b00000111; //  875 :   7 - 0x7
      11'h36C: dout <= 8'b00000111; //  876 :   7 - 0x7
      11'h36D: dout <= 8'b00000011; //  877 :   3 - 0x3
      11'h36E: dout <= 8'b00000010; //  878 :   2 - 0x2
      11'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout <= 8'b11100000; //  880 : 224 - 0xe0 -- Sprite 0x6e
      11'h371: dout <= 8'b11110000; //  881 : 240 - 0xf0
      11'h372: dout <= 8'b10100000; //  882 : 160 - 0xa0
      11'h373: dout <= 8'b11110000; //  883 : 240 - 0xf0
      11'h374: dout <= 8'b10010000; //  884 : 144 - 0x90
      11'h375: dout <= 8'b00110010; //  885 :  50 - 0x32
      11'h376: dout <= 8'b11100011; //  886 : 227 - 0xe3
      11'h377: dout <= 8'b00100001; //  887 :  33 - 0x21
      11'h378: dout <= 8'b00100000; //  888 :  32 - 0x20 -- Sprite 0x6f
      11'h379: dout <= 8'b01110000; //  889 : 112 - 0x70
      11'h37A: dout <= 8'b11110000; //  890 : 240 - 0xf0
      11'h37B: dout <= 8'b11111000; //  891 : 248 - 0xf8
      11'h37C: dout <= 8'b11111000; //  892 : 248 - 0xf8
      11'h37D: dout <= 8'b11110000; //  893 : 240 - 0xf0
      11'h37E: dout <= 8'b00110000; //  894 :  48 - 0x30
      11'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      11'h381: dout <= 8'b00000001; //  897 :   1 - 0x1
      11'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      11'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      11'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      11'h385: dout <= 8'b00011110; //  901 :  30 - 0x1e
      11'h386: dout <= 8'b01111111; //  902 : 127 - 0x7f
      11'h387: dout <= 8'b00111110; //  903 :  62 - 0x3e
      11'h388: dout <= 8'b00111100; //  904 :  60 - 0x3c -- Sprite 0x71
      11'h389: dout <= 8'b00111110; //  905 :  62 - 0x3e
      11'h38A: dout <= 8'b01111111; //  906 : 127 - 0x7f
      11'h38B: dout <= 8'b01111110; //  907 : 126 - 0x7e
      11'h38C: dout <= 8'b00011000; //  908 :  24 - 0x18
      11'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      11'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout <= 8'b11000000; //  912 : 192 - 0xc0 -- Sprite 0x72
      11'h391: dout <= 8'b11100000; //  913 : 224 - 0xe0
      11'h392: dout <= 8'b01000000; //  914 :  64 - 0x40
      11'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      11'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      11'h395: dout <= 8'b00111010; //  917 :  58 - 0x3a
      11'h396: dout <= 8'b11101111; //  918 : 239 - 0xef
      11'h397: dout <= 8'b01001011; //  919 :  75 - 0x4b
      11'h398: dout <= 8'b01011111; //  920 :  95 - 0x5f -- Sprite 0x73
      11'h399: dout <= 8'b01001011; //  921 :  75 - 0x4b
      11'h39A: dout <= 8'b11101111; //  922 : 239 - 0xef
      11'h39B: dout <= 8'b00111010; //  923 :  58 - 0x3a
      11'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      11'h39E: dout <= 8'b01100000; //  926 :  96 - 0x60
      11'h39F: dout <= 8'b11000000; //  927 : 192 - 0xc0
      11'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      11'h3A1: dout <= 8'b00001100; //  929 :  12 - 0xc
      11'h3A2: dout <= 8'b00001111; //  930 :  15 - 0xf
      11'h3A3: dout <= 8'b00011111; //  931 :  31 - 0x1f
      11'h3A4: dout <= 8'b00011111; //  932 :  31 - 0x1f
      11'h3A5: dout <= 8'b00001111; //  933 :  15 - 0xf
      11'h3A6: dout <= 8'b00001110; //  934 :  14 - 0xe
      11'h3A7: dout <= 8'b00000100; //  935 :   4 - 0x4
      11'h3A8: dout <= 8'b10000100; //  936 : 132 - 0x84 -- Sprite 0x75
      11'h3A9: dout <= 8'b11000111; //  937 : 199 - 0xc7
      11'h3AA: dout <= 8'b01001100; //  938 :  76 - 0x4c
      11'h3AB: dout <= 8'b00001001; //  939 :   9 - 0x9
      11'h3AC: dout <= 8'b00001111; //  940 :  15 - 0xf
      11'h3AD: dout <= 8'b00000101; //  941 :   5 - 0x5
      11'h3AE: dout <= 8'b00001111; //  942 :  15 - 0xf
      11'h3AF: dout <= 8'b00000111; //  943 :   7 - 0x7
      11'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x76
      11'h3B1: dout <= 8'b01000000; //  945 :  64 - 0x40
      11'h3B2: dout <= 8'b11000000; //  946 : 192 - 0xc0
      11'h3B3: dout <= 8'b11100000; //  947 : 224 - 0xe0
      11'h3B4: dout <= 8'b11100000; //  948 : 224 - 0xe0
      11'h3B5: dout <= 8'b11100000; //  949 : 224 - 0xe0
      11'h3B6: dout <= 8'b11100000; //  950 : 224 - 0xe0
      11'h3B7: dout <= 8'b01000010; //  951 :  66 - 0x42
      11'h3B8: dout <= 8'b01000011; //  952 :  67 - 0x43 -- Sprite 0x77
      11'h3B9: dout <= 8'b11000111; //  953 : 199 - 0xc7
      11'h3BA: dout <= 8'b01100010; //  954 :  98 - 0x62
      11'h3BB: dout <= 8'b00100000; //  955 :  32 - 0x20
      11'h3BC: dout <= 8'b11100000; //  956 : 224 - 0xe0
      11'h3BD: dout <= 8'b01000000; //  957 :  64 - 0x40
      11'h3BE: dout <= 8'b11100000; //  958 : 224 - 0xe0
      11'h3BF: dout <= 8'b11000000; //  959 : 192 - 0xc0
      11'h3C0: dout <= 8'b00000011; //  960 :   3 - 0x3 -- Sprite 0x78
      11'h3C1: dout <= 8'b00000100; //  961 :   4 - 0x4
      11'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout <= 8'b01011100; //  964 :  92 - 0x5c
      11'h3C5: dout <= 8'b11110111; //  965 : 247 - 0xf7
      11'h3C6: dout <= 8'b11010010; //  966 : 210 - 0xd2
      11'h3C7: dout <= 8'b11111010; //  967 : 250 - 0xfa
      11'h3C8: dout <= 8'b11010010; //  968 : 210 - 0xd2 -- Sprite 0x79
      11'h3C9: dout <= 8'b11110111; //  969 : 247 - 0xf7
      11'h3CA: dout <= 8'b01011100; //  970 :  92 - 0x5c
      11'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout <= 8'b00000010; //  973 :   2 - 0x2
      11'h3CE: dout <= 8'b00000111; //  974 :   7 - 0x7
      11'h3CF: dout <= 8'b00000011; //  975 :   3 - 0x3
      11'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      11'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout <= 8'b00011000; //  979 :  24 - 0x18
      11'h3D4: dout <= 8'b01111110; //  980 : 126 - 0x7e
      11'h3D5: dout <= 8'b11111110; //  981 : 254 - 0xfe
      11'h3D6: dout <= 8'b01111100; //  982 : 124 - 0x7c
      11'h3D7: dout <= 8'b00111100; //  983 :  60 - 0x3c
      11'h3D8: dout <= 8'b01111100; //  984 : 124 - 0x7c -- Sprite 0x7b
      11'h3D9: dout <= 8'b11111110; //  985 : 254 - 0xfe
      11'h3DA: dout <= 8'b01111000; //  986 : 120 - 0x78
      11'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout <= 8'b10000000; //  990 : 128 - 0x80
      11'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      11'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout <= 8'b00000001; //  994 :   1 - 0x1
      11'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      11'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      11'h3E5: dout <= 8'b00100000; //  997 :  32 - 0x20
      11'h3E6: dout <= 8'b01111100; //  998 : 124 - 0x7c
      11'h3E7: dout <= 8'b01111000; //  999 : 120 - 0x78
      11'h3E8: dout <= 8'b01111100; // 1000 : 124 - 0x7c -- Sprite 0x7d
      11'h3E9: dout <= 8'b11111110; // 1001 : 254 - 0xfe
      11'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout <= 8'b11111110; // 1003 : 254 - 0xfe
      11'h3EC: dout <= 8'b01111100; // 1004 : 124 - 0x7c
      11'h3ED: dout <= 8'b01100000; // 1005 :  96 - 0x60
      11'h3EE: dout <= 8'b11100000; // 1006 : 224 - 0xe0
      11'h3EF: dout <= 8'b11100001; // 1007 : 225 - 0xe1
      11'h3F0: dout <= 8'b01111100; // 1008 : 124 - 0x7c -- Sprite 0x7e
      11'h3F1: dout <= 8'b10000010; // 1009 : 130 - 0x82
      11'h3F2: dout <= 8'b00000001; // 1010 :   1 - 0x1
      11'h3F3: dout <= 8'b10000010; // 1011 : 130 - 0x82
      11'h3F4: dout <= 8'b01111100; // 1012 : 124 - 0x7c
      11'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout <= 8'b00010000; // 1016 :  16 - 0x10 -- Sprite 0x7f
      11'h3F9: dout <= 8'b00011001; // 1017 :  25 - 0x19
      11'h3FA: dout <= 8'b01011010; // 1018 :  90 - 0x5a
      11'h3FB: dout <= 8'b11011111; // 1019 : 223 - 0xdf
      11'h3FC: dout <= 8'b01001111; // 1020 :  79 - 0x4f
      11'h3FD: dout <= 8'b01110011; // 1021 : 115 - 0x73
      11'h3FE: dout <= 8'b11011011; // 1022 : 219 - 0xdb
      11'h3FF: dout <= 8'b00000010; // 1023 :   2 - 0x2
      11'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      11'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      11'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      11'h403: dout <= 8'b00000011; // 1027 :   3 - 0x3
      11'h404: dout <= 8'b00001100; // 1028 :  12 - 0xc
      11'h405: dout <= 8'b00010000; // 1029 :  16 - 0x10
      11'h406: dout <= 8'b00100010; // 1030 :  34 - 0x22
      11'h407: dout <= 8'b00100000; // 1031 :  32 - 0x20
      11'h408: dout <= 8'b00100001; // 1032 :  33 - 0x21 -- Sprite 0x81
      11'h409: dout <= 8'b00100011; // 1033 :  35 - 0x23
      11'h40A: dout <= 8'b00010000; // 1034 :  16 - 0x10
      11'h40B: dout <= 8'b00001100; // 1035 :  12 - 0xc
      11'h40C: dout <= 8'b00000011; // 1036 :   3 - 0x3
      11'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      11'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      11'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      11'h413: dout <= 8'b11000000; // 1043 : 192 - 0xc0
      11'h414: dout <= 8'b00110000; // 1044 :  48 - 0x30
      11'h415: dout <= 8'b00001000; // 1045 :   8 - 0x8
      11'h416: dout <= 8'b01100100; // 1046 : 100 - 0x64
      11'h417: dout <= 8'b11000100; // 1047 : 196 - 0xc4
      11'h418: dout <= 8'b10000100; // 1048 : 132 - 0x84 -- Sprite 0x83
      11'h419: dout <= 8'b00000100; // 1049 :   4 - 0x4
      11'h41A: dout <= 8'b00001000; // 1050 :   8 - 0x8
      11'h41B: dout <= 8'b00110000; // 1051 :  48 - 0x30
      11'h41C: dout <= 8'b11000000; // 1052 : 192 - 0xc0
      11'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      11'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      11'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      11'h423: dout <= 8'b00000011; // 1059 :   3 - 0x3
      11'h424: dout <= 8'b00001100; // 1060 :  12 - 0xc
      11'h425: dout <= 8'b00010000; // 1061 :  16 - 0x10
      11'h426: dout <= 8'b00100110; // 1062 :  38 - 0x26
      11'h427: dout <= 8'b00100011; // 1063 :  35 - 0x23
      11'h428: dout <= 8'b00100001; // 1064 :  33 - 0x21 -- Sprite 0x85
      11'h429: dout <= 8'b00100000; // 1065 :  32 - 0x20
      11'h42A: dout <= 8'b00010000; // 1066 :  16 - 0x10
      11'h42B: dout <= 8'b00001100; // 1067 :  12 - 0xc
      11'h42C: dout <= 8'b00000011; // 1068 :   3 - 0x3
      11'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      11'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      11'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      11'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      11'h433: dout <= 8'b11000000; // 1075 : 192 - 0xc0
      11'h434: dout <= 8'b00110000; // 1076 :  48 - 0x30
      11'h435: dout <= 8'b00001000; // 1077 :   8 - 0x8
      11'h436: dout <= 8'b01000100; // 1078 :  68 - 0x44
      11'h437: dout <= 8'b00000100; // 1079 :   4 - 0x4
      11'h438: dout <= 8'b10000100; // 1080 : 132 - 0x84 -- Sprite 0x87
      11'h439: dout <= 8'b11000100; // 1081 : 196 - 0xc4
      11'h43A: dout <= 8'b00001000; // 1082 :   8 - 0x8
      11'h43B: dout <= 8'b00110000; // 1083 :  48 - 0x30
      11'h43C: dout <= 8'b11000000; // 1084 : 192 - 0xc0
      11'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      11'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      11'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      11'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      11'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      11'h443: dout <= 8'b00000011; // 1091 :   3 - 0x3
      11'h444: dout <= 8'b00001100; // 1092 :  12 - 0xc
      11'h445: dout <= 8'b00010000; // 1093 :  16 - 0x10
      11'h446: dout <= 8'b00100000; // 1094 :  32 - 0x20
      11'h447: dout <= 8'b00100001; // 1095 :  33 - 0x21
      11'h448: dout <= 8'b00100011; // 1096 :  35 - 0x23 -- Sprite 0x89
      11'h449: dout <= 8'b00100110; // 1097 :  38 - 0x26
      11'h44A: dout <= 8'b00010000; // 1098 :  16 - 0x10
      11'h44B: dout <= 8'b00001100; // 1099 :  12 - 0xc
      11'h44C: dout <= 8'b00000011; // 1100 :   3 - 0x3
      11'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      11'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      11'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      11'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      11'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      11'h453: dout <= 8'b11000000; // 1107 : 192 - 0xc0
      11'h454: dout <= 8'b00110000; // 1108 :  48 - 0x30
      11'h455: dout <= 8'b00001000; // 1109 :   8 - 0x8
      11'h456: dout <= 8'b11000100; // 1110 : 196 - 0xc4
      11'h457: dout <= 8'b10000100; // 1111 : 132 - 0x84
      11'h458: dout <= 8'b00000100; // 1112 :   4 - 0x4 -- Sprite 0x8b
      11'h459: dout <= 8'b01000100; // 1113 :  68 - 0x44
      11'h45A: dout <= 8'b00001000; // 1114 :   8 - 0x8
      11'h45B: dout <= 8'b00110000; // 1115 :  48 - 0x30
      11'h45C: dout <= 8'b11000000; // 1116 : 192 - 0xc0
      11'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      11'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      11'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      11'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout <= 8'b00000011; // 1123 :   3 - 0x3
      11'h464: dout <= 8'b00001100; // 1124 :  12 - 0xc
      11'h465: dout <= 8'b00010000; // 1125 :  16 - 0x10
      11'h466: dout <= 8'b00100011; // 1126 :  35 - 0x23
      11'h467: dout <= 8'b00100001; // 1127 :  33 - 0x21
      11'h468: dout <= 8'b00100000; // 1128 :  32 - 0x20 -- Sprite 0x8d
      11'h469: dout <= 8'b00100010; // 1129 :  34 - 0x22
      11'h46A: dout <= 8'b00010000; // 1130 :  16 - 0x10
      11'h46B: dout <= 8'b00001100; // 1131 :  12 - 0xc
      11'h46C: dout <= 8'b00000011; // 1132 :   3 - 0x3
      11'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      11'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      11'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      11'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      11'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      11'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      11'h473: dout <= 8'b11000000; // 1139 : 192 - 0xc0
      11'h474: dout <= 8'b00110000; // 1140 :  48 - 0x30
      11'h475: dout <= 8'b00001000; // 1141 :   8 - 0x8
      11'h476: dout <= 8'b00000100; // 1142 :   4 - 0x4
      11'h477: dout <= 8'b10000100; // 1143 : 132 - 0x84
      11'h478: dout <= 8'b11000100; // 1144 : 196 - 0xc4 -- Sprite 0x8f
      11'h479: dout <= 8'b01100100; // 1145 : 100 - 0x64
      11'h47A: dout <= 8'b00001000; // 1146 :   8 - 0x8
      11'h47B: dout <= 8'b00110000; // 1147 :  48 - 0x30
      11'h47C: dout <= 8'b11000000; // 1148 : 192 - 0xc0
      11'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout <= 8'b00101111; // 1156 :  47 - 0x2f
      11'h485: dout <= 8'b00111111; // 1157 :  63 - 0x3f
      11'h486: dout <= 8'b01100000; // 1158 :  96 - 0x60
      11'h487: dout <= 8'b00100000; // 1159 :  32 - 0x20
      11'h488: dout <= 8'b00100000; // 1160 :  32 - 0x20 -- Sprite 0x91
      11'h489: dout <= 8'b01100000; // 1161 :  96 - 0x60
      11'h48A: dout <= 8'b00111111; // 1162 :  63 - 0x3f
      11'h48B: dout <= 8'b00101111; // 1163 :  47 - 0x2f
      11'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      11'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      11'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      11'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      11'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      11'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      11'h493: dout <= 8'b00000000; // 1171 :   0 - 0x0
      11'h494: dout <= 8'b11111010; // 1172 : 250 - 0xfa
      11'h495: dout <= 8'b11111110; // 1173 : 254 - 0xfe
      11'h496: dout <= 8'b00000011; // 1174 :   3 - 0x3
      11'h497: dout <= 8'b00000010; // 1175 :   2 - 0x2
      11'h498: dout <= 8'b00000010; // 1176 :   2 - 0x2 -- Sprite 0x93
      11'h499: dout <= 8'b00000011; // 1177 :   3 - 0x3
      11'h49A: dout <= 8'b11111110; // 1178 : 254 - 0xfe
      11'h49B: dout <= 8'b11111010; // 1179 : 250 - 0xfa
      11'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      11'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      11'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      11'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      11'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      11'h4A3: dout <= 8'b00001111; // 1187 :  15 - 0xf
      11'h4A4: dout <= 8'b00110000; // 1188 :  48 - 0x30
      11'h4A5: dout <= 8'b01100000; // 1189 :  96 - 0x60
      11'h4A6: dout <= 8'b00111111; // 1190 :  63 - 0x3f
      11'h4A7: dout <= 8'b01111111; // 1191 : 127 - 0x7f
      11'h4A8: dout <= 8'b01111111; // 1192 : 127 - 0x7f -- Sprite 0x95
      11'h4A9: dout <= 8'b00111111; // 1193 :  63 - 0x3f
      11'h4AA: dout <= 8'b01100000; // 1194 :  96 - 0x60
      11'h4AB: dout <= 8'b00110000; // 1195 :  48 - 0x30
      11'h4AC: dout <= 8'b00001111; // 1196 :  15 - 0xf
      11'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      11'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      11'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      11'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      11'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      11'h4B3: dout <= 8'b11111000; // 1203 : 248 - 0xf8
      11'h4B4: dout <= 8'b00000110; // 1204 :   6 - 0x6
      11'h4B5: dout <= 8'b00000011; // 1205 :   3 - 0x3
      11'h4B6: dout <= 8'b11111110; // 1206 : 254 - 0xfe
      11'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      11'h4B8: dout <= 8'b11111111; // 1208 : 255 - 0xff -- Sprite 0x97
      11'h4B9: dout <= 8'b11111110; // 1209 : 254 - 0xfe
      11'h4BA: dout <= 8'b00000011; // 1210 :   3 - 0x3
      11'h4BB: dout <= 8'b00000110; // 1211 :   6 - 0x6
      11'h4BC: dout <= 8'b11111000; // 1212 : 248 - 0xf8
      11'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      11'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      11'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      11'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      11'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      11'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout <= 8'b01000000; // 1219 :  64 - 0x40
      11'h4C4: dout <= 8'b00100000; // 1220 :  32 - 0x20
      11'h4C5: dout <= 8'b00000000; // 1221 :   0 - 0x0
      11'h4C6: dout <= 8'b00000000; // 1222 :   0 - 0x0
      11'h4C7: dout <= 8'b00000001; // 1223 :   1 - 0x1
      11'h4C8: dout <= 8'b00000011; // 1224 :   3 - 0x3 -- Sprite 0x99
      11'h4C9: dout <= 8'b00000111; // 1225 :   7 - 0x7
      11'h4CA: dout <= 8'b00000110; // 1226 :   6 - 0x6
      11'h4CB: dout <= 8'b00000110; // 1227 :   6 - 0x6
      11'h4CC: dout <= 8'b00000111; // 1228 :   7 - 0x7
      11'h4CD: dout <= 8'b00000011; // 1229 :   3 - 0x3
      11'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      11'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      11'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout <= 8'b01000000; // 1234 :  64 - 0x40
      11'h4D3: dout <= 8'b00000000; // 1235 :   0 - 0x0
      11'h4D4: dout <= 8'b00000000; // 1236 :   0 - 0x0
      11'h4D5: dout <= 8'b00001000; // 1237 :   8 - 0x8
      11'h4D6: dout <= 8'b00000000; // 1238 :   0 - 0x0
      11'h4D7: dout <= 8'b01000000; // 1239 :  64 - 0x40
      11'h4D8: dout <= 8'b11100000; // 1240 : 224 - 0xe0 -- Sprite 0x9b
      11'h4D9: dout <= 8'b11110000; // 1241 : 240 - 0xf0
      11'h4DA: dout <= 8'b11010000; // 1242 : 208 - 0xd0
      11'h4DB: dout <= 8'b11010000; // 1243 : 208 - 0xd0
      11'h4DC: dout <= 8'b11110000; // 1244 : 240 - 0xf0
      11'h4DD: dout <= 8'b11100000; // 1245 : 224 - 0xe0
      11'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      11'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      11'h4E1: dout <= 8'b00000000; // 1249 :   0 - 0x0
      11'h4E2: dout <= 8'b00000010; // 1250 :   2 - 0x2
      11'h4E3: dout <= 8'b00000000; // 1251 :   0 - 0x0
      11'h4E4: dout <= 8'b10000000; // 1252 : 128 - 0x80
      11'h4E5: dout <= 8'b00000000; // 1253 :   0 - 0x0
      11'h4E6: dout <= 8'b00000011; // 1254 :   3 - 0x3
      11'h4E7: dout <= 8'b00000111; // 1255 :   7 - 0x7
      11'h4E8: dout <= 8'b00000111; // 1256 :   7 - 0x7 -- Sprite 0x9d
      11'h4E9: dout <= 8'b00001111; // 1257 :  15 - 0xf
      11'h4EA: dout <= 8'b00001110; // 1258 :  14 - 0xe
      11'h4EB: dout <= 8'b00001110; // 1259 :  14 - 0xe
      11'h4EC: dout <= 8'b00001111; // 1260 :  15 - 0xf
      11'h4ED: dout <= 8'b00000111; // 1261 :   7 - 0x7
      11'h4EE: dout <= 8'b00000011; // 1262 :   3 - 0x3
      11'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout <= 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      11'h4F1: dout <= 8'b00000000; // 1265 :   0 - 0x0
      11'h4F2: dout <= 8'b00000000; // 1266 :   0 - 0x0
      11'h4F3: dout <= 8'b00001000; // 1267 :   8 - 0x8
      11'h4F4: dout <= 8'b00000000; // 1268 :   0 - 0x0
      11'h4F5: dout <= 8'b10000000; // 1269 : 128 - 0x80
      11'h4F6: dout <= 8'b00100100; // 1270 :  36 - 0x24
      11'h4F7: dout <= 8'b11000000; // 1271 : 192 - 0xc0
      11'h4F8: dout <= 8'b11110000; // 1272 : 240 - 0xf0 -- Sprite 0x9f
      11'h4F9: dout <= 8'b11111000; // 1273 : 248 - 0xf8
      11'h4FA: dout <= 8'b11011000; // 1274 : 216 - 0xd8
      11'h4FB: dout <= 8'b11011000; // 1275 : 216 - 0xd8
      11'h4FC: dout <= 8'b11111000; // 1276 : 248 - 0xf8
      11'h4FD: dout <= 8'b11110000; // 1277 : 240 - 0xf0
      11'h4FE: dout <= 8'b11000000; // 1278 : 192 - 0xc0
      11'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0xa0
      11'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      11'h502: dout <= 8'b00111000; // 1282 :  56 - 0x38
      11'h503: dout <= 8'b01101100; // 1283 : 108 - 0x6c
      11'h504: dout <= 8'b11000110; // 1284 : 198 - 0xc6
      11'h505: dout <= 8'b10000011; // 1285 : 131 - 0x83
      11'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      11'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      11'h508: dout <= 8'b11111111; // 1288 : 255 - 0xff -- Sprite 0xa1
      11'h509: dout <= 8'b11111111; // 1289 : 255 - 0xff
      11'h50A: dout <= 8'b00111000; // 1290 :  56 - 0x38
      11'h50B: dout <= 8'b01101100; // 1291 : 108 - 0x6c
      11'h50C: dout <= 8'b11000110; // 1292 : 198 - 0xc6
      11'h50D: dout <= 8'b10000011; // 1293 : 131 - 0x83
      11'h50E: dout <= 8'b11111111; // 1294 : 255 - 0xff
      11'h50F: dout <= 8'b11111111; // 1295 : 255 - 0xff
      11'h510: dout <= 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0xa2
      11'h511: dout <= 8'b00000000; // 1297 :   0 - 0x0
      11'h512: dout <= 8'b00000000; // 1298 :   0 - 0x0
      11'h513: dout <= 8'b00000000; // 1299 :   0 - 0x0
      11'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      11'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      11'h516: dout <= 8'b00000000; // 1302 :   0 - 0x0
      11'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout <= 8'b11111111; // 1304 : 255 - 0xff -- Sprite 0xa3
      11'h519: dout <= 8'b11111111; // 1305 : 255 - 0xff
      11'h51A: dout <= 8'b11111111; // 1306 : 255 - 0xff
      11'h51B: dout <= 8'b11111111; // 1307 : 255 - 0xff
      11'h51C: dout <= 8'b11111111; // 1308 : 255 - 0xff
      11'h51D: dout <= 8'b11111111; // 1309 : 255 - 0xff
      11'h51E: dout <= 8'b11111111; // 1310 : 255 - 0xff
      11'h51F: dout <= 8'b11111111; // 1311 : 255 - 0xff
      11'h520: dout <= 8'b11111111; // 1312 : 255 - 0xff -- Sprite 0xa4
      11'h521: dout <= 8'b11111111; // 1313 : 255 - 0xff
      11'h522: dout <= 8'b11111111; // 1314 : 255 - 0xff
      11'h523: dout <= 8'b11111111; // 1315 : 255 - 0xff
      11'h524: dout <= 8'b11111111; // 1316 : 255 - 0xff
      11'h525: dout <= 8'b11111111; // 1317 : 255 - 0xff
      11'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      11'h527: dout <= 8'b11111111; // 1319 : 255 - 0xff
      11'h528: dout <= 8'b11111111; // 1320 : 255 - 0xff -- Sprite 0xa5
      11'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      11'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      11'h52B: dout <= 8'b11111111; // 1323 : 255 - 0xff
      11'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      11'h52D: dout <= 8'b11111111; // 1325 : 255 - 0xff
      11'h52E: dout <= 8'b11111111; // 1326 : 255 - 0xff
      11'h52F: dout <= 8'b11111111; // 1327 : 255 - 0xff
      11'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0xa6
      11'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      11'h532: dout <= 8'b11111111; // 1330 : 255 - 0xff
      11'h533: dout <= 8'b11111111; // 1331 : 255 - 0xff
      11'h534: dout <= 8'b11111111; // 1332 : 255 - 0xff
      11'h535: dout <= 8'b11111111; // 1333 : 255 - 0xff
      11'h536: dout <= 8'b11111111; // 1334 : 255 - 0xff
      11'h537: dout <= 8'b11111111; // 1335 : 255 - 0xff
      11'h538: dout <= 8'b11111111; // 1336 : 255 - 0xff -- Sprite 0xa7
      11'h539: dout <= 8'b11111111; // 1337 : 255 - 0xff
      11'h53A: dout <= 8'b11111111; // 1338 : 255 - 0xff
      11'h53B: dout <= 8'b11111111; // 1339 : 255 - 0xff
      11'h53C: dout <= 8'b11111111; // 1340 : 255 - 0xff
      11'h53D: dout <= 8'b11111111; // 1341 : 255 - 0xff
      11'h53E: dout <= 8'b11111111; // 1342 : 255 - 0xff
      11'h53F: dout <= 8'b11111111; // 1343 : 255 - 0xff
      11'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      11'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      11'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      11'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      11'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      11'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      11'h546: dout <= 8'b00000001; // 1350 :   1 - 0x1
      11'h547: dout <= 8'b00000011; // 1351 :   3 - 0x3
      11'h548: dout <= 8'b00000111; // 1352 :   7 - 0x7 -- Sprite 0xa9
      11'h549: dout <= 8'b00000111; // 1353 :   7 - 0x7
      11'h54A: dout <= 8'b00000011; // 1354 :   3 - 0x3
      11'h54B: dout <= 8'b00100111; // 1355 :  39 - 0x27
      11'h54C: dout <= 8'b00011111; // 1356 :  31 - 0x1f
      11'h54D: dout <= 8'b00000111; // 1357 :   7 - 0x7
      11'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      11'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      11'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      11'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      11'h554: dout <= 8'b00000000; // 1364 :   0 - 0x0
      11'h555: dout <= 8'b11110000; // 1365 : 240 - 0xf0
      11'h556: dout <= 8'b11111000; // 1366 : 248 - 0xf8
      11'h557: dout <= 8'b10101100; // 1367 : 172 - 0xac
      11'h558: dout <= 8'b10101100; // 1368 : 172 - 0xac -- Sprite 0xab
      11'h559: dout <= 8'b11111000; // 1369 : 248 - 0xf8
      11'h55A: dout <= 8'b11111000; // 1370 : 248 - 0xf8
      11'h55B: dout <= 8'b11111000; // 1371 : 248 - 0xf8
      11'h55C: dout <= 8'b11110000; // 1372 : 240 - 0xf0
      11'h55D: dout <= 8'b11000000; // 1373 : 192 - 0xc0
      11'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      11'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      11'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      11'h566: dout <= 8'b00000001; // 1382 :   1 - 0x1
      11'h567: dout <= 8'b00000011; // 1383 :   3 - 0x3
      11'h568: dout <= 8'b00000111; // 1384 :   7 - 0x7 -- Sprite 0xad
      11'h569: dout <= 8'b00000111; // 1385 :   7 - 0x7
      11'h56A: dout <= 8'b00000111; // 1386 :   7 - 0x7
      11'h56B: dout <= 8'b00100111; // 1387 :  39 - 0x27
      11'h56C: dout <= 8'b00011111; // 1388 :  31 - 0x1f
      11'h56D: dout <= 8'b00000111; // 1389 :   7 - 0x7
      11'h56E: dout <= 8'b00000001; // 1390 :   1 - 0x1
      11'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      11'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      11'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      11'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      11'h575: dout <= 8'b11110000; // 1397 : 240 - 0xf0
      11'h576: dout <= 8'b11111000; // 1398 : 248 - 0xf8
      11'h577: dout <= 8'b10101100; // 1399 : 172 - 0xac
      11'h578: dout <= 8'b10101100; // 1400 : 172 - 0xac -- Sprite 0xaf
      11'h579: dout <= 8'b11111000; // 1401 : 248 - 0xf8
      11'h57A: dout <= 8'b11111000; // 1402 : 248 - 0xf8
      11'h57B: dout <= 8'b11111100; // 1403 : 252 - 0xfc
      11'h57C: dout <= 8'b11111100; // 1404 : 252 - 0xfc
      11'h57D: dout <= 8'b11111000; // 1405 : 248 - 0xf8
      11'h57E: dout <= 8'b11110000; // 1406 : 240 - 0xf0
      11'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      11'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0xb0
      11'h581: dout <= 8'b11111111; // 1409 : 255 - 0xff
      11'h582: dout <= 8'b11111111; // 1410 : 255 - 0xff
      11'h583: dout <= 8'b11111111; // 1411 : 255 - 0xff
      11'h584: dout <= 8'b11111111; // 1412 : 255 - 0xff
      11'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      11'h586: dout <= 8'b11111111; // 1414 : 255 - 0xff
      11'h587: dout <= 8'b11111111; // 1415 : 255 - 0xff
      11'h588: dout <= 8'b11111111; // 1416 : 255 - 0xff -- Sprite 0xb1
      11'h589: dout <= 8'b11111111; // 1417 : 255 - 0xff
      11'h58A: dout <= 8'b11111111; // 1418 : 255 - 0xff
      11'h58B: dout <= 8'b11111111; // 1419 : 255 - 0xff
      11'h58C: dout <= 8'b11111111; // 1420 : 255 - 0xff
      11'h58D: dout <= 8'b11111111; // 1421 : 255 - 0xff
      11'h58E: dout <= 8'b11111111; // 1422 : 255 - 0xff
      11'h58F: dout <= 8'b11111111; // 1423 : 255 - 0xff
      11'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0xb2
      11'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      11'h592: dout <= 8'b11111111; // 1426 : 255 - 0xff
      11'h593: dout <= 8'b11111111; // 1427 : 255 - 0xff
      11'h594: dout <= 8'b11111111; // 1428 : 255 - 0xff
      11'h595: dout <= 8'b11111111; // 1429 : 255 - 0xff
      11'h596: dout <= 8'b11111111; // 1430 : 255 - 0xff
      11'h597: dout <= 8'b11111111; // 1431 : 255 - 0xff
      11'h598: dout <= 8'b11111111; // 1432 : 255 - 0xff -- Sprite 0xb3
      11'h599: dout <= 8'b11111111; // 1433 : 255 - 0xff
      11'h59A: dout <= 8'b11111111; // 1434 : 255 - 0xff
      11'h59B: dout <= 8'b11111111; // 1435 : 255 - 0xff
      11'h59C: dout <= 8'b11111111; // 1436 : 255 - 0xff
      11'h59D: dout <= 8'b11111111; // 1437 : 255 - 0xff
      11'h59E: dout <= 8'b11111111; // 1438 : 255 - 0xff
      11'h59F: dout <= 8'b11111111; // 1439 : 255 - 0xff
      11'h5A0: dout <= 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0xb4
      11'h5A1: dout <= 8'b11111111; // 1441 : 255 - 0xff
      11'h5A2: dout <= 8'b11111111; // 1442 : 255 - 0xff
      11'h5A3: dout <= 8'b11111111; // 1443 : 255 - 0xff
      11'h5A4: dout <= 8'b11111111; // 1444 : 255 - 0xff
      11'h5A5: dout <= 8'b11111111; // 1445 : 255 - 0xff
      11'h5A6: dout <= 8'b11111111; // 1446 : 255 - 0xff
      11'h5A7: dout <= 8'b11111111; // 1447 : 255 - 0xff
      11'h5A8: dout <= 8'b11111111; // 1448 : 255 - 0xff -- Sprite 0xb5
      11'h5A9: dout <= 8'b11111111; // 1449 : 255 - 0xff
      11'h5AA: dout <= 8'b11111111; // 1450 : 255 - 0xff
      11'h5AB: dout <= 8'b11111111; // 1451 : 255 - 0xff
      11'h5AC: dout <= 8'b11111111; // 1452 : 255 - 0xff
      11'h5AD: dout <= 8'b11111111; // 1453 : 255 - 0xff
      11'h5AE: dout <= 8'b11111111; // 1454 : 255 - 0xff
      11'h5AF: dout <= 8'b11111111; // 1455 : 255 - 0xff
      11'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0xb6
      11'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      11'h5B2: dout <= 8'b11111111; // 1458 : 255 - 0xff
      11'h5B3: dout <= 8'b11111111; // 1459 : 255 - 0xff
      11'h5B4: dout <= 8'b11111111; // 1460 : 255 - 0xff
      11'h5B5: dout <= 8'b11111111; // 1461 : 255 - 0xff
      11'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      11'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      11'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- Sprite 0xb7
      11'h5B9: dout <= 8'b11111111; // 1465 : 255 - 0xff
      11'h5BA: dout <= 8'b11111111; // 1466 : 255 - 0xff
      11'h5BB: dout <= 8'b11111111; // 1467 : 255 - 0xff
      11'h5BC: dout <= 8'b11111111; // 1468 : 255 - 0xff
      11'h5BD: dout <= 8'b11111111; // 1469 : 255 - 0xff
      11'h5BE: dout <= 8'b11111111; // 1470 : 255 - 0xff
      11'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      11'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      11'h5C1: dout <= 8'b00000111; // 1473 :   7 - 0x7
      11'h5C2: dout <= 8'b00001000; // 1474 :   8 - 0x8
      11'h5C3: dout <= 8'b00010000; // 1475 :  16 - 0x10
      11'h5C4: dout <= 8'b00010000; // 1476 :  16 - 0x10
      11'h5C5: dout <= 8'b00100000; // 1477 :  32 - 0x20
      11'h5C6: dout <= 8'b00100000; // 1478 :  32 - 0x20
      11'h5C7: dout <= 8'b00100000; // 1479 :  32 - 0x20
      11'h5C8: dout <= 8'b00011111; // 1480 :  31 - 0x1f -- Sprite 0xb9
      11'h5C9: dout <= 8'b00111111; // 1481 :  63 - 0x3f
      11'h5CA: dout <= 8'b00111111; // 1482 :  63 - 0x3f
      11'h5CB: dout <= 8'b00111111; // 1483 :  63 - 0x3f
      11'h5CC: dout <= 8'b00111110; // 1484 :  62 - 0x3e
      11'h5CD: dout <= 8'b00111111; // 1485 :  63 - 0x3f
      11'h5CE: dout <= 8'b00111111; // 1486 :  63 - 0x3f
      11'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      11'h5D1: dout <= 8'b00000111; // 1489 :   7 - 0x7
      11'h5D2: dout <= 8'b00011111; // 1490 :  31 - 0x1f
      11'h5D3: dout <= 8'b00111111; // 1491 :  63 - 0x3f
      11'h5D4: dout <= 8'b01111111; // 1492 : 127 - 0x7f
      11'h5D5: dout <= 8'b11111111; // 1493 : 255 - 0xff
      11'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      11'h5D7: dout <= 8'b11011101; // 1495 : 221 - 0xdd
      11'h5D8: dout <= 8'b10001001; // 1496 : 137 - 0x89 -- Sprite 0xbb
      11'h5D9: dout <= 8'b00000001; // 1497 :   1 - 0x1
      11'h5DA: dout <= 8'b00000001; // 1498 :   1 - 0x1
      11'h5DB: dout <= 8'b00000001; // 1499 :   1 - 0x1
      11'h5DC: dout <= 8'b00000001; // 1500 :   1 - 0x1
      11'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      11'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      11'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      11'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      11'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      11'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      11'h5E4: dout <= 8'b00000000; // 1508 :   0 - 0x0
      11'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      11'h5E6: dout <= 8'b00000011; // 1510 :   3 - 0x3
      11'h5E7: dout <= 8'b00000111; // 1511 :   7 - 0x7
      11'h5E8: dout <= 8'b00001111; // 1512 :  15 - 0xf -- Sprite 0xbd
      11'h5E9: dout <= 8'b00001111; // 1513 :  15 - 0xf
      11'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      11'h5EB: dout <= 8'b00011111; // 1515 :  31 - 0x1f
      11'h5EC: dout <= 8'b01111111; // 1516 : 127 - 0x7f
      11'h5ED: dout <= 8'b00011100; // 1517 :  28 - 0x1c
      11'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout <= 8'b00000001; // 1520 :   1 - 0x1 -- Sprite 0xbe
      11'h5F1: dout <= 8'b00000010; // 1521 :   2 - 0x2
      11'h5F2: dout <= 8'b00011001; // 1522 :  25 - 0x19
      11'h5F3: dout <= 8'b00100100; // 1523 :  36 - 0x24
      11'h5F4: dout <= 8'b00011001; // 1524 :  25 - 0x19
      11'h5F5: dout <= 8'b00100010; // 1525 :  34 - 0x22
      11'h5F6: dout <= 8'b00010001; // 1526 :  17 - 0x11
      11'h5F7: dout <= 8'b00101100; // 1527 :  44 - 0x2c
      11'h5F8: dout <= 8'b00011111; // 1528 :  31 - 0x1f -- Sprite 0xbf
      11'h5F9: dout <= 8'b00000111; // 1529 :   7 - 0x7
      11'h5FA: dout <= 8'b00000011; // 1530 :   3 - 0x3
      11'h5FB: dout <= 8'b00000011; // 1531 :   3 - 0x3
      11'h5FC: dout <= 8'b00000001; // 1532 :   1 - 0x1
      11'h5FD: dout <= 8'b00000001; // 1533 :   1 - 0x1
      11'h5FE: dout <= 8'b00000001; // 1534 :   1 - 0x1
      11'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      11'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      11'h603: dout <= 8'b00000001; // 1539 :   1 - 0x1
      11'h604: dout <= 8'b00000011; // 1540 :   3 - 0x3
      11'h605: dout <= 8'b00000111; // 1541 :   7 - 0x7
      11'h606: dout <= 8'b00001101; // 1542 :  13 - 0xd
      11'h607: dout <= 8'b00011001; // 1543 :  25 - 0x19
      11'h608: dout <= 8'b00101001; // 1544 :  41 - 0x29 -- Sprite 0xc1
      11'h609: dout <= 8'b00011001; // 1545 :  25 - 0x19
      11'h60A: dout <= 8'b00001101; // 1546 :  13 - 0xd
      11'h60B: dout <= 8'b00000111; // 1547 :   7 - 0x7
      11'h60C: dout <= 8'b00000011; // 1548 :   3 - 0x3
      11'h60D: dout <= 8'b00000001; // 1549 :   1 - 0x1
      11'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      11'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout <= 8'b10000000; // 1555 : 128 - 0x80
      11'h614: dout <= 8'b11000000; // 1556 : 192 - 0xc0
      11'h615: dout <= 8'b11100000; // 1557 : 224 - 0xe0
      11'h616: dout <= 8'b10110000; // 1558 : 176 - 0xb0
      11'h617: dout <= 8'b10011000; // 1559 : 152 - 0x98
      11'h618: dout <= 8'b10010100; // 1560 : 148 - 0x94 -- Sprite 0xc3
      11'h619: dout <= 8'b10011000; // 1561 : 152 - 0x98
      11'h61A: dout <= 8'b10110000; // 1562 : 176 - 0xb0
      11'h61B: dout <= 8'b11100000; // 1563 : 224 - 0xe0
      11'h61C: dout <= 8'b11000000; // 1564 : 192 - 0xc0
      11'h61D: dout <= 8'b10000000; // 1565 : 128 - 0x80
      11'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      11'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout <= 8'b00000001; // 1575 :   1 - 0x1
      11'h628: dout <= 8'b00001111; // 1576 :  15 - 0xf -- Sprite 0xc5
      11'h629: dout <= 8'b01111001; // 1577 : 121 - 0x79
      11'h62A: dout <= 8'b10100001; // 1578 : 161 - 0xa1
      11'h62B: dout <= 8'b01111001; // 1579 : 121 - 0x79
      11'h62C: dout <= 8'b00001111; // 1580 :  15 - 0xf
      11'h62D: dout <= 8'b00000001; // 1581 :   1 - 0x1
      11'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      11'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      11'h631: dout <= 8'b00000000; // 1585 :   0 - 0x0
      11'h632: dout <= 8'b00000000; // 1586 :   0 - 0x0
      11'h633: dout <= 8'b00000000; // 1587 :   0 - 0x0
      11'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      11'h635: dout <= 8'b00000000; // 1589 :   0 - 0x0
      11'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      11'h637: dout <= 8'b10000000; // 1591 : 128 - 0x80
      11'h638: dout <= 8'b11110000; // 1592 : 240 - 0xf0 -- Sprite 0xc7
      11'h639: dout <= 8'b10011110; // 1593 : 158 - 0x9e
      11'h63A: dout <= 8'b10000101; // 1594 : 133 - 0x85
      11'h63B: dout <= 8'b10011110; // 1595 : 158 - 0x9e
      11'h63C: dout <= 8'b11110000; // 1596 : 240 - 0xf0
      11'h63D: dout <= 8'b10000000; // 1597 : 128 - 0x80
      11'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      11'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      11'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout <= 8'b00011110; // 1603 :  30 - 0x1e
      11'h644: dout <= 8'b00111111; // 1604 :  63 - 0x3f
      11'h645: dout <= 8'b00111111; // 1605 :  63 - 0x3f
      11'h646: dout <= 8'b00111111; // 1606 :  63 - 0x3f
      11'h647: dout <= 8'b00111111; // 1607 :  63 - 0x3f
      11'h648: dout <= 8'b00011111; // 1608 :  31 - 0x1f -- Sprite 0xc9
      11'h649: dout <= 8'b00001111; // 1609 :  15 - 0xf
      11'h64A: dout <= 8'b00000111; // 1610 :   7 - 0x7
      11'h64B: dout <= 8'b00000011; // 1611 :   3 - 0x3
      11'h64C: dout <= 8'b00000001; // 1612 :   1 - 0x1
      11'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      11'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      11'h653: dout <= 8'b00111100; // 1619 :  60 - 0x3c
      11'h654: dout <= 8'b01111110; // 1620 : 126 - 0x7e
      11'h655: dout <= 8'b11111110; // 1621 : 254 - 0xfe
      11'h656: dout <= 8'b11111110; // 1622 : 254 - 0xfe
      11'h657: dout <= 8'b11111110; // 1623 : 254 - 0xfe
      11'h658: dout <= 8'b11111100; // 1624 : 252 - 0xfc -- Sprite 0xcb
      11'h659: dout <= 8'b11111000; // 1625 : 248 - 0xf8
      11'h65A: dout <= 8'b11110000; // 1626 : 240 - 0xf0
      11'h65B: dout <= 8'b11100000; // 1627 : 224 - 0xe0
      11'h65C: dout <= 8'b11000000; // 1628 : 192 - 0xc0
      11'h65D: dout <= 8'b10000000; // 1629 : 128 - 0x80
      11'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout <= 8'b11111111; // 1632 : 255 - 0xff -- Sprite 0xcc
      11'h661: dout <= 8'b11111111; // 1633 : 255 - 0xff
      11'h662: dout <= 8'b11111111; // 1634 : 255 - 0xff
      11'h663: dout <= 8'b11111111; // 1635 : 255 - 0xff
      11'h664: dout <= 8'b11111111; // 1636 : 255 - 0xff
      11'h665: dout <= 8'b11111111; // 1637 : 255 - 0xff
      11'h666: dout <= 8'b11111111; // 1638 : 255 - 0xff
      11'h667: dout <= 8'b11111111; // 1639 : 255 - 0xff
      11'h668: dout <= 8'b11111111; // 1640 : 255 - 0xff -- Sprite 0xcd
      11'h669: dout <= 8'b11111111; // 1641 : 255 - 0xff
      11'h66A: dout <= 8'b11111111; // 1642 : 255 - 0xff
      11'h66B: dout <= 8'b11111111; // 1643 : 255 - 0xff
      11'h66C: dout <= 8'b11111111; // 1644 : 255 - 0xff
      11'h66D: dout <= 8'b11111111; // 1645 : 255 - 0xff
      11'h66E: dout <= 8'b11111111; // 1646 : 255 - 0xff
      11'h66F: dout <= 8'b11111111; // 1647 : 255 - 0xff
      11'h670: dout <= 8'b11111111; // 1648 : 255 - 0xff -- Sprite 0xce
      11'h671: dout <= 8'b11111111; // 1649 : 255 - 0xff
      11'h672: dout <= 8'b11111111; // 1650 : 255 - 0xff
      11'h673: dout <= 8'b11111111; // 1651 : 255 - 0xff
      11'h674: dout <= 8'b11111111; // 1652 : 255 - 0xff
      11'h675: dout <= 8'b11111111; // 1653 : 255 - 0xff
      11'h676: dout <= 8'b11111111; // 1654 : 255 - 0xff
      11'h677: dout <= 8'b11111111; // 1655 : 255 - 0xff
      11'h678: dout <= 8'b11111111; // 1656 : 255 - 0xff -- Sprite 0xcf
      11'h679: dout <= 8'b11111111; // 1657 : 255 - 0xff
      11'h67A: dout <= 8'b11111111; // 1658 : 255 - 0xff
      11'h67B: dout <= 8'b11111111; // 1659 : 255 - 0xff
      11'h67C: dout <= 8'b11111111; // 1660 : 255 - 0xff
      11'h67D: dout <= 8'b11111111; // 1661 : 255 - 0xff
      11'h67E: dout <= 8'b11111111; // 1662 : 255 - 0xff
      11'h67F: dout <= 8'b11111111; // 1663 : 255 - 0xff
      11'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      11'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      11'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      11'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      11'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      11'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      11'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      11'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      11'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      11'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      11'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      11'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      11'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      11'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      11'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      11'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      11'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- Sprite 0xd3
      11'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      11'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      11'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      11'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      11'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      11'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      11'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      11'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      11'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      11'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      11'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      11'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      11'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      11'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      11'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      11'h6AB: dout <= 8'b00000001; // 1707 :   1 - 0x1
      11'h6AC: dout <= 8'b00000011; // 1708 :   3 - 0x3
      11'h6AD: dout <= 8'b01100011; // 1709 :  99 - 0x63
      11'h6AE: dout <= 8'b00110001; // 1710 :  49 - 0x31
      11'h6AF: dout <= 8'b00011111; // 1711 :  31 - 0x1f
      11'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout <= 8'b11111100; // 1714 : 252 - 0xfc
      11'h6B3: dout <= 8'b11111110; // 1715 : 254 - 0xfe
      11'h6B4: dout <= 8'b11000000; // 1716 : 192 - 0xc0
      11'h6B5: dout <= 8'b01000000; // 1717 :  64 - 0x40
      11'h6B6: dout <= 8'b10000000; // 1718 : 128 - 0x80
      11'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      11'h6B8: dout <= 8'b01111111; // 1720 : 127 - 0x7f -- Sprite 0xd7
      11'h6B9: dout <= 8'b00111111; // 1721 :  63 - 0x3f
      11'h6BA: dout <= 8'b01010011; // 1722 :  83 - 0x53
      11'h6BB: dout <= 8'b00000111; // 1723 :   7 - 0x7
      11'h6BC: dout <= 8'b00001100; // 1724 :  12 - 0xc
      11'h6BD: dout <= 8'b00011011; // 1725 :  27 - 0x1b
      11'h6BE: dout <= 8'b00000111; // 1726 :   7 - 0x7
      11'h6BF: dout <= 8'b00000111; // 1727 :   7 - 0x7
      11'h6C0: dout <= 8'b00001111; // 1728 :  15 - 0xf -- Sprite 0xd8
      11'h6C1: dout <= 8'b00001111; // 1729 :  15 - 0xf
      11'h6C2: dout <= 8'b00000011; // 1730 :   3 - 0x3
      11'h6C3: dout <= 8'b00111000; // 1731 :  56 - 0x38
      11'h6C4: dout <= 8'b00111111; // 1732 :  63 - 0x3f
      11'h6C5: dout <= 8'b00001110; // 1733 :  14 - 0xe
      11'h6C6: dout <= 8'b00011100; // 1734 :  28 - 0x1c
      11'h6C7: dout <= 8'b00001110; // 1735 :  14 - 0xe
      11'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      11'h6C9: dout <= 8'b10010000; // 1737 : 144 - 0x90
      11'h6CA: dout <= 8'b11110000; // 1738 : 240 - 0xf0
      11'h6CB: dout <= 8'b11110000; // 1739 : 240 - 0xf0
      11'h6CC: dout <= 8'b00011000; // 1740 :  24 - 0x18
      11'h6CD: dout <= 8'b11111100; // 1741 : 252 - 0xfc
      11'h6CE: dout <= 8'b11110000; // 1742 : 240 - 0xf0
      11'h6CF: dout <= 8'b11111000; // 1743 : 248 - 0xf8
      11'h6D0: dout <= 8'b11111000; // 1744 : 248 - 0xf8 -- Sprite 0xda
      11'h6D1: dout <= 8'b11110000; // 1745 : 240 - 0xf0
      11'h6D2: dout <= 8'b10000111; // 1746 : 135 - 0x87
      11'h6D3: dout <= 8'b00111101; // 1747 :  61 - 0x3d
      11'h6D4: dout <= 8'b11111110; // 1748 : 254 - 0xfe
      11'h6D5: dout <= 8'b00011100; // 1749 :  28 - 0x1c
      11'h6D6: dout <= 8'b00001000; // 1750 :   8 - 0x8
      11'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout <= 8'b01111111; // 1752 : 127 - 0x7f -- Sprite 0xdb
      11'h6D9: dout <= 8'b00111111; // 1753 :  63 - 0x3f
      11'h6DA: dout <= 8'b01010011; // 1754 :  83 - 0x53
      11'h6DB: dout <= 8'b00000011; // 1755 :   3 - 0x3
      11'h6DC: dout <= 8'b00000001; // 1756 :   1 - 0x1
      11'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      11'h6DE: dout <= 8'b00000111; // 1758 :   7 - 0x7
      11'h6DF: dout <= 8'b00011111; // 1759 :  31 - 0x1f
      11'h6E0: dout <= 8'b11001111; // 1760 : 207 - 0xcf -- Sprite 0xdc
      11'h6E1: dout <= 8'b01100011; // 1761 :  99 - 0x63
      11'h6E2: dout <= 8'b00111000; // 1762 :  56 - 0x38
      11'h6E3: dout <= 8'b00111110; // 1763 :  62 - 0x3e
      11'h6E4: dout <= 8'b01111011; // 1764 : 123 - 0x7b
      11'h6E5: dout <= 8'b00110000; // 1765 :  48 - 0x30
      11'h6E6: dout <= 8'b00011000; // 1766 :  24 - 0x18
      11'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      11'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      11'h6E9: dout <= 8'b10010000; // 1769 : 144 - 0x90
      11'h6EA: dout <= 8'b11110000; // 1770 : 240 - 0xf0
      11'h6EB: dout <= 8'b11100000; // 1771 : 224 - 0xe0
      11'h6EC: dout <= 8'b11111000; // 1772 : 248 - 0xf8
      11'h6ED: dout <= 8'b00111000; // 1773 :  56 - 0x38
      11'h6EE: dout <= 8'b11110000; // 1774 : 240 - 0xf0
      11'h6EF: dout <= 8'b11110000; // 1775 : 240 - 0xf0
      11'h6F0: dout <= 8'b11111000; // 1776 : 248 - 0xf8 -- Sprite 0xde
      11'h6F1: dout <= 8'b11111000; // 1777 : 248 - 0xf8
      11'h6F2: dout <= 8'b11111000; // 1778 : 248 - 0xf8
      11'h6F3: dout <= 8'b00111000; // 1779 :  56 - 0x38
      11'h6F4: dout <= 8'b10000000; // 1780 : 128 - 0x80
      11'h6F5: dout <= 8'b11111000; // 1781 : 248 - 0xf8
      11'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      11'h6F7: dout <= 8'b01011100; // 1783 :  92 - 0x5c
      11'h6F8: dout <= 8'b11111111; // 1784 : 255 - 0xff -- Sprite 0xdf
      11'h6F9: dout <= 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout <= 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout <= 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout <= 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout <= 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout <= 8'b11111111; // 1791 : 255 - 0xff
      11'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0xe0
      11'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      11'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      11'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      11'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      11'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      11'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout <= 8'b11111111; // 1802 : 255 - 0xff
      11'h70B: dout <= 8'b11111111; // 1803 : 255 - 0xff
      11'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      11'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      11'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0xe2
      11'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      11'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      11'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      11'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      11'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      11'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      11'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      11'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      11'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      11'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0xe4
      11'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      11'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      11'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      11'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      11'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      11'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      11'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      11'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      11'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      11'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      11'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      11'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      11'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      11'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      11'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0xe6
      11'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      11'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      11'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      11'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      11'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      11'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      11'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      11'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      11'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      11'h73A: dout <= 8'b11111111; // 1850 : 255 - 0xff
      11'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      11'h73C: dout <= 8'b11111111; // 1852 : 255 - 0xff
      11'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      11'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      11'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      11'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      11'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      11'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      11'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      11'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      11'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout <= 8'b11111111; // 1864 : 255 - 0xff -- Sprite 0xe9
      11'h749: dout <= 8'b11111111; // 1865 : 255 - 0xff
      11'h74A: dout <= 8'b11111111; // 1866 : 255 - 0xff
      11'h74B: dout <= 8'b11111111; // 1867 : 255 - 0xff
      11'h74C: dout <= 8'b11111111; // 1868 : 255 - 0xff
      11'h74D: dout <= 8'b11111111; // 1869 : 255 - 0xff
      11'h74E: dout <= 8'b11111111; // 1870 : 255 - 0xff
      11'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      11'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      11'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      11'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      11'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      11'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      11'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      11'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      11'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      11'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff -- Sprite 0xeb
      11'h759: dout <= 8'b11111111; // 1881 : 255 - 0xff
      11'h75A: dout <= 8'b11111111; // 1882 : 255 - 0xff
      11'h75B: dout <= 8'b11111111; // 1883 : 255 - 0xff
      11'h75C: dout <= 8'b11111111; // 1884 : 255 - 0xff
      11'h75D: dout <= 8'b11111111; // 1885 : 255 - 0xff
      11'h75E: dout <= 8'b11111111; // 1886 : 255 - 0xff
      11'h75F: dout <= 8'b11111111; // 1887 : 255 - 0xff
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout <= 8'b00000001; // 1889 :   1 - 0x1
      11'h762: dout <= 8'b00000011; // 1890 :   3 - 0x3
      11'h763: dout <= 8'b00110011; // 1891 :  51 - 0x33
      11'h764: dout <= 8'b00011001; // 1892 :  25 - 0x19
      11'h765: dout <= 8'b00001111; // 1893 :  15 - 0xf
      11'h766: dout <= 8'b00111111; // 1894 :  63 - 0x3f
      11'h767: dout <= 8'b00011111; // 1895 :  31 - 0x1f
      11'h768: dout <= 8'b00101011; // 1896 :  43 - 0x2b -- Sprite 0xed
      11'h769: dout <= 8'b00000111; // 1897 :   7 - 0x7
      11'h76A: dout <= 8'b00000101; // 1898 :   5 - 0x5
      11'h76B: dout <= 8'b00001101; // 1899 :  13 - 0xd
      11'h76C: dout <= 8'b00001011; // 1900 :  11 - 0xb
      11'h76D: dout <= 8'b00011011; // 1901 :  27 - 0x1b
      11'h76E: dout <= 8'b00011011; // 1902 :  27 - 0x1b
      11'h76F: dout <= 8'b00000011; // 1903 :   3 - 0x3
      11'h770: dout <= 8'b00000001; // 1904 :   1 - 0x1 -- Sprite 0xee
      11'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout <= 8'b00000011; // 1906 :   3 - 0x3
      11'h773: dout <= 8'b00000101; // 1907 :   5 - 0x5
      11'h774: dout <= 8'b00001110; // 1908 :  14 - 0xe
      11'h775: dout <= 8'b00001101; // 1909 :  13 - 0xd
      11'h776: dout <= 8'b00000001; // 1910 :   1 - 0x1
      11'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout <= 8'b11111000; // 1912 : 248 - 0xf8 -- Sprite 0xef
      11'h779: dout <= 8'b11111100; // 1913 : 252 - 0xfc
      11'h77A: dout <= 8'b11000000; // 1914 : 192 - 0xc0
      11'h77B: dout <= 8'b01000000; // 1915 :  64 - 0x40
      11'h77C: dout <= 8'b10000000; // 1916 : 128 - 0x80
      11'h77D: dout <= 8'b10000000; // 1917 : 128 - 0x80
      11'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout <= 8'b10000000; // 1919 : 128 - 0x80
      11'h780: dout <= 8'b11010000; // 1920 : 208 - 0xd0 -- Sprite 0xf0
      11'h781: dout <= 8'b11111000; // 1921 : 248 - 0xf8
      11'h782: dout <= 8'b11111000; // 1922 : 248 - 0xf8
      11'h783: dout <= 8'b11101000; // 1923 : 232 - 0xe8
      11'h784: dout <= 8'b11001100; // 1924 : 204 - 0xcc
      11'h785: dout <= 8'b11100110; // 1925 : 230 - 0xe6
      11'h786: dout <= 8'b11111000; // 1926 : 248 - 0xf8
      11'h787: dout <= 8'b11111110; // 1927 : 254 - 0xfe
      11'h788: dout <= 8'b11111110; // 1928 : 254 - 0xfe -- Sprite 0xf1
      11'h789: dout <= 8'b11111110; // 1929 : 254 - 0xfe
      11'h78A: dout <= 8'b00000110; // 1930 :   6 - 0x6
      11'h78B: dout <= 8'b11111000; // 1931 : 248 - 0xf8
      11'h78C: dout <= 8'b00001110; // 1932 :  14 - 0xe
      11'h78D: dout <= 8'b10000000; // 1933 : 128 - 0x80
      11'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout <= 8'b00000001; // 1936 :   1 - 0x1 -- Sprite 0xf2
      11'h791: dout <= 8'b00001111; // 1937 :  15 - 0xf
      11'h792: dout <= 8'b00000111; // 1938 :   7 - 0x7
      11'h793: dout <= 8'b00011101; // 1939 :  29 - 0x1d
      11'h794: dout <= 8'b00111011; // 1940 :  59 - 0x3b
      11'h795: dout <= 8'b00000001; // 1941 :   1 - 0x1
      11'h796: dout <= 8'b00001111; // 1942 :  15 - 0xf
      11'h797: dout <= 8'b00000010; // 1943 :   2 - 0x2
      11'h798: dout <= 8'b00000010; // 1944 :   2 - 0x2 -- Sprite 0xf3
      11'h799: dout <= 8'b00000011; // 1945 :   3 - 0x3
      11'h79A: dout <= 8'b00000010; // 1946 :   2 - 0x2
      11'h79B: dout <= 8'b01110111; // 1947 : 119 - 0x77
      11'h79C: dout <= 8'b00010111; // 1948 :  23 - 0x17
      11'h79D: dout <= 8'b00000001; // 1949 :   1 - 0x1
      11'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout <= 8'b11100000; // 1952 : 224 - 0xe0 -- Sprite 0xf4
      11'h7A1: dout <= 8'b11110000; // 1953 : 240 - 0xf0
      11'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      11'h7A3: dout <= 8'b10110000; // 1955 : 176 - 0xb0
      11'h7A4: dout <= 8'b00110000; // 1956 :  48 - 0x30
      11'h7A5: dout <= 8'b01100000; // 1957 :  96 - 0x60
      11'h7A6: dout <= 8'b11110000; // 1958 : 240 - 0xf0
      11'h7A7: dout <= 8'b00010000; // 1959 :  16 - 0x10
      11'h7A8: dout <= 8'b00110000; // 1960 :  48 - 0x30 -- Sprite 0xf5
      11'h7A9: dout <= 8'b11110000; // 1961 : 240 - 0xf0
      11'h7AA: dout <= 8'b11010000; // 1962 : 208 - 0xd0
      11'h7AB: dout <= 8'b11111100; // 1963 : 252 - 0xfc
      11'h7AC: dout <= 8'b11111110; // 1964 : 254 - 0xfe
      11'h7AD: dout <= 8'b00001000; // 1965 :   8 - 0x8
      11'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout <= 8'b00010000; // 1969 :  16 - 0x10
      11'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout <= 8'b01110100; // 1971 : 116 - 0x74
      11'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      11'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      11'h7BA: dout <= 8'b00010000; // 1978 :  16 - 0x10
      11'h7BB: dout <= 8'b00010000; // 1979 :  16 - 0x10
      11'h7BC: dout <= 8'b00010000; // 1980 :  16 - 0x10
      11'h7BD: dout <= 8'b00010000; // 1981 :  16 - 0x10
      11'h7BE: dout <= 8'b00010000; // 1982 :  16 - 0x10
      11'h7BF: dout <= 8'b00010000; // 1983 :  16 - 0x10
      11'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      11'h7C1: dout <= 8'b00000100; // 1985 :   4 - 0x4
      11'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout <= 8'b00010100; // 1987 :  20 - 0x14
      11'h7C4: dout <= 8'b00000100; // 1988 :   4 - 0x4
      11'h7C5: dout <= 8'b00000100; // 1989 :   4 - 0x4
      11'h7C6: dout <= 8'b00000100; // 1990 :   4 - 0x4
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      11'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout <= 8'b00011111; // 1995 :  31 - 0x1f
      11'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      11'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout <= 8'b11111000; // 2003 : 248 - 0xf8
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      11'h7D9: dout <= 8'b00100000; // 2009 :  32 - 0x20
      11'h7DA: dout <= 8'b00100000; // 2010 :  32 - 0x20
      11'h7DB: dout <= 8'b00101000; // 2011 :  40 - 0x28
      11'h7DC: dout <= 8'b00100000; // 2012 :  32 - 0x20
      11'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout <= 8'b00100000; // 2014 :  32 - 0x20
      11'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      11'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout <= 8'b00001000; // 2018 :   8 - 0x8
      11'h7E3: dout <= 8'b00100101; // 2019 :  37 - 0x25
      11'h7E4: dout <= 8'b00010010; // 2020 :  18 - 0x12
      11'h7E5: dout <= 8'b01010011; // 2021 :  83 - 0x53
      11'h7E6: dout <= 8'b00110011; // 2022 :  51 - 0x33
      11'h7E7: dout <= 8'b00111001; // 2023 :  57 - 0x39
      11'h7E8: dout <= 8'b00001000; // 2024 :   8 - 0x8 -- Sprite 0xfd
      11'h7E9: dout <= 8'b10000000; // 2025 : 128 - 0x80
      11'h7EA: dout <= 8'b00110000; // 2026 :  48 - 0x30
      11'h7EB: dout <= 8'b10011100; // 2027 : 156 - 0x9c
      11'h7EC: dout <= 8'b11001010; // 2028 : 202 - 0xca
      11'h7ED: dout <= 8'b10111000; // 2029 : 184 - 0xb8
      11'h7EE: dout <= 8'b10011000; // 2030 : 152 - 0x98
      11'h7EF: dout <= 8'b01111000; // 2031 : 120 - 0x78
      11'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      11'h7F1: dout <= 8'b00001000; // 2033 :   8 - 0x8
      11'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout <= 8'b01000000; // 2035 :  64 - 0x40
      11'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout <= 8'b00110001; // 2037 :  49 - 0x31
      11'h7F6: dout <= 8'b00111101; // 2038 :  61 - 0x3d
      11'h7F7: dout <= 8'b00011001; // 2039 :  25 - 0x19
      11'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout <= 8'b10000000; // 2041 : 128 - 0x80
      11'h7FA: dout <= 8'b11000000; // 2042 : 192 - 0xc0
      11'h7FB: dout <= 8'b11000000; // 2043 : 192 - 0xc0
      11'h7FC: dout <= 8'b11000000; // 2044 : 192 - 0xc0
      11'h7FD: dout <= 8'b10001000; // 2045 : 136 - 0x88
      11'h7FE: dout <= 8'b10111000; // 2046 : 184 - 0xb8
      11'h7FF: dout <= 8'b10111000; // 2047 : 184 - 0xb8
    endcase
  end

endmodule
