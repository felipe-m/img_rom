---   Background Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG_BG_PLN0 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG_BG_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG_BG_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 0
    "00111000", --    0 -  0x0  :   56 - 0x38 -- Background 0x0
    "01001100", --    1 -  0x1  :   76 - 0x4c
    "11000110", --    2 -  0x2  :  198 - 0xc6
    "11000110", --    3 -  0x3  :  198 - 0xc6
    "11000110", --    4 -  0x4  :  198 - 0xc6
    "01100100", --    5 -  0x5  :  100 - 0x64
    "00111000", --    6 -  0x6  :   56 - 0x38
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00011000", --    8 -  0x8  :   24 - 0x18 -- Background 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "00011000", --   10 -  0xa  :   24 - 0x18
    "00011000", --   11 -  0xb  :   24 - 0x18
    "00011000", --   12 -  0xc  :   24 - 0x18
    "00011000", --   13 -  0xd  :   24 - 0x18
    "01111110", --   14 -  0xe  :  126 - 0x7e
    "00000000", --   15 -  0xf  :    0 - 0x0
    "01111100", --   16 - 0x10  :  124 - 0x7c -- Background 0x2
    "11000110", --   17 - 0x11  :  198 - 0xc6
    "00001110", --   18 - 0x12  :   14 - 0xe
    "00111100", --   19 - 0x13  :   60 - 0x3c
    "01111000", --   20 - 0x14  :  120 - 0x78
    "11100000", --   21 - 0x15  :  224 - 0xe0
    "11111110", --   22 - 0x16  :  254 - 0xfe
    "00000000", --   23 - 0x17  :    0 - 0x0
    "01111110", --   24 - 0x18  :  126 - 0x7e -- Background 0x3
    "00001100", --   25 - 0x19  :   12 - 0xc
    "00011000", --   26 - 0x1a  :   24 - 0x18
    "00111100", --   27 - 0x1b  :   60 - 0x3c
    "00000110", --   28 - 0x1c  :    6 - 0x6
    "11000110", --   29 - 0x1d  :  198 - 0xc6
    "01111100", --   30 - 0x1e  :  124 - 0x7c
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00011100", --   32 - 0x20  :   28 - 0x1c -- Background 0x4
    "00111100", --   33 - 0x21  :   60 - 0x3c
    "01101100", --   34 - 0x22  :  108 - 0x6c
    "11001100", --   35 - 0x23  :  204 - 0xcc
    "11111110", --   36 - 0x24  :  254 - 0xfe
    "00001100", --   37 - 0x25  :   12 - 0xc
    "00001100", --   38 - 0x26  :   12 - 0xc
    "00000000", --   39 - 0x27  :    0 - 0x0
    "11111100", --   40 - 0x28  :  252 - 0xfc -- Background 0x5
    "11000000", --   41 - 0x29  :  192 - 0xc0
    "11111100", --   42 - 0x2a  :  252 - 0xfc
    "00000110", --   43 - 0x2b  :    6 - 0x6
    "00000110", --   44 - 0x2c  :    6 - 0x6
    "11000110", --   45 - 0x2d  :  198 - 0xc6
    "01111100", --   46 - 0x2e  :  124 - 0x7c
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00111100", --   48 - 0x30  :   60 - 0x3c -- Background 0x6
    "01100000", --   49 - 0x31  :   96 - 0x60
    "11000000", --   50 - 0x32  :  192 - 0xc0
    "11111100", --   51 - 0x33  :  252 - 0xfc
    "11000110", --   52 - 0x34  :  198 - 0xc6
    "11000110", --   53 - 0x35  :  198 - 0xc6
    "01111100", --   54 - 0x36  :  124 - 0x7c
    "00000000", --   55 - 0x37  :    0 - 0x0
    "11111110", --   56 - 0x38  :  254 - 0xfe -- Background 0x7
    "11000110", --   57 - 0x39  :  198 - 0xc6
    "00001100", --   58 - 0x3a  :   12 - 0xc
    "00011000", --   59 - 0x3b  :   24 - 0x18
    "00110000", --   60 - 0x3c  :   48 - 0x30
    "00110000", --   61 - 0x3d  :   48 - 0x30
    "00110000", --   62 - 0x3e  :   48 - 0x30
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "01111000", --   64 - 0x40  :  120 - 0x78 -- Background 0x8
    "11000100", --   65 - 0x41  :  196 - 0xc4
    "11100100", --   66 - 0x42  :  228 - 0xe4
    "01111000", --   67 - 0x43  :  120 - 0x78
    "10000110", --   68 - 0x44  :  134 - 0x86
    "10000110", --   69 - 0x45  :  134 - 0x86
    "01111100", --   70 - 0x46  :  124 - 0x7c
    "00000000", --   71 - 0x47  :    0 - 0x0
    "01111100", --   72 - 0x48  :  124 - 0x7c -- Background 0x9
    "11000110", --   73 - 0x49  :  198 - 0xc6
    "11000110", --   74 - 0x4a  :  198 - 0xc6
    "01111110", --   75 - 0x4b  :  126 - 0x7e
    "00000110", --   76 - 0x4c  :    6 - 0x6
    "00001100", --   77 - 0x4d  :   12 - 0xc
    "01111000", --   78 - 0x4e  :  120 - 0x78
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00111000", --   80 - 0x50  :   56 - 0x38 -- Background 0xa
    "01101100", --   81 - 0x51  :  108 - 0x6c
    "11000110", --   82 - 0x52  :  198 - 0xc6
    "11000110", --   83 - 0x53  :  198 - 0xc6
    "11111110", --   84 - 0x54  :  254 - 0xfe
    "11000110", --   85 - 0x55  :  198 - 0xc6
    "11000110", --   86 - 0x56  :  198 - 0xc6
    "00000000", --   87 - 0x57  :    0 - 0x0
    "11111100", --   88 - 0x58  :  252 - 0xfc -- Background 0xb
    "11000110", --   89 - 0x59  :  198 - 0xc6
    "11000110", --   90 - 0x5a  :  198 - 0xc6
    "11111100", --   91 - 0x5b  :  252 - 0xfc
    "11000110", --   92 - 0x5c  :  198 - 0xc6
    "11000110", --   93 - 0x5d  :  198 - 0xc6
    "11111100", --   94 - 0x5e  :  252 - 0xfc
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00111100", --   96 - 0x60  :   60 - 0x3c -- Background 0xc
    "01100110", --   97 - 0x61  :  102 - 0x66
    "11000000", --   98 - 0x62  :  192 - 0xc0
    "11000000", --   99 - 0x63  :  192 - 0xc0
    "11000000", --  100 - 0x64  :  192 - 0xc0
    "01100110", --  101 - 0x65  :  102 - 0x66
    "00111100", --  102 - 0x66  :   60 - 0x3c
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11111000", --  104 - 0x68  :  248 - 0xf8 -- Background 0xd
    "11001100", --  105 - 0x69  :  204 - 0xcc
    "11000110", --  106 - 0x6a  :  198 - 0xc6
    "11000110", --  107 - 0x6b  :  198 - 0xc6
    "11000110", --  108 - 0x6c  :  198 - 0xc6
    "11001100", --  109 - 0x6d  :  204 - 0xcc
    "11111000", --  110 - 0x6e  :  248 - 0xf8
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11111110", --  112 - 0x70  :  254 - 0xfe -- Background 0xe
    "11000000", --  113 - 0x71  :  192 - 0xc0
    "11000000", --  114 - 0x72  :  192 - 0xc0
    "11111100", --  115 - 0x73  :  252 - 0xfc
    "11000000", --  116 - 0x74  :  192 - 0xc0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "11111110", --  118 - 0x76  :  254 - 0xfe
    "00000000", --  119 - 0x77  :    0 - 0x0
    "11111110", --  120 - 0x78  :  254 - 0xfe -- Background 0xf
    "11000000", --  121 - 0x79  :  192 - 0xc0
    "11000000", --  122 - 0x7a  :  192 - 0xc0
    "11111100", --  123 - 0x7b  :  252 - 0xfc
    "11000000", --  124 - 0x7c  :  192 - 0xc0
    "11000000", --  125 - 0x7d  :  192 - 0xc0
    "11000000", --  126 - 0x7e  :  192 - 0xc0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00111110", --  128 - 0x80  :   62 - 0x3e -- Background 0x10
    "01100000", --  129 - 0x81  :   96 - 0x60
    "11000000", --  130 - 0x82  :  192 - 0xc0
    "11011110", --  131 - 0x83  :  222 - 0xde
    "11000110", --  132 - 0x84  :  198 - 0xc6
    "01100110", --  133 - 0x85  :  102 - 0x66
    "01111110", --  134 - 0x86  :  126 - 0x7e
    "00000000", --  135 - 0x87  :    0 - 0x0
    "11000110", --  136 - 0x88  :  198 - 0xc6 -- Background 0x11
    "11000110", --  137 - 0x89  :  198 - 0xc6
    "11000110", --  138 - 0x8a  :  198 - 0xc6
    "11111110", --  139 - 0x8b  :  254 - 0xfe
    "11000110", --  140 - 0x8c  :  198 - 0xc6
    "11000110", --  141 - 0x8d  :  198 - 0xc6
    "11000110", --  142 - 0x8e  :  198 - 0xc6
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01111110", --  144 - 0x90  :  126 - 0x7e -- Background 0x12
    "00011000", --  145 - 0x91  :   24 - 0x18
    "00011000", --  146 - 0x92  :   24 - 0x18
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00011000", --  148 - 0x94  :   24 - 0x18
    "00011000", --  149 - 0x95  :   24 - 0x18
    "01111110", --  150 - 0x96  :  126 - 0x7e
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00011110", --  152 - 0x98  :   30 - 0x1e -- Background 0x13
    "00000110", --  153 - 0x99  :    6 - 0x6
    "00000110", --  154 - 0x9a  :    6 - 0x6
    "00000110", --  155 - 0x9b  :    6 - 0x6
    "11000110", --  156 - 0x9c  :  198 - 0xc6
    "11000110", --  157 - 0x9d  :  198 - 0xc6
    "01111100", --  158 - 0x9e  :  124 - 0x7c
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "11000110", --  160 - 0xa0  :  198 - 0xc6 -- Background 0x14
    "11001100", --  161 - 0xa1  :  204 - 0xcc
    "11011000", --  162 - 0xa2  :  216 - 0xd8
    "11110000", --  163 - 0xa3  :  240 - 0xf0
    "11111000", --  164 - 0xa4  :  248 - 0xf8
    "11011100", --  165 - 0xa5  :  220 - 0xdc
    "11001110", --  166 - 0xa6  :  206 - 0xce
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "01100000", --  168 - 0xa8  :   96 - 0x60 -- Background 0x15
    "01100000", --  169 - 0xa9  :   96 - 0x60
    "01100000", --  170 - 0xaa  :   96 - 0x60
    "01100000", --  171 - 0xab  :   96 - 0x60
    "01100000", --  172 - 0xac  :   96 - 0x60
    "01100000", --  173 - 0xad  :   96 - 0x60
    "01111110", --  174 - 0xae  :  126 - 0x7e
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11000110", --  176 - 0xb0  :  198 - 0xc6 -- Background 0x16
    "11101110", --  177 - 0xb1  :  238 - 0xee
    "11111110", --  178 - 0xb2  :  254 - 0xfe
    "11111110", --  179 - 0xb3  :  254 - 0xfe
    "11010110", --  180 - 0xb4  :  214 - 0xd6
    "11000110", --  181 - 0xb5  :  198 - 0xc6
    "11000110", --  182 - 0xb6  :  198 - 0xc6
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "11000110", --  184 - 0xb8  :  198 - 0xc6 -- Background 0x17
    "11100110", --  185 - 0xb9  :  230 - 0xe6
    "11110110", --  186 - 0xba  :  246 - 0xf6
    "11111110", --  187 - 0xbb  :  254 - 0xfe
    "11011110", --  188 - 0xbc  :  222 - 0xde
    "11001110", --  189 - 0xbd  :  206 - 0xce
    "11000110", --  190 - 0xbe  :  198 - 0xc6
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "01111100", --  192 - 0xc0  :  124 - 0x7c -- Background 0x18
    "11000110", --  193 - 0xc1  :  198 - 0xc6
    "11000110", --  194 - 0xc2  :  198 - 0xc6
    "11000110", --  195 - 0xc3  :  198 - 0xc6
    "11000110", --  196 - 0xc4  :  198 - 0xc6
    "11000110", --  197 - 0xc5  :  198 - 0xc6
    "01111100", --  198 - 0xc6  :  124 - 0x7c
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "11111100", --  200 - 0xc8  :  252 - 0xfc -- Background 0x19
    "11000110", --  201 - 0xc9  :  198 - 0xc6
    "11000110", --  202 - 0xca  :  198 - 0xc6
    "11000110", --  203 - 0xcb  :  198 - 0xc6
    "11111100", --  204 - 0xcc  :  252 - 0xfc
    "11000000", --  205 - 0xcd  :  192 - 0xc0
    "11000000", --  206 - 0xce  :  192 - 0xc0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "01111100", --  208 - 0xd0  :  124 - 0x7c -- Background 0x1a
    "11000110", --  209 - 0xd1  :  198 - 0xc6
    "11000110", --  210 - 0xd2  :  198 - 0xc6
    "11000110", --  211 - 0xd3  :  198 - 0xc6
    "11011110", --  212 - 0xd4  :  222 - 0xde
    "11001100", --  213 - 0xd5  :  204 - 0xcc
    "01111010", --  214 - 0xd6  :  122 - 0x7a
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "11111100", --  216 - 0xd8  :  252 - 0xfc -- Background 0x1b
    "11000110", --  217 - 0xd9  :  198 - 0xc6
    "11000110", --  218 - 0xda  :  198 - 0xc6
    "11001110", --  219 - 0xdb  :  206 - 0xce
    "11111000", --  220 - 0xdc  :  248 - 0xf8
    "11011100", --  221 - 0xdd  :  220 - 0xdc
    "11001110", --  222 - 0xde  :  206 - 0xce
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "01111000", --  224 - 0xe0  :  120 - 0x78 -- Background 0x1c
    "11001100", --  225 - 0xe1  :  204 - 0xcc
    "11000000", --  226 - 0xe2  :  192 - 0xc0
    "01111100", --  227 - 0xe3  :  124 - 0x7c
    "00000110", --  228 - 0xe4  :    6 - 0x6
    "11000110", --  229 - 0xe5  :  198 - 0xc6
    "01111100", --  230 - 0xe6  :  124 - 0x7c
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "01111110", --  232 - 0xe8  :  126 - 0x7e -- Background 0x1d
    "00011000", --  233 - 0xe9  :   24 - 0x18
    "00011000", --  234 - 0xea  :   24 - 0x18
    "00011000", --  235 - 0xeb  :   24 - 0x18
    "00011000", --  236 - 0xec  :   24 - 0x18
    "00011000", --  237 - 0xed  :   24 - 0x18
    "00011000", --  238 - 0xee  :   24 - 0x18
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11000110", --  240 - 0xf0  :  198 - 0xc6 -- Background 0x1e
    "11000110", --  241 - 0xf1  :  198 - 0xc6
    "11000110", --  242 - 0xf2  :  198 - 0xc6
    "11000110", --  243 - 0xf3  :  198 - 0xc6
    "11000110", --  244 - 0xf4  :  198 - 0xc6
    "11000110", --  245 - 0xf5  :  198 - 0xc6
    "01111100", --  246 - 0xf6  :  124 - 0x7c
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "11000110", --  248 - 0xf8  :  198 - 0xc6 -- Background 0x1f
    "11000110", --  249 - 0xf9  :  198 - 0xc6
    "11000110", --  250 - 0xfa  :  198 - 0xc6
    "11101110", --  251 - 0xfb  :  238 - 0xee
    "01111100", --  252 - 0xfc  :  124 - 0x7c
    "00111000", --  253 - 0xfd  :   56 - 0x38
    "00010000", --  254 - 0xfe  :   16 - 0x10
    "00000000", --  255 - 0xff  :    0 - 0x0
    "11000110", --  256 - 0x100  :  198 - 0xc6 -- Background 0x20
    "11000110", --  257 - 0x101  :  198 - 0xc6
    "11010110", --  258 - 0x102  :  214 - 0xd6
    "11111110", --  259 - 0x103  :  254 - 0xfe
    "11111110", --  260 - 0x104  :  254 - 0xfe
    "11101110", --  261 - 0x105  :  238 - 0xee
    "11000110", --  262 - 0x106  :  198 - 0xc6
    "00000000", --  263 - 0x107  :    0 - 0x0
    "11000110", --  264 - 0x108  :  198 - 0xc6 -- Background 0x21
    "11101110", --  265 - 0x109  :  238 - 0xee
    "01111100", --  266 - 0x10a  :  124 - 0x7c
    "00111000", --  267 - 0x10b  :   56 - 0x38
    "01111100", --  268 - 0x10c  :  124 - 0x7c
    "11101110", --  269 - 0x10d  :  238 - 0xee
    "11000110", --  270 - 0x10e  :  198 - 0xc6
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "01100110", --  272 - 0x110  :  102 - 0x66 -- Background 0x22
    "01100110", --  273 - 0x111  :  102 - 0x66
    "01100110", --  274 - 0x112  :  102 - 0x66
    "00111100", --  275 - 0x113  :   60 - 0x3c
    "00011000", --  276 - 0x114  :   24 - 0x18
    "00011000", --  277 - 0x115  :   24 - 0x18
    "00011000", --  278 - 0x116  :   24 - 0x18
    "00000000", --  279 - 0x117  :    0 - 0x0
    "11111110", --  280 - 0x118  :  254 - 0xfe -- Background 0x23
    "00001110", --  281 - 0x119  :   14 - 0xe
    "00011100", --  282 - 0x11a  :   28 - 0x1c
    "00111000", --  283 - 0x11b  :   56 - 0x38
    "01110000", --  284 - 0x11c  :  112 - 0x70
    "11100000", --  285 - 0x11d  :  224 - 0xe0
    "11111110", --  286 - 0x11e  :  254 - 0xfe
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- Background 0x25
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000110", --  298 - 0x12a  :    6 - 0x6
    "00001110", --  299 - 0x12b  :   14 - 0xe
    "00001000", --  300 - 0x12c  :    8 - 0x8
    "00001000", --  301 - 0x12d  :    8 - 0x8
    "00001000", --  302 - 0x12e  :    8 - 0x8
    "00001000", --  303 - 0x12f  :    8 - 0x8
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Background 0x26
    "01111000", --  305 - 0x131  :  120 - 0x78
    "01100101", --  306 - 0x132  :  101 - 0x65
    "01111001", --  307 - 0x133  :  121 - 0x79
    "01100101", --  308 - 0x134  :  101 - 0x65
    "01100101", --  309 - 0x135  :  101 - 0x65
    "01111000", --  310 - 0x136  :  120 - 0x78
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Background 0x27
    "11100100", --  313 - 0x139  :  228 - 0xe4
    "10010110", --  314 - 0x13a  :  150 - 0x96
    "10010110", --  315 - 0x13b  :  150 - 0x96
    "10010111", --  316 - 0x13c  :  151 - 0x97
    "10010110", --  317 - 0x13d  :  150 - 0x96
    "11100110", --  318 - 0x13e  :  230 - 0xe6
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "01011001", --  321 - 0x141  :   89 - 0x59
    "01011001", --  322 - 0x142  :   89 - 0x59
    "01011001", --  323 - 0x143  :   89 - 0x59
    "01011001", --  324 - 0x144  :   89 - 0x59
    "11011001", --  325 - 0x145  :  217 - 0xd9
    "01001110", --  326 - 0x146  :   78 - 0x4e
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Background 0x29
    "00111100", --  329 - 0x149  :   60 - 0x3c
    "01110000", --  330 - 0x14a  :  112 - 0x70
    "01110000", --  331 - 0x14b  :  112 - 0x70
    "00111100", --  332 - 0x14c  :   60 - 0x3c
    "00001100", --  333 - 0x14d  :   12 - 0xc
    "01111000", --  334 - 0x14e  :  120 - 0x78
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Background 0x2a
    "00000000", --  337 - 0x151  :    0 - 0x0
    "11000110", --  338 - 0x152  :  198 - 0xc6
    "11101110", --  339 - 0x153  :  238 - 0xee
    "00101000", --  340 - 0x154  :   40 - 0x28
    "00101000", --  341 - 0x155  :   40 - 0x28
    "00101000", --  342 - 0x156  :   40 - 0x28
    "00101000", --  343 - 0x157  :   40 - 0x28
    "00001000", --  344 - 0x158  :    8 - 0x8 -- Background 0x2b
    "00001000", --  345 - 0x159  :    8 - 0x8
    "00001000", --  346 - 0x15a  :    8 - 0x8
    "00001000", --  347 - 0x15b  :    8 - 0x8
    "00001110", --  348 - 0x15c  :   14 - 0xe
    "00000110", --  349 - 0x15d  :    6 - 0x6
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00101000", --  352 - 0x160  :   40 - 0x28 -- Background 0x2c
    "00101000", --  353 - 0x161  :   40 - 0x28
    "00101000", --  354 - 0x162  :   40 - 0x28
    "00101000", --  355 - 0x163  :   40 - 0x28
    "11101110", --  356 - 0x164  :  238 - 0xee
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Background 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "01100000", --  362 - 0x16a  :   96 - 0x60
    "01110000", --  363 - 0x16b  :  112 - 0x70
    "00010000", --  364 - 0x16c  :   16 - 0x10
    "00010000", --  365 - 0x16d  :   16 - 0x10
    "00010000", --  366 - 0x16e  :   16 - 0x10
    "00010000", --  367 - 0x16f  :   16 - 0x10
    "00011100", --  368 - 0x170  :   28 - 0x1c -- Background 0x2e
    "00111110", --  369 - 0x171  :   62 - 0x3e
    "00111100", --  370 - 0x172  :   60 - 0x3c
    "00111000", --  371 - 0x173  :   56 - 0x38
    "00110000", --  372 - 0x174  :   48 - 0x30
    "00000000", --  373 - 0x175  :    0 - 0x0
    "01100000", --  374 - 0x176  :   96 - 0x60
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00010000", --  376 - 0x178  :   16 - 0x10 -- Background 0x2f
    "00010000", --  377 - 0x179  :   16 - 0x10
    "00010000", --  378 - 0x17a  :   16 - 0x10
    "00010000", --  379 - 0x17b  :   16 - 0x10
    "01110000", --  380 - 0x17c  :  112 - 0x70
    "01100000", --  381 - 0x17d  :   96 - 0x60
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "11111111", --  384 - 0x180  :  255 - 0xff -- Background 0x30
    "11111111", --  385 - 0x181  :  255 - 0xff
    "00111000", --  386 - 0x182  :   56 - 0x38
    "01101100", --  387 - 0x183  :  108 - 0x6c
    "11000110", --  388 - 0x184  :  198 - 0xc6
    "10000011", --  389 - 0x185  :  131 - 0x83
    "11111111", --  390 - 0x186  :  255 - 0xff
    "11111111", --  391 - 0x187  :  255 - 0xff
    "11111111", --  392 - 0x188  :  255 - 0xff -- Background 0x31
    "00111000", --  393 - 0x189  :   56 - 0x38
    "01101100", --  394 - 0x18a  :  108 - 0x6c
    "11000110", --  395 - 0x18b  :  198 - 0xc6
    "10000011", --  396 - 0x18c  :  131 - 0x83
    "11111111", --  397 - 0x18d  :  255 - 0xff
    "11111111", --  398 - 0x18e  :  255 - 0xff
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00111000", --  400 - 0x190  :   56 - 0x38 -- Background 0x32
    "01101100", --  401 - 0x191  :  108 - 0x6c
    "11000110", --  402 - 0x192  :  198 - 0xc6
    "10000011", --  403 - 0x193  :  131 - 0x83
    "11111111", --  404 - 0x194  :  255 - 0xff
    "11111111", --  405 - 0x195  :  255 - 0xff
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "01101100", --  408 - 0x198  :  108 - 0x6c -- Background 0x33
    "11000110", --  409 - 0x199  :  198 - 0xc6
    "10000011", --  410 - 0x19a  :  131 - 0x83
    "11111111", --  411 - 0x19b  :  255 - 0xff
    "11111111", --  412 - 0x19c  :  255 - 0xff
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "11000110", --  416 - 0x1a0  :  198 - 0xc6 -- Background 0x34
    "10000011", --  417 - 0x1a1  :  131 - 0x83
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111111", --  419 - 0x1a3  :  255 - 0xff
    "00000000", --  420 - 0x1a4  :    0 - 0x0
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "10000011", --  424 - 0x1a8  :  131 - 0x83 -- Background 0x35
    "11111111", --  425 - 0x1a9  :  255 - 0xff
    "11111111", --  426 - 0x1aa  :  255 - 0xff
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "11111111", --  432 - 0x1b0  :  255 - 0xff -- Background 0x36
    "11111111", --  433 - 0x1b1  :  255 - 0xff
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "00000000", --  437 - 0x1b5  :    0 - 0x0
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "11111111", --  440 - 0x1b8  :  255 - 0xff -- Background 0x37
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "11111111", --  455 - 0x1c7  :  255 - 0xff
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Background 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "11111111", --  462 - 0x1ce  :  255 - 0xff
    "11111111", --  463 - 0x1cf  :  255 - 0xff
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "11111111", --  470 - 0x1d6  :  255 - 0xff
    "00111000", --  471 - 0x1d7  :   56 - 0x38
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "11111111", --  476 - 0x1dc  :  255 - 0xff
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "00111000", --  478 - 0x1de  :   56 - 0x38
    "01101100", --  479 - 0x1df  :  108 - 0x6c
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "00111000", --  485 - 0x1e5  :   56 - 0x38
    "01101100", --  486 - 0x1e6  :  108 - 0x6c
    "11000110", --  487 - 0x1e7  :  198 - 0xc6
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "11111111", --  490 - 0x1ea  :  255 - 0xff
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "00111000", --  492 - 0x1ec  :   56 - 0x38
    "01101100", --  493 - 0x1ed  :  108 - 0x6c
    "11000110", --  494 - 0x1ee  :  198 - 0xc6
    "10000011", --  495 - 0x1ef  :  131 - 0x83
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "00111000", --  499 - 0x1f3  :   56 - 0x38
    "01101100", --  500 - 0x1f4  :  108 - 0x6c
    "11000110", --  501 - 0x1f5  :  198 - 0xc6
    "10000011", --  502 - 0x1f6  :  131 - 0x83
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Background 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "11111111", --  519 - 0x207  :  255 - 0xff
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Background 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "11111111", --  525 - 0x20d  :  255 - 0xff
    "11111111", --  526 - 0x20e  :  255 - 0xff
    "00111000", --  527 - 0x20f  :   56 - 0x38
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Background 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111111", --  533 - 0x215  :  255 - 0xff
    "00111000", --  534 - 0x216  :   56 - 0x38
    "01101100", --  535 - 0x217  :  108 - 0x6c
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Background 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "00111000", --  541 - 0x21d  :   56 - 0x38
    "01101100", --  542 - 0x21e  :  108 - 0x6c
    "11000110", --  543 - 0x21f  :  198 - 0xc6
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Background 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111111", --  547 - 0x223  :  255 - 0xff
    "00111000", --  548 - 0x224  :   56 - 0x38
    "01101100", --  549 - 0x225  :  108 - 0x6c
    "11000110", --  550 - 0x226  :  198 - 0xc6
    "10000011", --  551 - 0x227  :  131 - 0x83
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Background 0x45
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "00111000", --  555 - 0x22b  :   56 - 0x38
    "01101100", --  556 - 0x22c  :  108 - 0x6c
    "11000110", --  557 - 0x22d  :  198 - 0xc6
    "10000011", --  558 - 0x22e  :  131 - 0x83
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "11111111", --  560 - 0x230  :  255 - 0xff -- Background 0x46
    "00111000", --  561 - 0x231  :   56 - 0x38
    "01101100", --  562 - 0x232  :  108 - 0x6c
    "11000110", --  563 - 0x233  :  198 - 0xc6
    "10000011", --  564 - 0x234  :  131 - 0x83
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00111000", --  568 - 0x238  :   56 - 0x38 -- Background 0x47
    "01101100", --  569 - 0x239  :  108 - 0x6c
    "11000110", --  570 - 0x23a  :  198 - 0xc6
    "10000011", --  571 - 0x23b  :  131 - 0x83
    "11111111", --  572 - 0x23c  :  255 - 0xff
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "01101100", --  576 - 0x240  :  108 - 0x6c -- Background 0x48
    "11000110", --  577 - 0x241  :  198 - 0xc6
    "10000011", --  578 - 0x242  :  131 - 0x83
    "11111111", --  579 - 0x243  :  255 - 0xff
    "11111111", --  580 - 0x244  :  255 - 0xff
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "11000110", --  584 - 0x248  :  198 - 0xc6 -- Background 0x49
    "10000011", --  585 - 0x249  :  131 - 0x83
    "11111111", --  586 - 0x24a  :  255 - 0xff
    "11111111", --  587 - 0x24b  :  255 - 0xff
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "10000011", --  592 - 0x250  :  131 - 0x83 -- Background 0x4a
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "11111111", --  600 - 0x258  :  255 - 0xff -- Background 0x4b
    "11111111", --  601 - 0x259  :  255 - 0xff
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "10111111", --  608 - 0x260  :  191 - 0xbf -- Background 0x4c
    "01011111", --  609 - 0x261  :   95 - 0x5f
    "01011111", --  610 - 0x262  :   95 - 0x5f
    "01011111", --  611 - 0x263  :   95 - 0x5f
    "00000000", --  612 - 0x264  :    0 - 0x0
    "01011111", --  613 - 0x265  :   95 - 0x5f
    "01010001", --  614 - 0x266  :   81 - 0x51
    "01010101", --  615 - 0x267  :   85 - 0x55
    "01010001", --  616 - 0x268  :   81 - 0x51 -- Background 0x4d
    "01011111", --  617 - 0x269  :   95 - 0x5f
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "01011111", --  619 - 0x26b  :   95 - 0x5f
    "01011111", --  620 - 0x26c  :   95 - 0x5f
    "01011111", --  621 - 0x26d  :   95 - 0x5f
    "01011111", --  622 - 0x26e  :   95 - 0x5f
    "10111111", --  623 - 0x26f  :  191 - 0xbf
    "11111111", --  624 - 0x270  :  255 - 0xff -- Background 0x4e
    "11111110", --  625 - 0x271  :  254 - 0xfe
    "11111110", --  626 - 0x272  :  254 - 0xfe
    "11111110", --  627 - 0x273  :  254 - 0xfe
    "00000000", --  628 - 0x274  :    0 - 0x0
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "00100110", --  630 - 0x276  :   38 - 0x26
    "00100110", --  631 - 0x277  :   38 - 0x26
    "00100010", --  632 - 0x278  :   34 - 0x22 -- Background 0x4f
    "11111110", --  633 - 0x279  :  254 - 0xfe
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "11111110", --  636 - 0x27c  :  254 - 0xfe
    "11111110", --  637 - 0x27d  :  254 - 0xfe
    "11111110", --  638 - 0x27e  :  254 - 0xfe
    "11111111", --  639 - 0x27f  :  255 - 0xff
    "00000111", --  640 - 0x280  :    7 - 0x7 -- Background 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00001111", --  642 - 0x282  :   15 - 0xf
    "00011111", --  643 - 0x283  :   31 - 0x1f
    "00011111", --  644 - 0x284  :   31 - 0x1f
    "00011111", --  645 - 0x285  :   31 - 0x1f
    "00011111", --  646 - 0x286  :   31 - 0x1f
    "00011111", --  647 - 0x287  :   31 - 0x1f
    "00011111", --  648 - 0x288  :   31 - 0x1f -- Background 0x51
    "00011111", --  649 - 0x289  :   31 - 0x1f
    "00011111", --  650 - 0x28a  :   31 - 0x1f
    "00011111", --  651 - 0x28b  :   31 - 0x1f
    "00011111", --  652 - 0x28c  :   31 - 0x1f
    "00001111", --  653 - 0x28d  :   15 - 0xf
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000111", --  655 - 0x28f  :    7 - 0x7
    "00000111", --  656 - 0x290  :    7 - 0x7 -- Background 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00001111", --  658 - 0x292  :   15 - 0xf
    "00011111", --  659 - 0x293  :   31 - 0x1f
    "00011111", --  660 - 0x294  :   31 - 0x1f
    "00011111", --  661 - 0x295  :   31 - 0x1f
    "00011111", --  662 - 0x296  :   31 - 0x1f
    "00011111", --  663 - 0x297  :   31 - 0x1f
    "00011111", --  664 - 0x298  :   31 - 0x1f -- Background 0x53
    "00011111", --  665 - 0x299  :   31 - 0x1f
    "00011111", --  666 - 0x29a  :   31 - 0x1f
    "00011111", --  667 - 0x29b  :   31 - 0x1f
    "00011111", --  668 - 0x29c  :   31 - 0x1f
    "00001111", --  669 - 0x29d  :   15 - 0xf
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000111", --  671 - 0x29f  :    7 - 0x7
    "11100000", --  672 - 0x2a0  :  224 - 0xe0 -- Background 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "11110001", --  674 - 0x2a2  :  241 - 0xf1
    "11111011", --  675 - 0x2a3  :  251 - 0xfb
    "11111011", --  676 - 0x2a4  :  251 - 0xfb
    "11111011", --  677 - 0x2a5  :  251 - 0xfb
    "11111011", --  678 - 0x2a6  :  251 - 0xfb
    "11111011", --  679 - 0x2a7  :  251 - 0xfb
    "11111011", --  680 - 0x2a8  :  251 - 0xfb -- Background 0x55
    "11111011", --  681 - 0x2a9  :  251 - 0xfb
    "11111011", --  682 - 0x2aa  :  251 - 0xfb
    "11111011", --  683 - 0x2ab  :  251 - 0xfb
    "11111011", --  684 - 0x2ac  :  251 - 0xfb
    "11110001", --  685 - 0x2ad  :  241 - 0xf1
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "11100000", --  687 - 0x2af  :  224 - 0xe0
    "11100000", --  688 - 0x2b0  :  224 - 0xe0 -- Background 0x56
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "11110001", --  690 - 0x2b2  :  241 - 0xf1
    "11111011", --  691 - 0x2b3  :  251 - 0xfb
    "11111011", --  692 - 0x2b4  :  251 - 0xfb
    "11111011", --  693 - 0x2b5  :  251 - 0xfb
    "11111011", --  694 - 0x2b6  :  251 - 0xfb
    "11111011", --  695 - 0x2b7  :  251 - 0xfb
    "11111011", --  696 - 0x2b8  :  251 - 0xfb -- Background 0x57
    "11111011", --  697 - 0x2b9  :  251 - 0xfb
    "11111011", --  698 - 0x2ba  :  251 - 0xfb
    "11111011", --  699 - 0x2bb  :  251 - 0xfb
    "11111011", --  700 - 0x2bc  :  251 - 0xfb
    "11110001", --  701 - 0x2bd  :  241 - 0xf1
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "11100000", --  703 - 0x2bf  :  224 - 0xe0
    "11111100", --  704 - 0x2c0  :  252 - 0xfc -- Background 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "11111110", --  706 - 0x2c2  :  254 - 0xfe
    "11111111", --  707 - 0x2c3  :  255 - 0xff
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11111111", --  710 - 0x2c6  :  255 - 0xff
    "11111111", --  711 - 0x2c7  :  255 - 0xff
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- Background 0x59
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "11111111", --  714 - 0x2ca  :  255 - 0xff
    "11111111", --  715 - 0x2cb  :  255 - 0xff
    "11111111", --  716 - 0x2cc  :  255 - 0xff
    "11111110", --  717 - 0x2cd  :  254 - 0xfe
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "11111100", --  719 - 0x2cf  :  252 - 0xfc
    "11111100", --  720 - 0x2d0  :  252 - 0xfc -- Background 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "11111110", --  722 - 0x2d2  :  254 - 0xfe
    "11111111", --  723 - 0x2d3  :  255 - 0xff
    "11111111", --  724 - 0x2d4  :  255 - 0xff
    "11111111", --  725 - 0x2d5  :  255 - 0xff
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "11111111", --  728 - 0x2d8  :  255 - 0xff -- Background 0x5b
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111110", --  733 - 0x2dd  :  254 - 0xfe
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "11111100", --  735 - 0x2df  :  252 - 0xfc
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00011111", --  738 - 0x2e2  :   31 - 0x1f
    "00010000", --  739 - 0x2e3  :   16 - 0x10
    "00010000", --  740 - 0x2e4  :   16 - 0x10
    "00011111", --  741 - 0x2e5  :   31 - 0x1f
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Background 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "11111000", --  746 - 0x2ea  :  248 - 0xf8
    "00001000", --  747 - 0x2eb  :    8 - 0x8
    "00001000", --  748 - 0x2ec  :    8 - 0x8
    "11111000", --  749 - 0x2ed  :  248 - 0xf8
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00000001", --  753 - 0x2f1  :    1 - 0x1
    "00000010", --  754 - 0x2f2  :    2 - 0x2
    "00000010", --  755 - 0x2f3  :    2 - 0x2
    "11110001", --  756 - 0x2f4  :  241 - 0xf1
    "00001000", --  757 - 0x2f5  :    8 - 0x8
    "00000100", --  758 - 0x2f6  :    4 - 0x4
    "00000011", --  759 - 0x2f7  :    3 - 0x3
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Background 0x5f
    "10000000", --  761 - 0x2f9  :  128 - 0x80
    "01000000", --  762 - 0x2fa  :   64 - 0x40
    "01000000", --  763 - 0x2fb  :   64 - 0x40
    "10001111", --  764 - 0x2fc  :  143 - 0x8f
    "00010000", --  765 - 0x2fd  :   16 - 0x10
    "00100000", --  766 - 0x2fe  :   32 - 0x20
    "11000000", --  767 - 0x2ff  :  192 - 0xc0
    "00000011", --  768 - 0x300  :    3 - 0x3 -- Background 0x60
    "00000100", --  769 - 0x301  :    4 - 0x4
    "00001000", --  770 - 0x302  :    8 - 0x8
    "11110001", --  771 - 0x303  :  241 - 0xf1
    "00000010", --  772 - 0x304  :    2 - 0x2
    "00000010", --  773 - 0x305  :    2 - 0x2
    "00000001", --  774 - 0x306  :    1 - 0x1
    "00000000", --  775 - 0x307  :    0 - 0x0
    "11000000", --  776 - 0x308  :  192 - 0xc0 -- Background 0x61
    "00100000", --  777 - 0x309  :   32 - 0x20
    "00010000", --  778 - 0x30a  :   16 - 0x10
    "10001111", --  779 - 0x30b  :  143 - 0x8f
    "01000000", --  780 - 0x30c  :   64 - 0x40
    "01000000", --  781 - 0x30d  :   64 - 0x40
    "10000000", --  782 - 0x30e  :  128 - 0x80
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "11111111", --  784 - 0x310  :  255 - 0xff -- Background 0x62
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11000011", --  786 - 0x312  :  195 - 0xc3
    "10000001", --  787 - 0x313  :  129 - 0x81
    "10000001", --  788 - 0x314  :  129 - 0x81
    "11000011", --  789 - 0x315  :  195 - 0xc3
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff -- Background 0x63
    "10011001", --  793 - 0x319  :  153 - 0x99
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "10000001", --  797 - 0x31d  :  129 - 0x81
    "10000001", --  798 - 0x31e  :  129 - 0x81
    "10000001", --  799 - 0x31f  :  129 - 0x81
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "01100000", --  804 - 0x324  :   96 - 0x60
    "01100000", --  805 - 0x325  :   96 - 0x60
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Background 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "01101100", --  812 - 0x32c  :  108 - 0x6c
    "01101100", --  813 - 0x32d  :  108 - 0x6c
    "00001000", --  814 - 0x32e  :    8 - 0x8
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00111100", --  816 - 0x330  :   60 - 0x3c -- Background 0x66
    "00011000", --  817 - 0x331  :   24 - 0x18
    "00011000", --  818 - 0x332  :   24 - 0x18
    "00011000", --  819 - 0x333  :   24 - 0x18
    "00011000", --  820 - 0x334  :   24 - 0x18
    "00011000", --  821 - 0x335  :   24 - 0x18
    "00111100", --  822 - 0x336  :   60 - 0x3c
    "00000000", --  823 - 0x337  :    0 - 0x0
    "11111111", --  824 - 0x338  :  255 - 0xff -- Background 0x67
    "01100110", --  825 - 0x339  :  102 - 0x66
    "01100110", --  826 - 0x33a  :  102 - 0x66
    "01100110", --  827 - 0x33b  :  102 - 0x66
    "01100110", --  828 - 0x33c  :  102 - 0x66
    "01100110", --  829 - 0x33d  :  102 - 0x66
    "01100110", --  830 - 0x33e  :  102 - 0x66
    "11111111", --  831 - 0x33f  :  255 - 0xff
    "00000011", --  832 - 0x340  :    3 - 0x3 -- Background 0x68
    "00000001", --  833 - 0x341  :    1 - 0x1
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "10000011", --  840 - 0x348  :  131 - 0x83 -- Background 0x69
    "11010001", --  841 - 0x349  :  209 - 0xd1
    "11100001", --  842 - 0x34a  :  225 - 0xe1
    "11010001", --  843 - 0x34b  :  209 - 0xd1
    "00000010", --  844 - 0x34c  :    2 - 0x2
    "10000100", --  845 - 0x34d  :  132 - 0x84
    "11110000", --  846 - 0x34e  :  240 - 0xf0
    "11001110", --  847 - 0x34f  :  206 - 0xce
    "11000000", --  848 - 0x350  :  192 - 0xc0 -- Background 0x6a
    "10000000", --  849 - 0x351  :  128 - 0x80
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "11000001", --  856 - 0x358  :  193 - 0xc1 -- Background 0x6b
    "10001011", --  857 - 0x359  :  139 - 0x8b
    "10000111", --  858 - 0x35a  :  135 - 0x87
    "10001011", --  859 - 0x35b  :  139 - 0x8b
    "01000000", --  860 - 0x35c  :   64 - 0x40
    "00100001", --  861 - 0x35d  :   33 - 0x21
    "00001111", --  862 - 0x35e  :   15 - 0xf
    "11010011", --  863 - 0x35f  :  211 - 0xd3
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "00011111", --  867 - 0x363  :   31 - 0x1f
    "00001111", --  868 - 0x364  :   15 - 0xf
    "00011110", --  869 - 0x365  :   30 - 0x1e
    "00111111", --  870 - 0x366  :   63 - 0x3f
    "01111111", --  871 - 0x367  :  127 - 0x7f
    "11111111", --  872 - 0x368  :  255 - 0xff -- Background 0x6d
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111000", --  875 - 0x36b  :  248 - 0xf8
    "11110000", --  876 - 0x36c  :  240 - 0xf0
    "01111000", --  877 - 0x36d  :  120 - 0x78
    "11111100", --  878 - 0x36e  :  252 - 0xfc
    "11111110", --  879 - 0x36f  :  254 - 0xfe
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00111100", --  885 - 0x375  :   60 - 0x3c
    "01000010", --  886 - 0x376  :   66 - 0x42
    "10000001", --  887 - 0x377  :  129 - 0x81
    "10000001", --  888 - 0x378  :  129 - 0x81 -- Background 0x6f
    "10111101", --  889 - 0x379  :  189 - 0xbd
    "01111110", --  890 - 0x37a  :  126 - 0x7e
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11100111", --  892 - 0x37c  :  231 - 0xe7
    "11111111", --  893 - 0x37d  :  255 - 0xff
    "11111111", --  894 - 0x37e  :  255 - 0xff
    "11111111", --  895 - 0x37f  :  255 - 0xff
    "00000001", --  896 - 0x380  :    1 - 0x1 -- Background 0x70
    "00000111", --  897 - 0x381  :    7 - 0x7
    "00011111", --  898 - 0x382  :   31 - 0x1f
    "00111111", --  899 - 0x383  :   63 - 0x3f
    "01111111", --  900 - 0x384  :  127 - 0x7f
    "11111111", --  901 - 0x385  :  255 - 0xff
    "11111111", --  902 - 0x386  :  255 - 0xff
    "11011101", --  903 - 0x387  :  221 - 0xdd
    "10001001", --  904 - 0x388  :  137 - 0x89 -- Background 0x71
    "00000001", --  905 - 0x389  :    1 - 0x1
    "00000001", --  906 - 0x38a  :    1 - 0x1
    "00000001", --  907 - 0x38b  :    1 - 0x1
    "00000001", --  908 - 0x38c  :    1 - 0x1
    "00000001", --  909 - 0x38d  :    1 - 0x1
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "10000000", --  912 - 0x390  :  128 - 0x80 -- Background 0x72
    "11100000", --  913 - 0x391  :  224 - 0xe0
    "11111000", --  914 - 0x392  :  248 - 0xf8
    "11111100", --  915 - 0x393  :  252 - 0xfc
    "11111110", --  916 - 0x394  :  254 - 0xfe
    "11111111", --  917 - 0x395  :  255 - 0xff
    "11111111", --  918 - 0x396  :  255 - 0xff
    "00111011", --  919 - 0x397  :   59 - 0x3b
    "00010001", --  920 - 0x398  :   17 - 0x11 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "01000000", --  925 - 0x39d  :   64 - 0x40
    "10000000", --  926 - 0x39e  :  128 - 0x80
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000001", --  928 - 0x3a0  :    1 - 0x1 -- Background 0x74
    "00000001", --  929 - 0x3a1  :    1 - 0x1
    "00000001", --  930 - 0x3a2  :    1 - 0x1
    "00000001", --  931 - 0x3a3  :    1 - 0x1
    "00000001", --  932 - 0x3a4  :    1 - 0x1
    "00000001", --  933 - 0x3a5  :    1 - 0x1
    "00000001", --  934 - 0x3a6  :    1 - 0x1
    "00000001", --  935 - 0x3a7  :    1 - 0x1
    "10000000", --  936 - 0x3a8  :  128 - 0x80 -- Background 0x75
    "10000000", --  937 - 0x3a9  :  128 - 0x80
    "10000000", --  938 - 0x3aa  :  128 - 0x80
    "10000000", --  939 - 0x3ab  :  128 - 0x80
    "10000000", --  940 - 0x3ac  :  128 - 0x80
    "10000000", --  941 - 0x3ad  :  128 - 0x80
    "10000000", --  942 - 0x3ae  :  128 - 0x80
    "10000000", --  943 - 0x3af  :  128 - 0x80
    "00000001", --  944 - 0x3b0  :    1 - 0x1 -- Background 0x76
    "00000011", --  945 - 0x3b1  :    3 - 0x3
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000011", --  948 - 0x3b4  :    3 - 0x3
    "00011001", --  949 - 0x3b5  :   25 - 0x19
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Background 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "01111100", --  954 - 0x3ba  :  124 - 0x7c
    "00000010", --  955 - 0x3bb  :    2 - 0x2
    "00000001", --  956 - 0x3bc  :    1 - 0x1
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000001", --  962 - 0x3c2  :    1 - 0x1
    "00000001", --  963 - 0x3c3  :    1 - 0x1
    "00000011", --  964 - 0x3c4  :    3 - 0x3
    "00000111", --  965 - 0x3c5  :    7 - 0x7
    "00000111", --  966 - 0x3c6  :    7 - 0x7
    "00001111", --  967 - 0x3c7  :   15 - 0xf
    "00001111", --  968 - 0x3c8  :   15 - 0xf -- Background 0x79
    "00000111", --  969 - 0x3c9  :    7 - 0x7
    "00001111", --  970 - 0x3ca  :   15 - 0xf
    "00000111", --  971 - 0x3cb  :    7 - 0x7
    "00000001", --  972 - 0x3cc  :    1 - 0x1
    "00010000", --  973 - 0x3cd  :   16 - 0x10
    "00100000", --  974 - 0x3ce  :   32 - 0x20
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "11111000", --  976 - 0x3d0  :  248 - 0xf8 -- Background 0x7a
    "11111110", --  977 - 0x3d1  :  254 - 0xfe
    "01111111", --  978 - 0x3d2  :  127 - 0x7f
    "00011111", --  979 - 0x3d3  :   31 - 0x1f
    "00001111", --  980 - 0x3d4  :   15 - 0xf
    "00011001", --  981 - 0x3d5  :   25 - 0x19
    "00110000", --  982 - 0x3d6  :   48 - 0x30
    "01110000", --  983 - 0x3d7  :  112 - 0x70
    "11111011", --  984 - 0x3d8  :  251 - 0xfb -- Background 0x7b
    "01110011", --  985 - 0x3d9  :  115 - 0x73
    "00100111", --  986 - 0x3da  :   39 - 0x27
    "00001111", --  987 - 0x3db  :   15 - 0xf
    "00011111", --  988 - 0x3dc  :   31 - 0x1f
    "00011111", --  989 - 0x3dd  :   31 - 0x1f
    "00111111", --  990 - 0x3de  :   63 - 0x3f
    "01111111", --  991 - 0x3df  :  127 - 0x7f
    "11111111", --  992 - 0x3e0  :  255 - 0xff -- Background 0x7c
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111110", --  996 - 0x3e4  :  254 - 0xfe
    "11111101", --  997 - 0x3e5  :  253 - 0xfd
    "11111000", --  998 - 0x3e6  :  248 - 0xf8
    "11110110", --  999 - 0x3e7  :  246 - 0xf6
    "11101111", -- 1000 - 0x3e8  :  239 - 0xef -- Background 0x7d
    "11001111", -- 1001 - 0x3e9  :  207 - 0xcf
    "10011111", -- 1002 - 0x3ea  :  159 - 0x9f
    "00011111", -- 1003 - 0x3eb  :   31 - 0x1f
    "00001111", -- 1004 - 0x3ec  :   15 - 0xf
    "00101101", -- 1005 - 0x3ed  :   45 - 0x2d
    "01010000", -- 1006 - 0x3ee  :   80 - 0x50
    "01000000", -- 1007 - 0x3ef  :   64 - 0x40
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "11100000", -- 1012 - 0x3f4  :  224 - 0xe0
    "11111110", -- 1013 - 0x3f5  :  254 - 0xfe
    "11111111", -- 1014 - 0x3f6  :  255 - 0xff
    "11110011", -- 1015 - 0x3f7  :  243 - 0xf3
    "11111011", -- 1016 - 0x3f8  :  251 - 0xfb -- Background 0x7f
    "11111011", -- 1017 - 0x3f9  :  251 - 0xfb
    "11111011", -- 1018 - 0x3fa  :  251 - 0xfb
    "11111011", -- 1019 - 0x3fb  :  251 - 0xfb
    "11111011", -- 1020 - 0x3fc  :  251 - 0xfb
    "11110011", -- 1021 - 0x3fd  :  243 - 0xf3
    "11110111", -- 1022 - 0x3fe  :  247 - 0xf7
    "11100111", -- 1023 - 0x3ff  :  231 - 0xe7
    "11001111", -- 1024 - 0x400  :  207 - 0xcf -- Background 0x80
    "10011111", -- 1025 - 0x401  :  159 - 0x9f
    "00111111", -- 1026 - 0x402  :   63 - 0x3f
    "00111111", -- 1027 - 0x403  :   63 - 0x3f
    "00111111", -- 1028 - 0x404  :   63 - 0x3f
    "00001111", -- 1029 - 0x405  :   15 - 0xf
    "00000011", -- 1030 - 0x406  :    3 - 0x3
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "11000000", -- 1032 - 0x408  :  192 - 0xc0 -- Background 0x81
    "11110000", -- 1033 - 0x409  :  240 - 0xf0
    "11111100", -- 1034 - 0x40a  :  252 - 0xfc
    "11110000", -- 1035 - 0x40b  :  240 - 0xf0
    "11110000", -- 1036 - 0x40c  :  240 - 0xf0
    "10011000", -- 1037 - 0x40d  :  152 - 0x98
    "00001000", -- 1038 - 0x40e  :    8 - 0x8
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x82
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "10000000", -- 1046 - 0x416  :  128 - 0x80
    "11000000", -- 1047 - 0x417  :  192 - 0xc0
    "11100000", -- 1048 - 0x418  :  224 - 0xe0 -- Background 0x83
    "11100000", -- 1049 - 0x419  :  224 - 0xe0
    "11110000", -- 1050 - 0x41a  :  240 - 0xf0
    "11110000", -- 1051 - 0x41b  :  240 - 0xf0
    "11110000", -- 1052 - 0x41c  :  240 - 0xf0
    "11110000", -- 1053 - 0x41d  :  240 - 0xf0
    "11111000", -- 1054 - 0x41e  :  248 - 0xf8
    "11111000", -- 1055 - 0x41f  :  248 - 0xf8
    "11111110", -- 1056 - 0x420  :  254 - 0xfe -- Background 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111111", -- 1061 - 0x425  :  255 - 0xff
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "00111111", -- 1064 - 0x428  :   63 - 0x3f -- Background 0x85
    "00011111", -- 1065 - 0x429  :   31 - 0x1f
    "00011111", -- 1066 - 0x42a  :   31 - 0x1f
    "00001111", -- 1067 - 0x42b  :   15 - 0xf
    "00000111", -- 1068 - 0x42c  :    7 - 0x7
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "11000000", -- 1074 - 0x432  :  192 - 0xc0
    "11100000", -- 1075 - 0x433  :  224 - 0xe0
    "11110000", -- 1076 - 0x434  :  240 - 0xf0
    "11110000", -- 1077 - 0x435  :  240 - 0xf0
    "11110000", -- 1078 - 0x436  :  240 - 0xf0
    "11111000", -- 1079 - 0x437  :  248 - 0xf8
    "11111001", -- 1080 - 0x438  :  249 - 0xf9 -- Background 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "00001110", -- 1085 - 0x43d  :   14 - 0xe
    "00000010", -- 1086 - 0x43e  :    2 - 0x2
    "00010100", -- 1087 - 0x43f  :   20 - 0x14
    "10000000", -- 1088 - 0x440  :  128 - 0x80 -- Background 0x88
    "10100000", -- 1089 - 0x441  :  160 - 0xa0
    "00100000", -- 1090 - 0x442  :   32 - 0x20
    "00100000", -- 1091 - 0x443  :   32 - 0x20
    "10100000", -- 1092 - 0x444  :  160 - 0xa0
    "10000000", -- 1093 - 0x445  :  128 - 0x80
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000001", -- 1096 - 0x448  :    1 - 0x1 -- Background 0x89
    "00000101", -- 1097 - 0x449  :    5 - 0x5
    "00000100", -- 1098 - 0x44a  :    4 - 0x4
    "00000100", -- 1099 - 0x44b  :    4 - 0x4
    "00000101", -- 1100 - 0x44c  :    5 - 0x5
    "00000001", -- 1101 - 0x44d  :    1 - 0x1
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000011", -- 1106 - 0x452  :    3 - 0x3
    "00000111", -- 1107 - 0x453  :    7 - 0x7
    "00001111", -- 1108 - 0x454  :   15 - 0xf
    "00001111", -- 1109 - 0x455  :   15 - 0xf
    "00001111", -- 1110 - 0x456  :   15 - 0xf
    "00001111", -- 1111 - 0x457  :   15 - 0xf
    "10011111", -- 1112 - 0x458  :  159 - 0x9f -- Background 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "01110000", -- 1117 - 0x45d  :  112 - 0x70
    "01000000", -- 1118 - 0x45e  :   64 - 0x40
    "00101000", -- 1119 - 0x45f  :   40 - 0x28
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000001", -- 1126 - 0x466  :    1 - 0x1
    "00000011", -- 1127 - 0x467  :    3 - 0x3
    "00000111", -- 1128 - 0x468  :    7 - 0x7 -- Background 0x8d
    "00000111", -- 1129 - 0x469  :    7 - 0x7
    "00001111", -- 1130 - 0x46a  :   15 - 0xf
    "00001111", -- 1131 - 0x46b  :   15 - 0xf
    "00001111", -- 1132 - 0x46c  :   15 - 0xf
    "00001111", -- 1133 - 0x46d  :   15 - 0xf
    "00011111", -- 1134 - 0x46e  :   31 - 0x1f
    "00011111", -- 1135 - 0x46f  :   31 - 0x1f
    "01111111", -- 1136 - 0x470  :  127 - 0x7f -- Background 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111111", -- 1138 - 0x472  :  255 - 0xff
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11111111", -- 1140 - 0x474  :  255 - 0xff
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "11111100", -- 1144 - 0x478  :  252 - 0xfc -- Background 0x8f
    "11111000", -- 1145 - 0x479  :  248 - 0xf8
    "11111000", -- 1146 - 0x47a  :  248 - 0xf8
    "11110000", -- 1147 - 0x47b  :  240 - 0xf0
    "11100000", -- 1148 - 0x47c  :  224 - 0xe0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000111", -- 1156 - 0x484  :    7 - 0x7
    "01111111", -- 1157 - 0x485  :  127 - 0x7f
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11001111", -- 1159 - 0x487  :  207 - 0xcf
    "11011111", -- 1160 - 0x488  :  223 - 0xdf -- Background 0x91
    "11011111", -- 1161 - 0x489  :  223 - 0xdf
    "11011111", -- 1162 - 0x48a  :  223 - 0xdf
    "11011111", -- 1163 - 0x48b  :  223 - 0xdf
    "11011111", -- 1164 - 0x48c  :  223 - 0xdf
    "11001111", -- 1165 - 0x48d  :  207 - 0xcf
    "11101111", -- 1166 - 0x48e  :  239 - 0xef
    "11100111", -- 1167 - 0x48f  :  231 - 0xe7
    "11110011", -- 1168 - 0x490  :  243 - 0xf3 -- Background 0x92
    "11111001", -- 1169 - 0x491  :  249 - 0xf9
    "11111100", -- 1170 - 0x492  :  252 - 0xfc
    "11111100", -- 1171 - 0x493  :  252 - 0xfc
    "11111100", -- 1172 - 0x494  :  252 - 0xfc
    "11110000", -- 1173 - 0x495  :  240 - 0xf0
    "11000000", -- 1174 - 0x496  :  192 - 0xc0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000011", -- 1176 - 0x498  :    3 - 0x3 -- Background 0x93
    "00001111", -- 1177 - 0x499  :   15 - 0xf
    "00111111", -- 1178 - 0x49a  :   63 - 0x3f
    "00001111", -- 1179 - 0x49b  :   15 - 0xf
    "00001111", -- 1180 - 0x49c  :   15 - 0xf
    "00011001", -- 1181 - 0x49d  :   25 - 0x19
    "00010000", -- 1182 - 0x49e  :   16 - 0x10
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00011111", -- 1184 - 0x4a0  :   31 - 0x1f -- Background 0x94
    "01111111", -- 1185 - 0x4a1  :  127 - 0x7f
    "11111110", -- 1186 - 0x4a2  :  254 - 0xfe
    "11111000", -- 1187 - 0x4a3  :  248 - 0xf8
    "11110000", -- 1188 - 0x4a4  :  240 - 0xf0
    "10011000", -- 1189 - 0x4a5  :  152 - 0x98
    "00001100", -- 1190 - 0x4a6  :   12 - 0xc
    "00001110", -- 1191 - 0x4a7  :   14 - 0xe
    "11011111", -- 1192 - 0x4a8  :  223 - 0xdf -- Background 0x95
    "11001110", -- 1193 - 0x4a9  :  206 - 0xce
    "11100100", -- 1194 - 0x4aa  :  228 - 0xe4
    "11110000", -- 1195 - 0x4ab  :  240 - 0xf0
    "11111000", -- 1196 - 0x4ac  :  248 - 0xf8
    "11111000", -- 1197 - 0x4ad  :  248 - 0xf8
    "11111100", -- 1198 - 0x4ae  :  252 - 0xfc
    "11111110", -- 1199 - 0x4af  :  254 - 0xfe
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Background 0x96
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "01111111", -- 1204 - 0x4b4  :  127 - 0x7f
    "10111111", -- 1205 - 0x4b5  :  191 - 0xbf
    "00011111", -- 1206 - 0x4b6  :   31 - 0x1f
    "01101111", -- 1207 - 0x4b7  :  111 - 0x6f
    "11110111", -- 1208 - 0x4b8  :  247 - 0xf7 -- Background 0x97
    "11110011", -- 1209 - 0x4b9  :  243 - 0xf3
    "11111001", -- 1210 - 0x4ba  :  249 - 0xf9
    "11111000", -- 1211 - 0x4bb  :  248 - 0xf8
    "11110000", -- 1212 - 0x4bc  :  240 - 0xf0
    "10110100", -- 1213 - 0x4bd  :  180 - 0xb4
    "00001010", -- 1214 - 0x4be  :   10 - 0xa
    "00000010", -- 1215 - 0x4bf  :    2 - 0x2
    "10000000", -- 1216 - 0x4c0  :  128 - 0x80 -- Background 0x98
    "11000000", -- 1217 - 0x4c1  :  192 - 0xc0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "11000000", -- 1220 - 0x4c4  :  192 - 0xc0
    "10011000", -- 1221 - 0x4c5  :  152 - 0x98
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00111110", -- 1226 - 0x4ca  :   62 - 0x3e
    "01000000", -- 1227 - 0x4cb  :   64 - 0x40
    "10000000", -- 1228 - 0x4cc  :  128 - 0x80
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "10000000", -- 1234 - 0x4d2  :  128 - 0x80
    "10000000", -- 1235 - 0x4d3  :  128 - 0x80
    "11000000", -- 1236 - 0x4d4  :  192 - 0xc0
    "11100000", -- 1237 - 0x4d5  :  224 - 0xe0
    "11100000", -- 1238 - 0x4d6  :  224 - 0xe0
    "11110000", -- 1239 - 0x4d7  :  240 - 0xf0
    "11110000", -- 1240 - 0x4d8  :  240 - 0xf0 -- Background 0x9b
    "11100000", -- 1241 - 0x4d9  :  224 - 0xe0
    "11110000", -- 1242 - 0x4da  :  240 - 0xf0
    "11100000", -- 1243 - 0x4db  :  224 - 0xe0
    "10000000", -- 1244 - 0x4dc  :  128 - 0x80
    "00001000", -- 1245 - 0x4dd  :    8 - 0x8
    "00000100", -- 1246 - 0x4de  :    4 - 0x4
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000001", -- 1250 - 0x4e2  :    1 - 0x1
    "00000011", -- 1251 - 0x4e3  :    3 - 0x3
    "00000011", -- 1252 - 0x4e4  :    3 - 0x3
    "00000011", -- 1253 - 0x4e5  :    3 - 0x3
    "00000111", -- 1254 - 0x4e6  :    7 - 0x7
    "00000111", -- 1255 - 0x4e7  :    7 - 0x7
    "00000111", -- 1256 - 0x4e8  :    7 - 0x7 -- Background 0x9d
    "00000011", -- 1257 - 0x4e9  :    3 - 0x3
    "00000011", -- 1258 - 0x4ea  :    3 - 0x3
    "00000011", -- 1259 - 0x4eb  :    3 - 0x3
    "00000011", -- 1260 - 0x4ec  :    3 - 0x3
    "00000011", -- 1261 - 0x4ed  :    3 - 0x3
    "00000011", -- 1262 - 0x4ee  :    3 - 0x3
    "00000001", -- 1263 - 0x4ef  :    1 - 0x1
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Background 0x9e
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000001", -- 1269 - 0x4f5  :    1 - 0x1
    "00000010", -- 1270 - 0x4f6  :    2 - 0x2
    "00000100", -- 1271 - 0x4f7  :    4 - 0x4
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00011100", -- 1278 - 0x4fe  :   28 - 0x1c
    "00111011", -- 1279 - 0x4ff  :   59 - 0x3b
    "01111110", -- 1280 - 0x500  :  126 - 0x7e -- Background 0xa0
    "11111110", -- 1281 - 0x501  :  254 - 0xfe
    "11111111", -- 1282 - 0x502  :  255 - 0xff
    "11111111", -- 1283 - 0x503  :  255 - 0xff
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111101", -- 1286 - 0x506  :  253 - 0xfd
    "11111001", -- 1287 - 0x507  :  249 - 0xf9
    "11110011", -- 1288 - 0x508  :  243 - 0xf3 -- Background 0xa1
    "11110111", -- 1289 - 0x509  :  247 - 0xf7
    "11110110", -- 1290 - 0x50a  :  246 - 0xf6
    "11101110", -- 1291 - 0x50b  :  238 - 0xee
    "11111101", -- 1292 - 0x50c  :  253 - 0xfd
    "11111100", -- 1293 - 0x50d  :  252 - 0xfc
    "11111000", -- 1294 - 0x50e  :  248 - 0xf8
    "11100001", -- 1295 - 0x50f  :  225 - 0xe1
    "11010011", -- 1296 - 0x510  :  211 - 0xd3 -- Background 0xa2
    "11001011", -- 1297 - 0x511  :  203 - 0xcb
    "11000011", -- 1298 - 0x512  :  195 - 0xc3
    "11100001", -- 1299 - 0x513  :  225 - 0xe1
    "11111001", -- 1300 - 0x514  :  249 - 0xf9
    "00111001", -- 1301 - 0x515  :   57 - 0x39
    "01000010", -- 1302 - 0x516  :   66 - 0x42
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000111", -- 1304 - 0x518  :    7 - 0x7 -- Background 0xa3
    "00001111", -- 1305 - 0x519  :   15 - 0xf
    "00011001", -- 1306 - 0x51a  :   25 - 0x19
    "00110000", -- 1307 - 0x51b  :   48 - 0x30
    "01100011", -- 1308 - 0x51c  :   99 - 0x63
    "01110010", -- 1309 - 0x51d  :  114 - 0x72
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "00000001", -- 1311 - 0x51f  :    1 - 0x1
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Background 0xa4
    "00011111", -- 1313 - 0x521  :   31 - 0x1f
    "00100000", -- 1314 - 0x522  :   32 - 0x20
    "11000000", -- 1315 - 0x523  :  192 - 0xc0
    "11000000", -- 1316 - 0x524  :  192 - 0xc0
    "11110000", -- 1317 - 0x525  :  240 - 0xf0
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11111111", -- 1319 - 0x527  :  255 - 0xff
    "10101011", -- 1320 - 0x528  :  171 - 0xab -- Background 0xa5
    "11000001", -- 1321 - 0x529  :  193 - 0xc1
    "10000001", -- 1322 - 0x52a  :  129 - 0x81
    "10010001", -- 1323 - 0x52b  :  145 - 0x91
    "10000010", -- 1324 - 0x52c  :  130 - 0x82
    "11111100", -- 1325 - 0x52d  :  252 - 0xfc
    "11100000", -- 1326 - 0x52e  :  224 - 0xe0
    "11001110", -- 1327 - 0x52f  :  206 - 0xce
    "11100101", -- 1328 - 0x530  :  229 - 0xe5 -- Background 0xa6
    "11011010", -- 1329 - 0x531  :  218 - 0xda
    "11110000", -- 1330 - 0x532  :  240 - 0xf0
    "11100000", -- 1331 - 0x533  :  224 - 0xe0
    "11000000", -- 1332 - 0x534  :  192 - 0xc0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "11110000", -- 1336 - 0x538  :  240 - 0xf0 -- Background 0xa7
    "11111000", -- 1337 - 0x539  :  248 - 0xf8
    "11001100", -- 1338 - 0x53a  :  204 - 0xcc
    "10000110", -- 1339 - 0x53b  :  134 - 0x86
    "01100010", -- 1340 - 0x53c  :   98 - 0x62
    "00100110", -- 1341 - 0x53d  :   38 - 0x26
    "00000110", -- 1342 - 0x53e  :    6 - 0x6
    "11000000", -- 1343 - 0x53f  :  192 - 0xc0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Background 0xa8
    "11111100", -- 1345 - 0x541  :  252 - 0xfc
    "00000110", -- 1346 - 0x542  :    6 - 0x6
    "00000011", -- 1347 - 0x543  :    3 - 0x3
    "00000001", -- 1348 - 0x544  :    1 - 0x1
    "00000111", -- 1349 - 0x545  :    7 - 0x7
    "11111111", -- 1350 - 0x546  :  255 - 0xff
    "11111111", -- 1351 - 0x547  :  255 - 0xff
    "11010101", -- 1352 - 0x548  :  213 - 0xd5 -- Background 0xa9
    "10000011", -- 1353 - 0x549  :  131 - 0x83
    "10000001", -- 1354 - 0x54a  :  129 - 0x81
    "10001001", -- 1355 - 0x54b  :  137 - 0x89
    "01000001", -- 1356 - 0x54c  :   65 - 0x41
    "00111111", -- 1357 - 0x54d  :   63 - 0x3f
    "00000111", -- 1358 - 0x54e  :    7 - 0x7
    "11010011", -- 1359 - 0x54f  :  211 - 0xd3
    "01101111", -- 1360 - 0x550  :  111 - 0x6f -- Background 0xaa
    "11011011", -- 1361 - 0x551  :  219 - 0xdb
    "00001111", -- 1362 - 0x552  :   15 - 0xf
    "00000111", -- 1363 - 0x553  :    7 - 0x7
    "00000011", -- 1364 - 0x554  :    3 - 0x3
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Background 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00111000", -- 1374 - 0x55e  :   56 - 0x38
    "11011100", -- 1375 - 0x55f  :  220 - 0xdc
    "01111110", -- 1376 - 0x560  :  126 - 0x7e -- Background 0xac
    "01111111", -- 1377 - 0x561  :  127 - 0x7f
    "01111111", -- 1378 - 0x562  :  127 - 0x7f
    "11111111", -- 1379 - 0x563  :  255 - 0xff
    "11111111", -- 1380 - 0x564  :  255 - 0xff
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "10111111", -- 1382 - 0x566  :  191 - 0xbf
    "10011111", -- 1383 - 0x567  :  159 - 0x9f
    "11001111", -- 1384 - 0x568  :  207 - 0xcf -- Background 0xad
    "11101111", -- 1385 - 0x569  :  239 - 0xef
    "01101111", -- 1386 - 0x56a  :  111 - 0x6f
    "01110111", -- 1387 - 0x56b  :  119 - 0x77
    "10111111", -- 1388 - 0x56c  :  191 - 0xbf
    "00111111", -- 1389 - 0x56d  :   63 - 0x3f
    "00011111", -- 1390 - 0x56e  :   31 - 0x1f
    "10000111", -- 1391 - 0x56f  :  135 - 0x87
    "11001011", -- 1392 - 0x570  :  203 - 0xcb -- Background 0xae
    "11010011", -- 1393 - 0x571  :  211 - 0xd3
    "11000011", -- 1394 - 0x572  :  195 - 0xc3
    "10000111", -- 1395 - 0x573  :  135 - 0x87
    "10011111", -- 1396 - 0x574  :  159 - 0x9f
    "10011100", -- 1397 - 0x575  :  156 - 0x9c
    "01000010", -- 1398 - 0x576  :   66 - 0x42
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "10000000", -- 1402 - 0x57a  :  128 - 0x80
    "11000000", -- 1403 - 0x57b  :  192 - 0xc0
    "11000000", -- 1404 - 0x57c  :  192 - 0xc0
    "11000000", -- 1405 - 0x57d  :  192 - 0xc0
    "11100000", -- 1406 - 0x57e  :  224 - 0xe0
    "11100000", -- 1407 - 0x57f  :  224 - 0xe0
    "11100000", -- 1408 - 0x580  :  224 - 0xe0 -- Background 0xb0
    "11000000", -- 1409 - 0x581  :  192 - 0xc0
    "11000000", -- 1410 - 0x582  :  192 - 0xc0
    "11000000", -- 1411 - 0x583  :  192 - 0xc0
    "11000000", -- 1412 - 0x584  :  192 - 0xc0
    "11000000", -- 1413 - 0x585  :  192 - 0xc0
    "11000000", -- 1414 - 0x586  :  192 - 0xc0
    "10000000", -- 1415 - 0x587  :  128 - 0x80
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "10000000", -- 1421 - 0x58d  :  128 - 0x80
    "01000000", -- 1422 - 0x58e  :   64 - 0x40
    "00100000", -- 1423 - 0x58f  :   32 - 0x20
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000001", -- 1427 - 0x593  :    1 - 0x1
    "00000011", -- 1428 - 0x594  :    3 - 0x3
    "00000111", -- 1429 - 0x595  :    7 - 0x7
    "00000111", -- 1430 - 0x596  :    7 - 0x7
    "00000111", -- 1431 - 0x597  :    7 - 0x7
    "00000011", -- 1432 - 0x598  :    3 - 0x3 -- Background 0xb3
    "00000001", -- 1433 - 0x599  :    1 - 0x1
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000001", -- 1438 - 0x59e  :    1 - 0x1
    "00000001", -- 1439 - 0x59f  :    1 - 0x1
    "00000001", -- 1440 - 0x5a0  :    1 - 0x1 -- Background 0xb4
    "00000001", -- 1441 - 0x5a1  :    1 - 0x1
    "00000111", -- 1442 - 0x5a2  :    7 - 0x7
    "00000011", -- 1443 - 0x5a3  :    3 - 0x3
    "00000100", -- 1444 - 0x5a4  :    4 - 0x4
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000111", -- 1455 - 0x5af  :    7 - 0x7
    "00001110", -- 1456 - 0x5b0  :   14 - 0xe -- Background 0xb6
    "00111110", -- 1457 - 0x5b1  :   62 - 0x3e
    "01111111", -- 1458 - 0x5b2  :  127 - 0x7f
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11101111", -- 1461 - 0x5b5  :  239 - 0xef
    "11110111", -- 1462 - 0x5b6  :  247 - 0xf7
    "11111000", -- 1463 - 0x5b7  :  248 - 0xf8
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- Background 0xb7
    "11111111", -- 1465 - 0x5b9  :  255 - 0xff
    "11111111", -- 1466 - 0x5ba  :  255 - 0xff
    "00011111", -- 1467 - 0x5bb  :   31 - 0x1f
    "00011111", -- 1468 - 0x5bc  :   31 - 0x1f
    "01111111", -- 1469 - 0x5bd  :  127 - 0x7f
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "11111110", -- 1471 - 0x5bf  :  254 - 0xfe
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Background 0xb8
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111100", -- 1475 - 0x5c3  :  252 - 0xfc
    "11111000", -- 1476 - 0x5c4  :  248 - 0xf8
    "10000000", -- 1477 - 0x5c5  :  128 - 0x80
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00110000", -- 1480 - 0x5c8  :   48 - 0x30 -- Background 0xb9
    "01111111", -- 1481 - 0x5c9  :  127 - 0x7f
    "01111111", -- 1482 - 0x5ca  :  127 - 0x7f
    "00111111", -- 1483 - 0x5cb  :   63 - 0x3f
    "10000111", -- 1484 - 0x5cc  :  135 - 0x87
    "11110000", -- 1485 - 0x5cd  :  240 - 0xf0
    "11111111", -- 1486 - 0x5ce  :  255 - 0xff
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11100101", -- 1488 - 0x5d0  :  229 - 0xe5 -- Background 0xba
    "11011010", -- 1489 - 0x5d1  :  218 - 0xda
    "11000000", -- 1490 - 0x5d2  :  192 - 0xc0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000110", -- 1496 - 0x5d8  :    6 - 0x6 -- Background 0xbb
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111110", -- 1499 - 0x5db  :  254 - 0xfe
    "11110001", -- 1500 - 0x5dc  :  241 - 0xf1
    "00000111", -- 1501 - 0x5dd  :    7 - 0x7
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0xbc
    "00000001", -- 1505 - 0x5e1  :    1 - 0x1
    "00000010", -- 1506 - 0x5e2  :    2 - 0x2
    "00000111", -- 1507 - 0x5e3  :    7 - 0x7
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00100000", -- 1510 - 0x5e6  :   32 - 0x20
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "01111111", -- 1512 - 0x5e8  :  127 - 0x7f -- Background 0xbd
    "01111111", -- 1513 - 0x5e9  :  127 - 0x7f
    "01111111", -- 1514 - 0x5ea  :  127 - 0x7f
    "11111111", -- 1515 - 0x5eb  :  255 - 0xff
    "11111111", -- 1516 - 0x5ec  :  255 - 0xff
    "11111111", -- 1517 - 0x5ed  :  255 - 0xff
    "11111111", -- 1518 - 0x5ee  :  255 - 0xff
    "11111110", -- 1519 - 0x5ef  :  254 - 0xfe
    "11111100", -- 1520 - 0x5f0  :  252 - 0xfc -- Background 0xbe
    "10111000", -- 1521 - 0x5f1  :  184 - 0xb8
    "01111000", -- 1522 - 0x5f2  :  120 - 0x78
    "01111000", -- 1523 - 0x5f3  :  120 - 0x78
    "10110000", -- 1524 - 0x5f4  :  176 - 0xb0
    "01111000", -- 1525 - 0x5f5  :  120 - 0x78
    "11111100", -- 1526 - 0x5f6  :  252 - 0xfc
    "11111110", -- 1527 - 0x5f7  :  254 - 0xfe
    "11111111", -- 1528 - 0x5f8  :  255 - 0xff -- Background 0xbf
    "11111111", -- 1529 - 0x5f9  :  255 - 0xff
    "11111111", -- 1530 - 0x5fa  :  255 - 0xff
    "11111111", -- 1531 - 0x5fb  :  255 - 0xff
    "11111111", -- 1532 - 0x5fc  :  255 - 0xff
    "10011100", -- 1533 - 0x5fd  :  156 - 0x9c
    "01000010", -- 1534 - 0x5fe  :   66 - 0x42
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00100000", -- 1538 - 0x602  :   32 - 0x20
    "01000000", -- 1539 - 0x603  :   64 - 0x40
    "10001010", -- 1540 - 0x604  :  138 - 0x8a
    "00011110", -- 1541 - 0x605  :   30 - 0x1e
    "01111110", -- 1542 - 0x606  :  126 - 0x7e
    "10111110", -- 1543 - 0x607  :  190 - 0xbe
    "11011111", -- 1544 - 0x608  :  223 - 0xdf -- Background 0xc1
    "11111111", -- 1545 - 0x609  :  255 - 0xff
    "11111110", -- 1546 - 0x60a  :  254 - 0xfe
    "11111100", -- 1547 - 0x60b  :  252 - 0xfc
    "11110000", -- 1548 - 0x60c  :  240 - 0xf0
    "11100000", -- 1549 - 0x60d  :  224 - 0xe0
    "10000000", -- 1550 - 0x60e  :  128 - 0x80
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000100", -- 1554 - 0x612  :    4 - 0x4
    "00000010", -- 1555 - 0x613  :    2 - 0x2
    "01010001", -- 1556 - 0x614  :   81 - 0x51
    "01111000", -- 1557 - 0x615  :  120 - 0x78
    "01111110", -- 1558 - 0x616  :  126 - 0x7e
    "11111101", -- 1559 - 0x617  :  253 - 0xfd
    "11111011", -- 1560 - 0x618  :  251 - 0xfb -- Background 0xc3
    "11111111", -- 1561 - 0x619  :  255 - 0xff
    "01111111", -- 1562 - 0x61a  :  127 - 0x7f
    "00111111", -- 1563 - 0x61b  :   63 - 0x3f
    "00001111", -- 1564 - 0x61c  :   15 - 0xf
    "00000111", -- 1565 - 0x61d  :    7 - 0x7
    "00000001", -- 1566 - 0x61e  :    1 - 0x1
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Background 0xc4
    "10000000", -- 1569 - 0x621  :  128 - 0x80
    "01000000", -- 1570 - 0x622  :   64 - 0x40
    "11100000", -- 1571 - 0x623  :  224 - 0xe0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000100", -- 1574 - 0x626  :    4 - 0x4
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "11111110", -- 1576 - 0x628  :  254 - 0xfe -- Background 0xc5
    "11111110", -- 1577 - 0x629  :  254 - 0xfe
    "11111110", -- 1578 - 0x62a  :  254 - 0xfe
    "11111111", -- 1579 - 0x62b  :  255 - 0xff
    "11111111", -- 1580 - 0x62c  :  255 - 0xff
    "11111111", -- 1581 - 0x62d  :  255 - 0xff
    "11111111", -- 1582 - 0x62e  :  255 - 0xff
    "01111111", -- 1583 - 0x62f  :  127 - 0x7f
    "00111111", -- 1584 - 0x630  :   63 - 0x3f -- Background 0xc6
    "00011101", -- 1585 - 0x631  :   29 - 0x1d
    "00011110", -- 1586 - 0x632  :   30 - 0x1e
    "00011110", -- 1587 - 0x633  :   30 - 0x1e
    "00001101", -- 1588 - 0x634  :   13 - 0xd
    "00011110", -- 1589 - 0x635  :   30 - 0x1e
    "00111111", -- 1590 - 0x636  :   63 - 0x3f
    "01111111", -- 1591 - 0x637  :  127 - 0x7f
    "11111111", -- 1592 - 0x638  :  255 - 0xff -- Background 0xc7
    "11111111", -- 1593 - 0x639  :  255 - 0xff
    "11111111", -- 1594 - 0x63a  :  255 - 0xff
    "11111111", -- 1595 - 0x63b  :  255 - 0xff
    "11111111", -- 1596 - 0x63c  :  255 - 0xff
    "00111001", -- 1597 - 0x63d  :   57 - 0x39
    "01000010", -- 1598 - 0x63e  :   66 - 0x42
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "01101111", -- 1600 - 0x640  :  111 - 0x6f -- Background 0xc8
    "11011011", -- 1601 - 0x641  :  219 - 0xdb
    "00000011", -- 1602 - 0x642  :    3 - 0x3
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "11100000", -- 1615 - 0x64f  :  224 - 0xe0
    "01110000", -- 1616 - 0x650  :  112 - 0x70 -- Background 0xca
    "01111100", -- 1617 - 0x651  :  124 - 0x7c
    "01111110", -- 1618 - 0x652  :  126 - 0x7e
    "11111111", -- 1619 - 0x653  :  255 - 0xff
    "11111111", -- 1620 - 0x654  :  255 - 0xff
    "11110111", -- 1621 - 0x655  :  247 - 0xf7
    "11101111", -- 1622 - 0x656  :  239 - 0xef
    "00011111", -- 1623 - 0x657  :   31 - 0x1f
    "11111111", -- 1624 - 0x658  :  255 - 0xff -- Background 0xcb
    "11111111", -- 1625 - 0x659  :  255 - 0xff
    "11111111", -- 1626 - 0x65a  :  255 - 0xff
    "11111000", -- 1627 - 0x65b  :  248 - 0xf8
    "11111000", -- 1628 - 0x65c  :  248 - 0xf8
    "11111110", -- 1629 - 0x65d  :  254 - 0xfe
    "11111111", -- 1630 - 0x65e  :  255 - 0xff
    "11111111", -- 1631 - 0x65f  :  255 - 0xff
    "11111111", -- 1632 - 0x660  :  255 - 0xff -- Background 0xcc
    "11111111", -- 1633 - 0x661  :  255 - 0xff
    "11111111", -- 1634 - 0x662  :  255 - 0xff
    "00111111", -- 1635 - 0x663  :   63 - 0x3f
    "00011110", -- 1636 - 0x664  :   30 - 0x1e
    "00000001", -- 1637 - 0x665  :    1 - 0x1
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "10000000", -- 1643 - 0x66b  :  128 - 0x80
    "11000000", -- 1644 - 0x66c  :  192 - 0xc0
    "11100000", -- 1645 - 0x66d  :  224 - 0xe0
    "11100000", -- 1646 - 0x66e  :  224 - 0xe0
    "11100000", -- 1647 - 0x66f  :  224 - 0xe0
    "11000000", -- 1648 - 0x670  :  192 - 0xc0 -- Background 0xce
    "10000000", -- 1649 - 0x671  :  128 - 0x80
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "10000000", -- 1654 - 0x676  :  128 - 0x80
    "10000000", -- 1655 - 0x677  :  128 - 0x80
    "10000000", -- 1656 - 0x678  :  128 - 0x80 -- Background 0xcf
    "10000000", -- 1657 - 0x679  :  128 - 0x80
    "11100000", -- 1658 - 0x67a  :  224 - 0xe0
    "11000000", -- 1659 - 0x67b  :  192 - 0xc0
    "00100000", -- 1660 - 0x67c  :   32 - 0x20
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00011111", -- 1664 - 0x680  :   31 - 0x1f -- Background 0xd0
    "00000110", -- 1665 - 0x681  :    6 - 0x6
    "00000110", -- 1666 - 0x682  :    6 - 0x6
    "00000110", -- 1667 - 0x683  :    6 - 0x6
    "00000110", -- 1668 - 0x684  :    6 - 0x6
    "00000110", -- 1669 - 0x685  :    6 - 0x6
    "00000110", -- 1670 - 0x686  :    6 - 0x6
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00111001", -- 1672 - 0x688  :   57 - 0x39 -- Background 0xd1
    "01100101", -- 1673 - 0x689  :  101 - 0x65
    "01100101", -- 1674 - 0x68a  :  101 - 0x65
    "01100101", -- 1675 - 0x68b  :  101 - 0x65
    "01100101", -- 1676 - 0x68c  :  101 - 0x65
    "01100101", -- 1677 - 0x68d  :  101 - 0x65
    "00111001", -- 1678 - 0x68e  :   57 - 0x39
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "11100000", -- 1680 - 0x690  :  224 - 0xe0 -- Background 0xd2
    "10110000", -- 1681 - 0x691  :  176 - 0xb0
    "10110000", -- 1682 - 0x692  :  176 - 0xb0
    "10110110", -- 1683 - 0x693  :  182 - 0xb6
    "11100110", -- 1684 - 0x694  :  230 - 0xe6
    "10000000", -- 1685 - 0x695  :  128 - 0x80
    "10000000", -- 1686 - 0x696  :  128 - 0x80
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00111100", -- 1688 - 0x698  :   60 - 0x3c -- Background 0xd3
    "01000010", -- 1689 - 0x699  :   66 - 0x42
    "10011001", -- 1690 - 0x69a  :  153 - 0x99
    "10100001", -- 1691 - 0x69b  :  161 - 0xa1
    "10100001", -- 1692 - 0x69c  :  161 - 0xa1
    "10011001", -- 1693 - 0x69d  :  153 - 0x99
    "01000010", -- 1694 - 0x69e  :   66 - 0x42
    "00111100", -- 1695 - 0x69f  :   60 - 0x3c
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000011", -- 1699 - 0x6a3  :    3 - 0x3
    "00000110", -- 1700 - 0x6a4  :    6 - 0x6
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000001", -- 1702 - 0x6a6  :    1 - 0x1
    "00000111", -- 1703 - 0x6a7  :    7 - 0x7
    "00001111", -- 1704 - 0x6a8  :   15 - 0xf -- Background 0xd5
    "00011111", -- 1705 - 0x6a9  :   31 - 0x1f
    "00111111", -- 1706 - 0x6aa  :   63 - 0x3f
    "01111111", -- 1707 - 0x6ab  :  127 - 0x7f
    "01111111", -- 1708 - 0x6ac  :  127 - 0x7f
    "01111111", -- 1709 - 0x6ad  :  127 - 0x7f
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "01111111", -- 1711 - 0x6af  :  127 - 0x7f
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "10000000", -- 1715 - 0x6b3  :  128 - 0x80
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "10100000", -- 1719 - 0x6b7  :  160 - 0xa0
    "11100000", -- 1720 - 0x6b8  :  224 - 0xe0 -- Background 0xd7
    "11110000", -- 1721 - 0x6b9  :  240 - 0xf0
    "11100000", -- 1722 - 0x6ba  :  224 - 0xe0
    "11011101", -- 1723 - 0x6bb  :  221 - 0xdd
    "11111010", -- 1724 - 0x6bc  :  250 - 0xfa
    "11101011", -- 1725 - 0x6bd  :  235 - 0xeb
    "10000000", -- 1726 - 0x6be  :  128 - 0x80
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000011", -- 1731 - 0x6c3  :    3 - 0x3
    "00000110", -- 1732 - 0x6c4  :    6 - 0x6
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000001", -- 1734 - 0x6c6  :    1 - 0x1
    "00000001", -- 1735 - 0x6c7  :    1 - 0x1
    "00001011", -- 1736 - 0x6c8  :   11 - 0xb -- Background 0xd9
    "00000111", -- 1737 - 0x6c9  :    7 - 0x7
    "00000011", -- 1738 - 0x6ca  :    3 - 0x3
    "01011101", -- 1739 - 0x6cb  :   93 - 0x5d
    "10101111", -- 1740 - 0x6cc  :  175 - 0xaf
    "01010011", -- 1741 - 0x6cd  :   83 - 0x53
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "10000000", -- 1747 - 0x6d3  :  128 - 0x80
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "01100000", -- 1750 - 0x6d6  :   96 - 0x60
    "11110000", -- 1751 - 0x6d7  :  240 - 0xf0
    "11111000", -- 1752 - 0x6d8  :  248 - 0xf8 -- Background 0xdb
    "11111100", -- 1753 - 0x6d9  :  252 - 0xfc
    "11111100", -- 1754 - 0x6da  :  252 - 0xfc
    "11111110", -- 1755 - 0x6db  :  254 - 0xfe
    "11111110", -- 1756 - 0x6dc  :  254 - 0xfe
    "11111111", -- 1757 - 0x6dd  :  255 - 0xff
    "11111111", -- 1758 - 0x6de  :  255 - 0xff
    "01111110", -- 1759 - 0x6df  :  126 - 0x7e
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00100001", -- 1766 - 0x6e6  :   33 - 0x21
    "00111111", -- 1767 - 0x6e7  :   63 - 0x3f
    "00111111", -- 1768 - 0x6e8  :   63 - 0x3f -- Background 0xdd
    "00011111", -- 1769 - 0x6e9  :   31 - 0x1f
    "00011111", -- 1770 - 0x6ea  :   31 - 0x1f
    "00001111", -- 1771 - 0x6eb  :   15 - 0xf
    "00000111", -- 1772 - 0x6ec  :    7 - 0x7
    "00000011", -- 1773 - 0x6ed  :    3 - 0x3
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00111110", -- 1776 - 0x6f0  :   62 - 0x3e -- Background 0xde
    "00011110", -- 1777 - 0x6f1  :   30 - 0x1e
    "00011110", -- 1778 - 0x6f2  :   30 - 0x1e
    "00001110", -- 1779 - 0x6f3  :   14 - 0xe
    "00001111", -- 1780 - 0x6f4  :   15 - 0xf
    "00011111", -- 1781 - 0x6f5  :   31 - 0x1f
    "10011111", -- 1782 - 0x6f6  :  159 - 0x9f
    "10011111", -- 1783 - 0x6f7  :  159 - 0x9f
    "11011111", -- 1784 - 0x6f8  :  223 - 0xdf -- Background 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11111111", -- 1788 - 0x6fc  :  255 - 0xff
    "11011111", -- 1789 - 0x6fd  :  223 - 0xdf
    "11100111", -- 1790 - 0x6fe  :  231 - 0xe7
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00100000", -- 1792 - 0x700  :   32 - 0x20 -- Background 0xe0
    "00001111", -- 1793 - 0x701  :   15 - 0xf
    "00110000", -- 1794 - 0x702  :   48 - 0x30
    "01000000", -- 1795 - 0x703  :   64 - 0x40
    "10011000", -- 1796 - 0x704  :  152 - 0x98
    "00111110", -- 1797 - 0x705  :   62 - 0x3e
    "00011111", -- 1798 - 0x706  :   31 - 0x1f
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "10000001", -- 1800 - 0x708  :  129 - 0x81 -- Background 0xe1
    "00110110", -- 1801 - 0x709  :   54 - 0x36
    "00101110", -- 1802 - 0x70a  :   46 - 0x2e
    "10101111", -- 1803 - 0x70b  :  175 - 0xaf
    "10101110", -- 1804 - 0x70c  :  174 - 0xae
    "11010001", -- 1805 - 0x70d  :  209 - 0xd1
    "11101111", -- 1806 - 0x70e  :  239 - 0xef
    "10000111", -- 1807 - 0x70f  :  135 - 0x87
    "00000010", -- 1808 - 0x710  :    2 - 0x2 -- Background 0xe2
    "11111000", -- 1809 - 0x711  :  248 - 0xf8
    "00000110", -- 1810 - 0x712  :    6 - 0x6
    "00000001", -- 1811 - 0x713  :    1 - 0x1
    "00001100", -- 1812 - 0x714  :   12 - 0xc
    "00111110", -- 1813 - 0x715  :   62 - 0x3e
    "11111100", -- 1814 - 0x716  :  252 - 0xfc
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "11000000", -- 1816 - 0x718  :  192 - 0xc0 -- Background 0xe3
    "00110110", -- 1817 - 0x719  :   54 - 0x36
    "00111110", -- 1818 - 0x71a  :   62 - 0x3e
    "01111010", -- 1819 - 0x71b  :  122 - 0x7a
    "10110110", -- 1820 - 0x71c  :  182 - 0xb6
    "11001101", -- 1821 - 0x71d  :  205 - 0xcd
    "11111011", -- 1822 - 0x71e  :  251 - 0xfb
    "11110000", -- 1823 - 0x71f  :  240 - 0xf0
    "00111110", -- 1824 - 0x720  :   62 - 0x3e -- Background 0xe4
    "00111100", -- 1825 - 0x721  :   60 - 0x3c
    "00111100", -- 1826 - 0x722  :   60 - 0x3c
    "00111000", -- 1827 - 0x723  :   56 - 0x38
    "11111000", -- 1828 - 0x724  :  248 - 0xf8
    "01111100", -- 1829 - 0x725  :  124 - 0x7c
    "01111110", -- 1830 - 0x726  :  126 - 0x7e
    "01111000", -- 1831 - 0x727  :  120 - 0x78
    "11111000", -- 1832 - 0x728  :  248 - 0xf8 -- Background 0xe5
    "01111111", -- 1833 - 0x729  :  127 - 0x7f
    "01111111", -- 1834 - 0x72a  :  127 - 0x7f
    "11111110", -- 1835 - 0x72b  :  254 - 0xfe
    "11111111", -- 1836 - 0x72c  :  255 - 0xff
    "11111111", -- 1837 - 0x72d  :  255 - 0xff
    "11110011", -- 1838 - 0x72e  :  243 - 0xf3
    "10000001", -- 1839 - 0x72f  :  129 - 0x81
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00010000", -- 1843 - 0x733  :   16 - 0x10
    "01000000", -- 1844 - 0x734  :   64 - 0x40
    "00100000", -- 1845 - 0x735  :   32 - 0x20
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000110", -- 1848 - 0x738  :    6 - 0x6 -- Background 0xe7
    "00001110", -- 1849 - 0x739  :   14 - 0xe
    "01111110", -- 1850 - 0x73a  :  126 - 0x7e
    "11111110", -- 1851 - 0x73b  :  254 - 0xfe
    "11111110", -- 1852 - 0x73c  :  254 - 0xfe
    "11111100", -- 1853 - 0x73d  :  252 - 0xfc
    "11111000", -- 1854 - 0x73e  :  248 - 0xf8
    "11110000", -- 1855 - 0x73f  :  240 - 0xf0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000001", -- 1863 - 0x747  :    1 - 0x1
    "00000010", -- 1864 - 0x748  :    2 - 0x2 -- Background 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00001000", -- 1866 - 0x74a  :    8 - 0x8
    "00000001", -- 1867 - 0x74b  :    1 - 0x1
    "00010011", -- 1868 - 0x74c  :   19 - 0x13
    "00000001", -- 1869 - 0x74d  :    1 - 0x1
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Background 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Background 0xeb
    "01000011", -- 1881 - 0x759  :   67 - 0x43
    "01111111", -- 1882 - 0x75a  :  127 - 0x7f
    "01111111", -- 1883 - 0x75b  :  127 - 0x7f
    "01111111", -- 1884 - 0x75c  :  127 - 0x7f
    "00111111", -- 1885 - 0x75d  :   63 - 0x3f
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "11000000", -- 1894 - 0x766  :  192 - 0xc0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00010000", -- 1896 - 0x768  :   16 - 0x10 -- Background 0xed
    "00111000", -- 1897 - 0x769  :   56 - 0x38
    "10111111", -- 1898 - 0x76a  :  191 - 0xbf
    "11111111", -- 1899 - 0x76b  :  255 - 0xff
    "11111111", -- 1900 - 0x76c  :  255 - 0xff
    "11111111", -- 1901 - 0x76d  :  255 - 0xff
    "11111111", -- 1902 - 0x76e  :  255 - 0xff
    "11111111", -- 1903 - 0x76f  :  255 - 0xff
    "01111110", -- 1904 - 0x770  :  126 - 0x7e -- Background 0xee
    "00011110", -- 1905 - 0x771  :   30 - 0x1e
    "00011110", -- 1906 - 0x772  :   30 - 0x1e
    "00001110", -- 1907 - 0x773  :   14 - 0xe
    "00001111", -- 1908 - 0x774  :   15 - 0xf
    "00011110", -- 1909 - 0x775  :   30 - 0x1e
    "00011110", -- 1910 - 0x776  :   30 - 0x1e
    "00111110", -- 1911 - 0x777  :   62 - 0x3e
    "01111111", -- 1912 - 0x778  :  127 - 0x7f -- Background 0xef
    "01111111", -- 1913 - 0x779  :  127 - 0x7f
    "10111111", -- 1914 - 0x77a  :  191 - 0xbf
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111111", -- 1916 - 0x77c  :  255 - 0xff
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11100111", -- 1918 - 0x77e  :  231 - 0xe7
    "11000000", -- 1919 - 0x77f  :  192 - 0xc0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00010000", -- 1922 - 0x782  :   16 - 0x10
    "11111101", -- 1923 - 0x783  :  253 - 0xfd
    "11111010", -- 1924 - 0x784  :  250 - 0xfa
    "11101011", -- 1925 - 0x785  :  235 - 0xeb
    "10000000", -- 1926 - 0x786  :  128 - 0x80
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00100000", -- 1928 - 0x788  :   32 - 0x20 -- Background 0xf1
    "00011111", -- 1929 - 0x789  :   31 - 0x1f
    "01100000", -- 1930 - 0x78a  :   96 - 0x60
    "10001110", -- 1931 - 0x78b  :  142 - 0x8e
    "00111111", -- 1932 - 0x78c  :   63 - 0x3f
    "01111111", -- 1933 - 0x78d  :  127 - 0x7f
    "01111111", -- 1934 - 0x78e  :  127 - 0x7f
    "01111100", -- 1935 - 0x78f  :  124 - 0x7c
    "00111001", -- 1936 - 0x790  :   57 - 0x39 -- Background 0xf2
    "00110110", -- 1937 - 0x791  :   54 - 0x36
    "00101110", -- 1938 - 0x792  :   46 - 0x2e
    "10101111", -- 1939 - 0x793  :  175 - 0xaf
    "10101110", -- 1940 - 0x794  :  174 - 0xae
    "11010001", -- 1941 - 0x795  :  209 - 0xd1
    "11101111", -- 1942 - 0x796  :  239 - 0xef
    "10000111", -- 1943 - 0x797  :  135 - 0x87
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000100", -- 1946 - 0x79a  :    4 - 0x4
    "01011111", -- 1947 - 0x79b  :   95 - 0x5f
    "10101111", -- 1948 - 0x79c  :  175 - 0xaf
    "01010011", -- 1949 - 0x79d  :   83 - 0x53
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000010", -- 1952 - 0x7a0  :    2 - 0x2 -- Background 0xf4
    "11111100", -- 1953 - 0x7a1  :  252 - 0xfc
    "00000011", -- 1954 - 0x7a2  :    3 - 0x3
    "00111000", -- 1955 - 0x7a3  :   56 - 0x38
    "11111110", -- 1956 - 0x7a4  :  254 - 0xfe
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "00011110", -- 1959 - 0x7a7  :   30 - 0x1e
    "11000000", -- 1960 - 0x7a8  :  192 - 0xc0 -- Background 0xf5
    "00110110", -- 1961 - 0x7a9  :   54 - 0x36
    "00111110", -- 1962 - 0x7aa  :   62 - 0x3e
    "01111010", -- 1963 - 0x7ab  :  122 - 0x7a
    "10110110", -- 1964 - 0x7ac  :  182 - 0xb6
    "11001101", -- 1965 - 0x7ad  :  205 - 0xcd
    "11111011", -- 1966 - 0x7ae  :  251 - 0xfb
    "11110000", -- 1967 - 0x7af  :  240 - 0xf0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00001110", -- 1973 - 0x7b5  :   14 - 0xe
    "00001000", -- 1974 - 0x7b6  :    8 - 0x8
    "00001000", -- 1975 - 0x7b7  :    8 - 0x8
    "00011111", -- 1976 - 0x7b8  :   31 - 0x1f -- Background 0xf7
    "00111111", -- 1977 - 0x7b9  :   63 - 0x3f
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "01111111", -- 1983 - 0x7bf  :  127 - 0x7f
    "00111111", -- 1984 - 0x7c0  :   63 - 0x3f -- Background 0xf8
    "00111110", -- 1985 - 0x7c1  :   62 - 0x3e
    "00111100", -- 1986 - 0x7c2  :   60 - 0x3c
    "10111000", -- 1987 - 0x7c3  :  184 - 0xb8
    "01111000", -- 1988 - 0x7c4  :  120 - 0x78
    "01111000", -- 1989 - 0x7c5  :  120 - 0x78
    "01111110", -- 1990 - 0x7c6  :  126 - 0x7e
    "01111110", -- 1991 - 0x7c7  :  126 - 0x7e
    "11111101", -- 1992 - 0x7c8  :  253 - 0xfd -- Background 0xf9
    "01111001", -- 1993 - 0x7c9  :  121 - 0x79
    "01111011", -- 1994 - 0x7ca  :  123 - 0x7b
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11110011", -- 1998 - 0x7ce  :  243 - 0xf3
    "10000000", -- 1999 - 0x7cf  :  128 - 0x80
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00010000", -- 2008 - 0x7d8  :   16 - 0x10 -- Background 0xfb
    "10000100", -- 2009 - 0x7d9  :  132 - 0x84
    "11100000", -- 2010 - 0x7da  :  224 - 0xe0
    "11000000", -- 2011 - 0x7db  :  192 - 0xc0
    "10000000", -- 2012 - 0x7dc  :  128 - 0x80
    "10000000", -- 2013 - 0x7dd  :  128 - 0x80
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Background 0xfc
    "01001000", -- 2017 - 0x7e1  :   72 - 0x48
    "00100000", -- 2018 - 0x7e2  :   32 - 0x20
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000100", -- 2021 - 0x7e5  :    4 - 0x4
    "00001110", -- 2022 - 0x7e6  :   14 - 0xe
    "11111110", -- 2023 - 0x7e7  :  254 - 0xfe
    "11111110", -- 2024 - 0x7e8  :  254 - 0xfe -- Background 0xfd
    "11111100", -- 2025 - 0x7e9  :  252 - 0xfc
    "11111100", -- 2026 - 0x7ea  :  252 - 0xfc
    "11111000", -- 2027 - 0x7eb  :  248 - 0xf8
    "11110000", -- 2028 - 0x7ec  :  240 - 0xf0
    "11100000", -- 2029 - 0x7ed  :  224 - 0xe0
    "10000000", -- 2030 - 0x7ee  :  128 - 0x80
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00001111", -- 2032 - 0x7f0  :   15 - 0xf -- Background 0xfe
    "00000110", -- 2033 - 0x7f1  :    6 - 0x6
    "00000110", -- 2034 - 0x7f2  :    6 - 0x6
    "00000110", -- 2035 - 0x7f3  :    6 - 0x6
    "00000110", -- 2036 - 0x7f4  :    6 - 0x6
    "00000110", -- 2037 - 0x7f5  :    6 - 0x6
    "00001111", -- 2038 - 0x7f6  :   15 - 0xf
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "11110000", -- 2040 - 0x7f8  :  240 - 0xf0 -- Background 0xff
    "01100000", -- 2041 - 0x7f9  :   96 - 0x60
    "01100000", -- 2042 - 0x7fa  :   96 - 0x60
    "01100110", -- 2043 - 0x7fb  :  102 - 0x66
    "01100110", -- 2044 - 0x7fc  :  102 - 0x66
    "01100000", -- 2045 - 0x7fd  :   96 - 0x60
    "11110000", -- 2046 - 0x7fe  :  240 - 0xf0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
