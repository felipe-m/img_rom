---   Background Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG_BG is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG_BG;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG_BG is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table both color planes
    "00111000", --    0 -  0x0  :   56 - 0x38 -- Background 0x0
    "01001100", --    1 -  0x1  :   76 - 0x4c
    "11000110", --    2 -  0x2  :  198 - 0xc6
    "11000110", --    3 -  0x3  :  198 - 0xc6
    "11000110", --    4 -  0x4  :  198 - 0xc6
    "01100100", --    5 -  0x5  :  100 - 0x64
    "00111000", --    6 -  0x6  :   56 - 0x38
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00011000", --   16 - 0x10  :   24 - 0x18 -- Background 0x1
    "00111000", --   17 - 0x11  :   56 - 0x38
    "00011000", --   18 - 0x12  :   24 - 0x18
    "00011000", --   19 - 0x13  :   24 - 0x18
    "00011000", --   20 - 0x14  :   24 - 0x18
    "00011000", --   21 - 0x15  :   24 - 0x18
    "01111110", --   22 - 0x16  :  126 - 0x7e
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "01111100", --   32 - 0x20  :  124 - 0x7c -- Background 0x2
    "11000110", --   33 - 0x21  :  198 - 0xc6
    "00001110", --   34 - 0x22  :   14 - 0xe
    "00111100", --   35 - 0x23  :   60 - 0x3c
    "01111000", --   36 - 0x24  :  120 - 0x78
    "11100000", --   37 - 0x25  :  224 - 0xe0
    "11111110", --   38 - 0x26  :  254 - 0xfe
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "01111110", --   48 - 0x30  :  126 - 0x7e -- Background 0x3
    "00001100", --   49 - 0x31  :   12 - 0xc
    "00011000", --   50 - 0x32  :   24 - 0x18
    "00111100", --   51 - 0x33  :   60 - 0x3c
    "00000110", --   52 - 0x34  :    6 - 0x6
    "11000110", --   53 - 0x35  :  198 - 0xc6
    "01111100", --   54 - 0x36  :  124 - 0x7c
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- plane 1
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00011100", --   64 - 0x40  :   28 - 0x1c -- Background 0x4
    "00111100", --   65 - 0x41  :   60 - 0x3c
    "01101100", --   66 - 0x42  :  108 - 0x6c
    "11001100", --   67 - 0x43  :  204 - 0xcc
    "11111110", --   68 - 0x44  :  254 - 0xfe
    "00001100", --   69 - 0x45  :   12 - 0xc
    "00001100", --   70 - 0x46  :   12 - 0xc
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- plane 1
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "11111100", --   80 - 0x50  :  252 - 0xfc -- Background 0x5
    "11000000", --   81 - 0x51  :  192 - 0xc0
    "11111100", --   82 - 0x52  :  252 - 0xfc
    "00000110", --   83 - 0x53  :    6 - 0x6
    "00000110", --   84 - 0x54  :    6 - 0x6
    "11000110", --   85 - 0x55  :  198 - 0xc6
    "01111100", --   86 - 0x56  :  124 - 0x7c
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- plane 1
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00111100", --   96 - 0x60  :   60 - 0x3c -- Background 0x6
    "01100000", --   97 - 0x61  :   96 - 0x60
    "11000000", --   98 - 0x62  :  192 - 0xc0
    "11111100", --   99 - 0x63  :  252 - 0xfc
    "11000110", --  100 - 0x64  :  198 - 0xc6
    "11000110", --  101 - 0x65  :  198 - 0xc6
    "01111100", --  102 - 0x66  :  124 - 0x7c
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- plane 1
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11111110", --  112 - 0x70  :  254 - 0xfe -- Background 0x7
    "11000110", --  113 - 0x71  :  198 - 0xc6
    "00001100", --  114 - 0x72  :   12 - 0xc
    "00011000", --  115 - 0x73  :   24 - 0x18
    "00110000", --  116 - 0x74  :   48 - 0x30
    "00110000", --  117 - 0x75  :   48 - 0x30
    "00110000", --  118 - 0x76  :   48 - 0x30
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- plane 1
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "01111000", --  128 - 0x80  :  120 - 0x78 -- Background 0x8
    "11000100", --  129 - 0x81  :  196 - 0xc4
    "11100100", --  130 - 0x82  :  228 - 0xe4
    "01111000", --  131 - 0x83  :  120 - 0x78
    "10000110", --  132 - 0x84  :  134 - 0x86
    "10000110", --  133 - 0x85  :  134 - 0x86
    "01111100", --  134 - 0x86  :  124 - 0x7c
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- plane 1
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01111100", --  144 - 0x90  :  124 - 0x7c -- Background 0x9
    "11000110", --  145 - 0x91  :  198 - 0xc6
    "11000110", --  146 - 0x92  :  198 - 0xc6
    "01111110", --  147 - 0x93  :  126 - 0x7e
    "00000110", --  148 - 0x94  :    6 - 0x6
    "00001100", --  149 - 0x95  :   12 - 0xc
    "01111000", --  150 - 0x96  :  120 - 0x78
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- plane 1
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00111000", --  160 - 0xa0  :   56 - 0x38 -- Background 0xa
    "01101100", --  161 - 0xa1  :  108 - 0x6c
    "11000110", --  162 - 0xa2  :  198 - 0xc6
    "11000110", --  163 - 0xa3  :  198 - 0xc6
    "11111110", --  164 - 0xa4  :  254 - 0xfe
    "11000110", --  165 - 0xa5  :  198 - 0xc6
    "11000110", --  166 - 0xa6  :  198 - 0xc6
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- plane 1
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11111100", --  176 - 0xb0  :  252 - 0xfc -- Background 0xb
    "11000110", --  177 - 0xb1  :  198 - 0xc6
    "11000110", --  178 - 0xb2  :  198 - 0xc6
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11000110", --  180 - 0xb4  :  198 - 0xc6
    "11000110", --  181 - 0xb5  :  198 - 0xc6
    "11111100", --  182 - 0xb6  :  252 - 0xfc
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- plane 1
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00111100", --  192 - 0xc0  :   60 - 0x3c -- Background 0xc
    "01100110", --  193 - 0xc1  :  102 - 0x66
    "11000000", --  194 - 0xc2  :  192 - 0xc0
    "11000000", --  195 - 0xc3  :  192 - 0xc0
    "11000000", --  196 - 0xc4  :  192 - 0xc0
    "01100110", --  197 - 0xc5  :  102 - 0x66
    "00111100", --  198 - 0xc6  :   60 - 0x3c
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- plane 1
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "11111000", --  208 - 0xd0  :  248 - 0xf8 -- Background 0xd
    "11001100", --  209 - 0xd1  :  204 - 0xcc
    "11000110", --  210 - 0xd2  :  198 - 0xc6
    "11000110", --  211 - 0xd3  :  198 - 0xc6
    "11000110", --  212 - 0xd4  :  198 - 0xc6
    "11001100", --  213 - 0xd5  :  204 - 0xcc
    "11111000", --  214 - 0xd6  :  248 - 0xf8
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- plane 1
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "11111110", --  224 - 0xe0  :  254 - 0xfe -- Background 0xe
    "11000000", --  225 - 0xe1  :  192 - 0xc0
    "11000000", --  226 - 0xe2  :  192 - 0xc0
    "11111100", --  227 - 0xe3  :  252 - 0xfc
    "11000000", --  228 - 0xe4  :  192 - 0xc0
    "11000000", --  229 - 0xe5  :  192 - 0xc0
    "11111110", --  230 - 0xe6  :  254 - 0xfe
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- plane 1
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11111110", --  240 - 0xf0  :  254 - 0xfe -- Background 0xf
    "11000000", --  241 - 0xf1  :  192 - 0xc0
    "11000000", --  242 - 0xf2  :  192 - 0xc0
    "11111100", --  243 - 0xf3  :  252 - 0xfc
    "11000000", --  244 - 0xf4  :  192 - 0xc0
    "11000000", --  245 - 0xf5  :  192 - 0xc0
    "11000000", --  246 - 0xf6  :  192 - 0xc0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- plane 1
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00111110", --  256 - 0x100  :   62 - 0x3e -- Background 0x10
    "01100000", --  257 - 0x101  :   96 - 0x60
    "11000000", --  258 - 0x102  :  192 - 0xc0
    "11011110", --  259 - 0x103  :  222 - 0xde
    "11000110", --  260 - 0x104  :  198 - 0xc6
    "01100110", --  261 - 0x105  :  102 - 0x66
    "01111110", --  262 - 0x106  :  126 - 0x7e
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- plane 1
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "11000110", --  272 - 0x110  :  198 - 0xc6 -- Background 0x11
    "11000110", --  273 - 0x111  :  198 - 0xc6
    "11000110", --  274 - 0x112  :  198 - 0xc6
    "11111110", --  275 - 0x113  :  254 - 0xfe
    "11000110", --  276 - 0x114  :  198 - 0xc6
    "11000110", --  277 - 0x115  :  198 - 0xc6
    "11000110", --  278 - 0x116  :  198 - 0xc6
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- plane 1
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "01111110", --  288 - 0x120  :  126 - 0x7e -- Background 0x12
    "00011000", --  289 - 0x121  :   24 - 0x18
    "00011000", --  290 - 0x122  :   24 - 0x18
    "00011000", --  291 - 0x123  :   24 - 0x18
    "00011000", --  292 - 0x124  :   24 - 0x18
    "00011000", --  293 - 0x125  :   24 - 0x18
    "01111110", --  294 - 0x126  :  126 - 0x7e
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- plane 1
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00011110", --  304 - 0x130  :   30 - 0x1e -- Background 0x13
    "00000110", --  305 - 0x131  :    6 - 0x6
    "00000110", --  306 - 0x132  :    6 - 0x6
    "00000110", --  307 - 0x133  :    6 - 0x6
    "11000110", --  308 - 0x134  :  198 - 0xc6
    "11000110", --  309 - 0x135  :  198 - 0xc6
    "01111100", --  310 - 0x136  :  124 - 0x7c
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- plane 1
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "11000110", --  320 - 0x140  :  198 - 0xc6 -- Background 0x14
    "11001100", --  321 - 0x141  :  204 - 0xcc
    "11011000", --  322 - 0x142  :  216 - 0xd8
    "11110000", --  323 - 0x143  :  240 - 0xf0
    "11111000", --  324 - 0x144  :  248 - 0xf8
    "11011100", --  325 - 0x145  :  220 - 0xdc
    "11001110", --  326 - 0x146  :  206 - 0xce
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- plane 1
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "01100000", --  336 - 0x150  :   96 - 0x60 -- Background 0x15
    "01100000", --  337 - 0x151  :   96 - 0x60
    "01100000", --  338 - 0x152  :   96 - 0x60
    "01100000", --  339 - 0x153  :   96 - 0x60
    "01100000", --  340 - 0x154  :   96 - 0x60
    "01100000", --  341 - 0x155  :   96 - 0x60
    "01111110", --  342 - 0x156  :  126 - 0x7e
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0 -- plane 1
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "11000110", --  352 - 0x160  :  198 - 0xc6 -- Background 0x16
    "11101110", --  353 - 0x161  :  238 - 0xee
    "11111110", --  354 - 0x162  :  254 - 0xfe
    "11111110", --  355 - 0x163  :  254 - 0xfe
    "11010110", --  356 - 0x164  :  214 - 0xd6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "11000110", --  358 - 0x166  :  198 - 0xc6
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- plane 1
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "11000110", --  368 - 0x170  :  198 - 0xc6 -- Background 0x17
    "11100110", --  369 - 0x171  :  230 - 0xe6
    "11110110", --  370 - 0x172  :  246 - 0xf6
    "11111110", --  371 - 0x173  :  254 - 0xfe
    "11011110", --  372 - 0x174  :  222 - 0xde
    "11001110", --  373 - 0x175  :  206 - 0xce
    "11000110", --  374 - 0x176  :  198 - 0xc6
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- plane 1
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "01111100", --  384 - 0x180  :  124 - 0x7c -- Background 0x18
    "11000110", --  385 - 0x181  :  198 - 0xc6
    "11000110", --  386 - 0x182  :  198 - 0xc6
    "11000110", --  387 - 0x183  :  198 - 0xc6
    "11000110", --  388 - 0x184  :  198 - 0xc6
    "11000110", --  389 - 0x185  :  198 - 0xc6
    "01111100", --  390 - 0x186  :  124 - 0x7c
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- plane 1
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "11111100", --  400 - 0x190  :  252 - 0xfc -- Background 0x19
    "11000110", --  401 - 0x191  :  198 - 0xc6
    "11000110", --  402 - 0x192  :  198 - 0xc6
    "11000110", --  403 - 0x193  :  198 - 0xc6
    "11111100", --  404 - 0x194  :  252 - 0xfc
    "11000000", --  405 - 0x195  :  192 - 0xc0
    "11000000", --  406 - 0x196  :  192 - 0xc0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- plane 1
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "01111100", --  416 - 0x1a0  :  124 - 0x7c -- Background 0x1a
    "11000110", --  417 - 0x1a1  :  198 - 0xc6
    "11000110", --  418 - 0x1a2  :  198 - 0xc6
    "11000110", --  419 - 0x1a3  :  198 - 0xc6
    "11011110", --  420 - 0x1a4  :  222 - 0xde
    "11001100", --  421 - 0x1a5  :  204 - 0xcc
    "01111010", --  422 - 0x1a6  :  122 - 0x7a
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- plane 1
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "11111100", --  432 - 0x1b0  :  252 - 0xfc -- Background 0x1b
    "11000110", --  433 - 0x1b1  :  198 - 0xc6
    "11000110", --  434 - 0x1b2  :  198 - 0xc6
    "11001110", --  435 - 0x1b3  :  206 - 0xce
    "11111000", --  436 - 0x1b4  :  248 - 0xf8
    "11011100", --  437 - 0x1b5  :  220 - 0xdc
    "11001110", --  438 - 0x1b6  :  206 - 0xce
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- plane 1
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "01111000", --  448 - 0x1c0  :  120 - 0x78 -- Background 0x1c
    "11001100", --  449 - 0x1c1  :  204 - 0xcc
    "11000000", --  450 - 0x1c2  :  192 - 0xc0
    "01111100", --  451 - 0x1c3  :  124 - 0x7c
    "00000110", --  452 - 0x1c4  :    6 - 0x6
    "11000110", --  453 - 0x1c5  :  198 - 0xc6
    "01111100", --  454 - 0x1c6  :  124 - 0x7c
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- plane 1
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "01111110", --  464 - 0x1d0  :  126 - 0x7e -- Background 0x1d
    "00011000", --  465 - 0x1d1  :   24 - 0x18
    "00011000", --  466 - 0x1d2  :   24 - 0x18
    "00011000", --  467 - 0x1d3  :   24 - 0x18
    "00011000", --  468 - 0x1d4  :   24 - 0x18
    "00011000", --  469 - 0x1d5  :   24 - 0x18
    "00011000", --  470 - 0x1d6  :   24 - 0x18
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- plane 1
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "11000110", --  480 - 0x1e0  :  198 - 0xc6 -- Background 0x1e
    "11000110", --  481 - 0x1e1  :  198 - 0xc6
    "11000110", --  482 - 0x1e2  :  198 - 0xc6
    "11000110", --  483 - 0x1e3  :  198 - 0xc6
    "11000110", --  484 - 0x1e4  :  198 - 0xc6
    "11000110", --  485 - 0x1e5  :  198 - 0xc6
    "01111100", --  486 - 0x1e6  :  124 - 0x7c
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- plane 1
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "11000110", --  496 - 0x1f0  :  198 - 0xc6 -- Background 0x1f
    "11000110", --  497 - 0x1f1  :  198 - 0xc6
    "11000110", --  498 - 0x1f2  :  198 - 0xc6
    "11101110", --  499 - 0x1f3  :  238 - 0xee
    "01111100", --  500 - 0x1f4  :  124 - 0x7c
    "00111000", --  501 - 0x1f5  :   56 - 0x38
    "00010000", --  502 - 0x1f6  :   16 - 0x10
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- plane 1
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "11000110", --  512 - 0x200  :  198 - 0xc6 -- Background 0x20
    "11000110", --  513 - 0x201  :  198 - 0xc6
    "11010110", --  514 - 0x202  :  214 - 0xd6
    "11111110", --  515 - 0x203  :  254 - 0xfe
    "11111110", --  516 - 0x204  :  254 - 0xfe
    "11101110", --  517 - 0x205  :  238 - 0xee
    "11000110", --  518 - 0x206  :  198 - 0xc6
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "11000110", --  528 - 0x210  :  198 - 0xc6 -- Background 0x21
    "11101110", --  529 - 0x211  :  238 - 0xee
    "01111100", --  530 - 0x212  :  124 - 0x7c
    "00111000", --  531 - 0x213  :   56 - 0x38
    "01111100", --  532 - 0x214  :  124 - 0x7c
    "11101110", --  533 - 0x215  :  238 - 0xee
    "11000110", --  534 - 0x216  :  198 - 0xc6
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- plane 1
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01100110", --  544 - 0x220  :  102 - 0x66 -- Background 0x22
    "01100110", --  545 - 0x221  :  102 - 0x66
    "01100110", --  546 - 0x222  :  102 - 0x66
    "00111100", --  547 - 0x223  :   60 - 0x3c
    "00011000", --  548 - 0x224  :   24 - 0x18
    "00011000", --  549 - 0x225  :   24 - 0x18
    "00011000", --  550 - 0x226  :   24 - 0x18
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- plane 1
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "11111110", --  560 - 0x230  :  254 - 0xfe -- Background 0x23
    "00001110", --  561 - 0x231  :   14 - 0xe
    "00011100", --  562 - 0x232  :   28 - 0x1c
    "00111000", --  563 - 0x233  :   56 - 0x38
    "01110000", --  564 - 0x234  :  112 - 0x70
    "11100000", --  565 - 0x235  :  224 - 0xe0
    "11111110", --  566 - 0x236  :  254 - 0xfe
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- plane 1
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x24
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- plane 1
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Background 0x25
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000110", --  594 - 0x252  :    6 - 0x6
    "00001110", --  595 - 0x253  :   14 - 0xe
    "00001000", --  596 - 0x254  :    8 - 0x8
    "00001000", --  597 - 0x255  :    8 - 0x8
    "00001000", --  598 - 0x256  :    8 - 0x8
    "00001000", --  599 - 0x257  :    8 - 0x8
    "00000000", --  600 - 0x258  :    0 - 0x0 -- plane 1
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x26
    "01111000", --  609 - 0x261  :  120 - 0x78
    "01100101", --  610 - 0x262  :  101 - 0x65
    "01111001", --  611 - 0x263  :  121 - 0x79
    "01100101", --  612 - 0x264  :  101 - 0x65
    "01100101", --  613 - 0x265  :  101 - 0x65
    "01111000", --  614 - 0x266  :  120 - 0x78
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- plane 1
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x27
    "11100100", --  625 - 0x271  :  228 - 0xe4
    "10010110", --  626 - 0x272  :  150 - 0x96
    "10010110", --  627 - 0x273  :  150 - 0x96
    "10010111", --  628 - 0x274  :  151 - 0x97
    "10010110", --  629 - 0x275  :  150 - 0x96
    "11100110", --  630 - 0x276  :  230 - 0xe6
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- plane 1
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x28
    "01011001", --  641 - 0x281  :   89 - 0x59
    "01011001", --  642 - 0x282  :   89 - 0x59
    "01011001", --  643 - 0x283  :   89 - 0x59
    "01011001", --  644 - 0x284  :   89 - 0x59
    "11011001", --  645 - 0x285  :  217 - 0xd9
    "01001110", --  646 - 0x286  :   78 - 0x4e
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x29
    "00111100", --  657 - 0x291  :   60 - 0x3c
    "01110000", --  658 - 0x292  :  112 - 0x70
    "01110000", --  659 - 0x293  :  112 - 0x70
    "00111100", --  660 - 0x294  :   60 - 0x3c
    "00001100", --  661 - 0x295  :   12 - 0xc
    "01111000", --  662 - 0x296  :  120 - 0x78
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- plane 1
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Background 0x2a
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "11000110", --  674 - 0x2a2  :  198 - 0xc6
    "11101110", --  675 - 0x2a3  :  238 - 0xee
    "00101000", --  676 - 0x2a4  :   40 - 0x28
    "00101000", --  677 - 0x2a5  :   40 - 0x28
    "00101000", --  678 - 0x2a6  :   40 - 0x28
    "00101000", --  679 - 0x2a7  :   40 - 0x28
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- plane 1
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00001000", --  688 - 0x2b0  :    8 - 0x8 -- Background 0x2b
    "00001000", --  689 - 0x2b1  :    8 - 0x8
    "00001000", --  690 - 0x2b2  :    8 - 0x8
    "00001000", --  691 - 0x2b3  :    8 - 0x8
    "00001110", --  692 - 0x2b4  :   14 - 0xe
    "00000110", --  693 - 0x2b5  :    6 - 0x6
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- plane 1
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00101000", --  704 - 0x2c0  :   40 - 0x28 -- Background 0x2c
    "00101000", --  705 - 0x2c1  :   40 - 0x28
    "00101000", --  706 - 0x2c2  :   40 - 0x28
    "00101000", --  707 - 0x2c3  :   40 - 0x28
    "11101110", --  708 - 0x2c4  :  238 - 0xee
    "11000110", --  709 - 0x2c5  :  198 - 0xc6
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- plane 1
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Background 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "01100000", --  722 - 0x2d2  :   96 - 0x60
    "01110000", --  723 - 0x2d3  :  112 - 0x70
    "00010000", --  724 - 0x2d4  :   16 - 0x10
    "00010000", --  725 - 0x2d5  :   16 - 0x10
    "00010000", --  726 - 0x2d6  :   16 - 0x10
    "00010000", --  727 - 0x2d7  :   16 - 0x10
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- plane 1
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00011100", --  736 - 0x2e0  :   28 - 0x1c -- Background 0x2e
    "00111110", --  737 - 0x2e1  :   62 - 0x3e
    "00111100", --  738 - 0x2e2  :   60 - 0x3c
    "00111000", --  739 - 0x2e3  :   56 - 0x38
    "00110000", --  740 - 0x2e4  :   48 - 0x30
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "01100000", --  742 - 0x2e6  :   96 - 0x60
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- plane 1
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00010000", --  752 - 0x2f0  :   16 - 0x10 -- Background 0x2f
    "00010000", --  753 - 0x2f1  :   16 - 0x10
    "00010000", --  754 - 0x2f2  :   16 - 0x10
    "00010000", --  755 - 0x2f3  :   16 - 0x10
    "01110000", --  756 - 0x2f4  :  112 - 0x70
    "01100000", --  757 - 0x2f5  :   96 - 0x60
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- plane 1
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "11111111", --  768 - 0x300  :  255 - 0xff -- Background 0x30
    "11111111", --  769 - 0x301  :  255 - 0xff
    "00111000", --  770 - 0x302  :   56 - 0x38
    "01101100", --  771 - 0x303  :  108 - 0x6c
    "11000110", --  772 - 0x304  :  198 - 0xc6
    "10000011", --  773 - 0x305  :  131 - 0x83
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "00000000", --  776 - 0x308  :    0 - 0x0 -- plane 1
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "11111111", --  784 - 0x310  :  255 - 0xff -- Background 0x31
    "00111000", --  785 - 0x311  :   56 - 0x38
    "01101100", --  786 - 0x312  :  108 - 0x6c
    "11000110", --  787 - 0x313  :  198 - 0xc6
    "10000011", --  788 - 0x314  :  131 - 0x83
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- plane 1
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00111000", --  800 - 0x320  :   56 - 0x38 -- Background 0x32
    "01101100", --  801 - 0x321  :  108 - 0x6c
    "11000110", --  802 - 0x322  :  198 - 0xc6
    "10000011", --  803 - 0x323  :  131 - 0x83
    "11111111", --  804 - 0x324  :  255 - 0xff
    "11111111", --  805 - 0x325  :  255 - 0xff
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- plane 1
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "01101100", --  816 - 0x330  :  108 - 0x6c -- Background 0x33
    "11000110", --  817 - 0x331  :  198 - 0xc6
    "10000011", --  818 - 0x332  :  131 - 0x83
    "11111111", --  819 - 0x333  :  255 - 0xff
    "11111111", --  820 - 0x334  :  255 - 0xff
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- plane 1
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "11000110", --  832 - 0x340  :  198 - 0xc6 -- Background 0x34
    "10000011", --  833 - 0x341  :  131 - 0x83
    "11111111", --  834 - 0x342  :  255 - 0xff
    "11111111", --  835 - 0x343  :  255 - 0xff
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- plane 1
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "10000011", --  848 - 0x350  :  131 - 0x83 -- Background 0x35
    "11111111", --  849 - 0x351  :  255 - 0xff
    "11111111", --  850 - 0x352  :  255 - 0xff
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- plane 1
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x36
    "11111111", --  865 - 0x361  :  255 - 0xff
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- plane 1
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "11111111", --  880 - 0x370  :  255 - 0xff -- Background 0x37
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- plane 1
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "11111111", --  903 - 0x387  :  255 - 0xff
    "00000000", --  904 - 0x388  :    0 - 0x0 -- plane 1
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x39
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "11111111", --  918 - 0x396  :  255 - 0xff
    "11111111", --  919 - 0x397  :  255 - 0xff
    "00000000", --  920 - 0x398  :    0 - 0x0 -- plane 1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "11111111", --  933 - 0x3a5  :  255 - 0xff
    "11111111", --  934 - 0x3a6  :  255 - 0xff
    "00111000", --  935 - 0x3a7  :   56 - 0x38
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "11111111", --  948 - 0x3b4  :  255 - 0xff
    "11111111", --  949 - 0x3b5  :  255 - 0xff
    "00111000", --  950 - 0x3b6  :   56 - 0x38
    "01101100", --  951 - 0x3b7  :  108 - 0x6c
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- plane 1
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "00111000", --  965 - 0x3c5  :   56 - 0x38
    "01101100", --  966 - 0x3c6  :  108 - 0x6c
    "11000110", --  967 - 0x3c7  :  198 - 0xc6
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "00111000", --  980 - 0x3d4  :   56 - 0x38
    "01101100", --  981 - 0x3d5  :  108 - 0x6c
    "11000110", --  982 - 0x3d6  :  198 - 0xc6
    "10000011", --  983 - 0x3d7  :  131 - 0x83
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- plane 1
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x3e
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "00111000", --  995 - 0x3e3  :   56 - 0x38
    "01101100", --  996 - 0x3e4  :  108 - 0x6c
    "11000110", --  997 - 0x3e5  :  198 - 0xc6
    "10000011", --  998 - 0x3e6  :  131 - 0x83
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "10000001", -- 1016 - 0x3f8  :  129 - 0x81 -- plane 1
    "11111111", -- 1017 - 0x3f9  :  255 - 0xff
    "10000001", -- 1018 - 0x3fa  :  129 - 0x81
    "10000001", -- 1019 - 0x3fb  :  129 - 0x81
    "10000001", -- 1020 - 0x3fc  :  129 - 0x81
    "11111111", -- 1021 - 0x3fd  :  255 - 0xff
    "10000001", -- 1022 - 0x3fe  :  129 - 0x81
    "10000001", -- 1023 - 0x3ff  :  129 - 0x81
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "11111111", -- 1031 - 0x407  :  255 - 0xff
    "10000001", -- 1032 - 0x408  :  129 - 0x81 -- plane 1
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "10000001", -- 1034 - 0x40a  :  129 - 0x81
    "10000001", -- 1035 - 0x40b  :  129 - 0x81
    "10000001", -- 1036 - 0x40c  :  129 - 0x81
    "11111111", -- 1037 - 0x40d  :  255 - 0xff
    "10000001", -- 1038 - 0x40e  :  129 - 0x81
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x41
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "11111111", -- 1045 - 0x415  :  255 - 0xff
    "11111111", -- 1046 - 0x416  :  255 - 0xff
    "00111000", -- 1047 - 0x417  :   56 - 0x38
    "10000001", -- 1048 - 0x418  :  129 - 0x81 -- plane 1
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "10000001", -- 1050 - 0x41a  :  129 - 0x81
    "10000001", -- 1051 - 0x41b  :  129 - 0x81
    "10000001", -- 1052 - 0x41c  :  129 - 0x81
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Background 0x42
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111111", -- 1061 - 0x425  :  255 - 0xff
    "00111000", -- 1062 - 0x426  :   56 - 0x38
    "01101100", -- 1063 - 0x427  :  108 - 0x6c
    "10000001", -- 1064 - 0x428  :  129 - 0x81 -- plane 1
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "10000001", -- 1066 - 0x42a  :  129 - 0x81
    "10000001", -- 1067 - 0x42b  :  129 - 0x81
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x43
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "00111000", -- 1077 - 0x435  :   56 - 0x38
    "01101100", -- 1078 - 0x436  :  108 - 0x6c
    "11000110", -- 1079 - 0x437  :  198 - 0xc6
    "10000001", -- 1080 - 0x438  :  129 - 0x81 -- plane 1
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "10000001", -- 1082 - 0x43a  :  129 - 0x81
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x44
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "11111111", -- 1090 - 0x442  :  255 - 0xff
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "00111000", -- 1092 - 0x444  :   56 - 0x38
    "01101100", -- 1093 - 0x445  :  108 - 0x6c
    "11000110", -- 1094 - 0x446  :  198 - 0xc6
    "10000011", -- 1095 - 0x447  :  131 - 0x83
    "10000001", -- 1096 - 0x448  :  129 - 0x81 -- plane 1
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x45
    "11111111", -- 1105 - 0x451  :  255 - 0xff
    "11111111", -- 1106 - 0x452  :  255 - 0xff
    "00111000", -- 1107 - 0x453  :   56 - 0x38
    "01101100", -- 1108 - 0x454  :  108 - 0x6c
    "11000110", -- 1109 - 0x455  :  198 - 0xc6
    "10000011", -- 1110 - 0x456  :  131 - 0x83
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "10000001", -- 1112 - 0x458  :  129 - 0x81 -- plane 1
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Background 0x46
    "00111000", -- 1121 - 0x461  :   56 - 0x38
    "01101100", -- 1122 - 0x462  :  108 - 0x6c
    "11000110", -- 1123 - 0x463  :  198 - 0xc6
    "10000011", -- 1124 - 0x464  :  131 - 0x83
    "11111111", -- 1125 - 0x465  :  255 - 0xff
    "11111111", -- 1126 - 0x466  :  255 - 0xff
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0 -- plane 1
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "10000001", -- 1135 - 0x46f  :  129 - 0x81
    "00111000", -- 1136 - 0x470  :   56 - 0x38 -- Background 0x47
    "01101100", -- 1137 - 0x471  :  108 - 0x6c
    "11000110", -- 1138 - 0x472  :  198 - 0xc6
    "10000011", -- 1139 - 0x473  :  131 - 0x83
    "11111111", -- 1140 - 0x474  :  255 - 0xff
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0 -- plane 1
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "10000001", -- 1150 - 0x47e  :  129 - 0x81
    "10000001", -- 1151 - 0x47f  :  129 - 0x81
    "01101100", -- 1152 - 0x480  :  108 - 0x6c -- Background 0x48
    "11000110", -- 1153 - 0x481  :  198 - 0xc6
    "10000011", -- 1154 - 0x482  :  131 - 0x83
    "11111111", -- 1155 - 0x483  :  255 - 0xff
    "11111111", -- 1156 - 0x484  :  255 - 0xff
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- plane 1
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "10000001", -- 1166 - 0x48e  :  129 - 0x81
    "10000001", -- 1167 - 0x48f  :  129 - 0x81
    "11000110", -- 1168 - 0x490  :  198 - 0xc6 -- Background 0x49
    "10000011", -- 1169 - 0x491  :  131 - 0x83
    "11111111", -- 1170 - 0x492  :  255 - 0xff
    "11111111", -- 1171 - 0x493  :  255 - 0xff
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- plane 1
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "10000001", -- 1180 - 0x49c  :  129 - 0x81
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "10000001", -- 1182 - 0x49e  :  129 - 0x81
    "10000001", -- 1183 - 0x49f  :  129 - 0x81
    "10000011", -- 1184 - 0x4a0  :  131 - 0x83 -- Background 0x4a
    "11111111", -- 1185 - 0x4a1  :  255 - 0xff
    "11111111", -- 1186 - 0x4a2  :  255 - 0xff
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "10000001", -- 1195 - 0x4ab  :  129 - 0x81
    "10000001", -- 1196 - 0x4ac  :  129 - 0x81
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "10000001", -- 1198 - 0x4ae  :  129 - 0x81
    "10000001", -- 1199 - 0x4af  :  129 - 0x81
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Background 0x4b
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "10000001", -- 1210 - 0x4ba  :  129 - 0x81
    "10000001", -- 1211 - 0x4bb  :  129 - 0x81
    "10000001", -- 1212 - 0x4bc  :  129 - 0x81
    "11111111", -- 1213 - 0x4bd  :  255 - 0xff
    "10000001", -- 1214 - 0x4be  :  129 - 0x81
    "10000001", -- 1215 - 0x4bf  :  129 - 0x81
    "10111111", -- 1216 - 0x4c0  :  191 - 0xbf -- Background 0x4c
    "01011111", -- 1217 - 0x4c1  :   95 - 0x5f
    "01011111", -- 1218 - 0x4c2  :   95 - 0x5f
    "01011111", -- 1219 - 0x4c3  :   95 - 0x5f
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "01011111", -- 1221 - 0x4c5  :   95 - 0x5f
    "01010001", -- 1222 - 0x4c6  :   81 - 0x51
    "01010101", -- 1223 - 0x4c7  :   85 - 0x55
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- plane 1
    "01111111", -- 1225 - 0x4c9  :  127 - 0x7f
    "01111111", -- 1226 - 0x4ca  :  127 - 0x7f
    "01111111", -- 1227 - 0x4cb  :  127 - 0x7f
    "01111111", -- 1228 - 0x4cc  :  127 - 0x7f
    "01111111", -- 1229 - 0x4cd  :  127 - 0x7f
    "01111111", -- 1230 - 0x4ce  :  127 - 0x7f
    "01111111", -- 1231 - 0x4cf  :  127 - 0x7f
    "01010001", -- 1232 - 0x4d0  :   81 - 0x51 -- Background 0x4d
    "01011111", -- 1233 - 0x4d1  :   95 - 0x5f
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "01011111", -- 1235 - 0x4d3  :   95 - 0x5f
    "01011111", -- 1236 - 0x4d4  :   95 - 0x5f
    "01011111", -- 1237 - 0x4d5  :   95 - 0x5f
    "01011111", -- 1238 - 0x4d6  :   95 - 0x5f
    "10111111", -- 1239 - 0x4d7  :  191 - 0xbf
    "01111111", -- 1240 - 0x4d8  :  127 - 0x7f -- plane 1
    "01111111", -- 1241 - 0x4d9  :  127 - 0x7f
    "01111111", -- 1242 - 0x4da  :  127 - 0x7f
    "01111111", -- 1243 - 0x4db  :  127 - 0x7f
    "01110010", -- 1244 - 0x4dc  :  114 - 0x72
    "01111111", -- 1245 - 0x4dd  :  127 - 0x7f
    "01111111", -- 1246 - 0x4de  :  127 - 0x7f
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Background 0x4e
    "11111110", -- 1249 - 0x4e1  :  254 - 0xfe
    "11111110", -- 1250 - 0x4e2  :  254 - 0xfe
    "11111110", -- 1251 - 0x4e3  :  254 - 0xfe
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "11111110", -- 1253 - 0x4e5  :  254 - 0xfe
    "00100110", -- 1254 - 0x4e6  :   38 - 0x26
    "00100110", -- 1255 - 0x4e7  :   38 - 0x26
    "11111111", -- 1256 - 0x4e8  :  255 - 0xff -- plane 1
    "11111110", -- 1257 - 0x4e9  :  254 - 0xfe
    "11111110", -- 1258 - 0x4ea  :  254 - 0xfe
    "11111110", -- 1259 - 0x4eb  :  254 - 0xfe
    "11111110", -- 1260 - 0x4ec  :  254 - 0xfe
    "11111110", -- 1261 - 0x4ed  :  254 - 0xfe
    "11111110", -- 1262 - 0x4ee  :  254 - 0xfe
    "11111110", -- 1263 - 0x4ef  :  254 - 0xfe
    "00100010", -- 1264 - 0x4f0  :   34 - 0x22 -- Background 0x4f
    "11111110", -- 1265 - 0x4f1  :  254 - 0xfe
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "11111110", -- 1267 - 0x4f3  :  254 - 0xfe
    "11111110", -- 1268 - 0x4f4  :  254 - 0xfe
    "11111110", -- 1269 - 0x4f5  :  254 - 0xfe
    "11111110", -- 1270 - 0x4f6  :  254 - 0xfe
    "11111111", -- 1271 - 0x4f7  :  255 - 0xff
    "11111110", -- 1272 - 0x4f8  :  254 - 0xfe -- plane 1
    "11111110", -- 1273 - 0x4f9  :  254 - 0xfe
    "11111110", -- 1274 - 0x4fa  :  254 - 0xfe
    "11111110", -- 1275 - 0x4fb  :  254 - 0xfe
    "01001010", -- 1276 - 0x4fc  :   74 - 0x4a
    "11111110", -- 1277 - 0x4fd  :  254 - 0xfe
    "11111110", -- 1278 - 0x4fe  :  254 - 0xfe
    "11111111", -- 1279 - 0x4ff  :  255 - 0xff
    "00000111", -- 1280 - 0x500  :    7 - 0x7 -- Background 0x50
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00001111", -- 1282 - 0x502  :   15 - 0xf
    "00011111", -- 1283 - 0x503  :   31 - 0x1f
    "00011111", -- 1284 - 0x504  :   31 - 0x1f
    "00011111", -- 1285 - 0x505  :   31 - 0x1f
    "00011111", -- 1286 - 0x506  :   31 - 0x1f
    "00011111", -- 1287 - 0x507  :   31 - 0x1f
    "00000101", -- 1288 - 0x508  :    5 - 0x5 -- plane 1
    "00001111", -- 1289 - 0x509  :   15 - 0xf
    "00001011", -- 1290 - 0x50a  :   11 - 0xb
    "00011011", -- 1291 - 0x50b  :   27 - 0x1b
    "00010011", -- 1292 - 0x50c  :   19 - 0x13
    "00010011", -- 1293 - 0x50d  :   19 - 0x13
    "00010011", -- 1294 - 0x50e  :   19 - 0x13
    "00010011", -- 1295 - 0x50f  :   19 - 0x13
    "00011111", -- 1296 - 0x510  :   31 - 0x1f -- Background 0x51
    "00011111", -- 1297 - 0x511  :   31 - 0x1f
    "00011111", -- 1298 - 0x512  :   31 - 0x1f
    "00011111", -- 1299 - 0x513  :   31 - 0x1f
    "00011111", -- 1300 - 0x514  :   31 - 0x1f
    "00001111", -- 1301 - 0x515  :   15 - 0xf
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000111", -- 1303 - 0x517  :    7 - 0x7
    "00010011", -- 1304 - 0x518  :   19 - 0x13 -- plane 1
    "00010011", -- 1305 - 0x519  :   19 - 0x13
    "00010011", -- 1306 - 0x51a  :   19 - 0x13
    "00010011", -- 1307 - 0x51b  :   19 - 0x13
    "00011011", -- 1308 - 0x51c  :   27 - 0x1b
    "00001011", -- 1309 - 0x51d  :   11 - 0xb
    "00001111", -- 1310 - 0x51e  :   15 - 0xf
    "00000101", -- 1311 - 0x51f  :    5 - 0x5
    "00000111", -- 1312 - 0x520  :    7 - 0x7 -- Background 0x52
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00001111", -- 1314 - 0x522  :   15 - 0xf
    "00011111", -- 1315 - 0x523  :   31 - 0x1f
    "00011111", -- 1316 - 0x524  :   31 - 0x1f
    "00011111", -- 1317 - 0x525  :   31 - 0x1f
    "00011111", -- 1318 - 0x526  :   31 - 0x1f
    "00011111", -- 1319 - 0x527  :   31 - 0x1f
    "00000101", -- 1320 - 0x528  :    5 - 0x5 -- plane 1
    "00001111", -- 1321 - 0x529  :   15 - 0xf
    "00001011", -- 1322 - 0x52a  :   11 - 0xb
    "00011011", -- 1323 - 0x52b  :   27 - 0x1b
    "00010011", -- 1324 - 0x52c  :   19 - 0x13
    "00010011", -- 1325 - 0x52d  :   19 - 0x13
    "00010011", -- 1326 - 0x52e  :   19 - 0x13
    "00010011", -- 1327 - 0x52f  :   19 - 0x13
    "00011111", -- 1328 - 0x530  :   31 - 0x1f -- Background 0x53
    "00011111", -- 1329 - 0x531  :   31 - 0x1f
    "00011111", -- 1330 - 0x532  :   31 - 0x1f
    "00011111", -- 1331 - 0x533  :   31 - 0x1f
    "00011111", -- 1332 - 0x534  :   31 - 0x1f
    "00001111", -- 1333 - 0x535  :   15 - 0xf
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000111", -- 1335 - 0x537  :    7 - 0x7
    "00010011", -- 1336 - 0x538  :   19 - 0x13 -- plane 1
    "00010011", -- 1337 - 0x539  :   19 - 0x13
    "00010011", -- 1338 - 0x53a  :   19 - 0x13
    "00010011", -- 1339 - 0x53b  :   19 - 0x13
    "00011011", -- 1340 - 0x53c  :   27 - 0x1b
    "00001011", -- 1341 - 0x53d  :   11 - 0xb
    "00001111", -- 1342 - 0x53e  :   15 - 0xf
    "00000101", -- 1343 - 0x53f  :    5 - 0x5
    "11100000", -- 1344 - 0x540  :  224 - 0xe0 -- Background 0x54
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "11110001", -- 1346 - 0x542  :  241 - 0xf1
    "11111011", -- 1347 - 0x543  :  251 - 0xfb
    "11111011", -- 1348 - 0x544  :  251 - 0xfb
    "11111011", -- 1349 - 0x545  :  251 - 0xfb
    "11111011", -- 1350 - 0x546  :  251 - 0xfb
    "11111011", -- 1351 - 0x547  :  251 - 0xfb
    "10100000", -- 1352 - 0x548  :  160 - 0xa0 -- plane 1
    "11110001", -- 1353 - 0x549  :  241 - 0xf1
    "11010001", -- 1354 - 0x54a  :  209 - 0xd1
    "11011011", -- 1355 - 0x54b  :  219 - 0xdb
    "11001010", -- 1356 - 0x54c  :  202 - 0xca
    "11001010", -- 1357 - 0x54d  :  202 - 0xca
    "11001010", -- 1358 - 0x54e  :  202 - 0xca
    "11001010", -- 1359 - 0x54f  :  202 - 0xca
    "11111011", -- 1360 - 0x550  :  251 - 0xfb -- Background 0x55
    "11111011", -- 1361 - 0x551  :  251 - 0xfb
    "11111011", -- 1362 - 0x552  :  251 - 0xfb
    "11111011", -- 1363 - 0x553  :  251 - 0xfb
    "11111011", -- 1364 - 0x554  :  251 - 0xfb
    "11110001", -- 1365 - 0x555  :  241 - 0xf1
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "11100000", -- 1367 - 0x557  :  224 - 0xe0
    "11001010", -- 1368 - 0x558  :  202 - 0xca -- plane 1
    "11001010", -- 1369 - 0x559  :  202 - 0xca
    "11001010", -- 1370 - 0x55a  :  202 - 0xca
    "11001010", -- 1371 - 0x55b  :  202 - 0xca
    "11011011", -- 1372 - 0x55c  :  219 - 0xdb
    "11010001", -- 1373 - 0x55d  :  209 - 0xd1
    "11110001", -- 1374 - 0x55e  :  241 - 0xf1
    "10100000", -- 1375 - 0x55f  :  160 - 0xa0
    "11100000", -- 1376 - 0x560  :  224 - 0xe0 -- Background 0x56
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "11110001", -- 1378 - 0x562  :  241 - 0xf1
    "11111011", -- 1379 - 0x563  :  251 - 0xfb
    "11111011", -- 1380 - 0x564  :  251 - 0xfb
    "11111011", -- 1381 - 0x565  :  251 - 0xfb
    "11111011", -- 1382 - 0x566  :  251 - 0xfb
    "11111011", -- 1383 - 0x567  :  251 - 0xfb
    "10100000", -- 1384 - 0x568  :  160 - 0xa0 -- plane 1
    "11110001", -- 1385 - 0x569  :  241 - 0xf1
    "11010001", -- 1386 - 0x56a  :  209 - 0xd1
    "11011011", -- 1387 - 0x56b  :  219 - 0xdb
    "11001010", -- 1388 - 0x56c  :  202 - 0xca
    "11001010", -- 1389 - 0x56d  :  202 - 0xca
    "11001010", -- 1390 - 0x56e  :  202 - 0xca
    "11001010", -- 1391 - 0x56f  :  202 - 0xca
    "11111011", -- 1392 - 0x570  :  251 - 0xfb -- Background 0x57
    "11111011", -- 1393 - 0x571  :  251 - 0xfb
    "11111011", -- 1394 - 0x572  :  251 - 0xfb
    "11111011", -- 1395 - 0x573  :  251 - 0xfb
    "11111011", -- 1396 - 0x574  :  251 - 0xfb
    "11110001", -- 1397 - 0x575  :  241 - 0xf1
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "11100000", -- 1399 - 0x577  :  224 - 0xe0
    "11001010", -- 1400 - 0x578  :  202 - 0xca -- plane 1
    "11001010", -- 1401 - 0x579  :  202 - 0xca
    "11001010", -- 1402 - 0x57a  :  202 - 0xca
    "11001010", -- 1403 - 0x57b  :  202 - 0xca
    "11011011", -- 1404 - 0x57c  :  219 - 0xdb
    "11010001", -- 1405 - 0x57d  :  209 - 0xd1
    "11110000", -- 1406 - 0x57e  :  240 - 0xf0
    "10100000", -- 1407 - 0x57f  :  160 - 0xa0
    "11111100", -- 1408 - 0x580  :  252 - 0xfc -- Background 0x58
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "11111110", -- 1410 - 0x582  :  254 - 0xfe
    "11111111", -- 1411 - 0x583  :  255 - 0xff
    "11111111", -- 1412 - 0x584  :  255 - 0xff
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "10110100", -- 1416 - 0x588  :  180 - 0xb4 -- plane 1
    "11111110", -- 1417 - 0x589  :  254 - 0xfe
    "01111010", -- 1418 - 0x58a  :  122 - 0x7a
    "01111011", -- 1419 - 0x58b  :  123 - 0x7b
    "01111001", -- 1420 - 0x58c  :  121 - 0x79
    "01111001", -- 1421 - 0x58d  :  121 - 0x79
    "01111001", -- 1422 - 0x58e  :  121 - 0x79
    "01111001", -- 1423 - 0x58f  :  121 - 0x79
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Background 0x59
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "11111111", -- 1426 - 0x592  :  255 - 0xff
    "11111111", -- 1427 - 0x593  :  255 - 0xff
    "11111111", -- 1428 - 0x594  :  255 - 0xff
    "11111110", -- 1429 - 0x595  :  254 - 0xfe
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "11111100", -- 1431 - 0x597  :  252 - 0xfc
    "01111001", -- 1432 - 0x598  :  121 - 0x79 -- plane 1
    "01111001", -- 1433 - 0x599  :  121 - 0x79
    "01111001", -- 1434 - 0x59a  :  121 - 0x79
    "01111001", -- 1435 - 0x59b  :  121 - 0x79
    "01111011", -- 1436 - 0x59c  :  123 - 0x7b
    "01111010", -- 1437 - 0x59d  :  122 - 0x7a
    "11111110", -- 1438 - 0x59e  :  254 - 0xfe
    "10110100", -- 1439 - 0x59f  :  180 - 0xb4
    "11111100", -- 1440 - 0x5a0  :  252 - 0xfc -- Background 0x5a
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "11111110", -- 1442 - 0x5a2  :  254 - 0xfe
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "11111111", -- 1445 - 0x5a5  :  255 - 0xff
    "11111111", -- 1446 - 0x5a6  :  255 - 0xff
    "11111111", -- 1447 - 0x5a7  :  255 - 0xff
    "10110100", -- 1448 - 0x5a8  :  180 - 0xb4 -- plane 1
    "11111110", -- 1449 - 0x5a9  :  254 - 0xfe
    "01111010", -- 1450 - 0x5aa  :  122 - 0x7a
    "01111011", -- 1451 - 0x5ab  :  123 - 0x7b
    "01111001", -- 1452 - 0x5ac  :  121 - 0x79
    "01111001", -- 1453 - 0x5ad  :  121 - 0x79
    "01111001", -- 1454 - 0x5ae  :  121 - 0x79
    "01111001", -- 1455 - 0x5af  :  121 - 0x79
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Background 0x5b
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11111110", -- 1461 - 0x5b5  :  254 - 0xfe
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "11111100", -- 1463 - 0x5b7  :  252 - 0xfc
    "01111001", -- 1464 - 0x5b8  :  121 - 0x79 -- plane 1
    "01111001", -- 1465 - 0x5b9  :  121 - 0x79
    "01111001", -- 1466 - 0x5ba  :  121 - 0x79
    "01111001", -- 1467 - 0x5bb  :  121 - 0x79
    "01111011", -- 1468 - 0x5bc  :  123 - 0x7b
    "01111010", -- 1469 - 0x5bd  :  122 - 0x7a
    "11111110", -- 1470 - 0x5be  :  254 - 0xfe
    "10110100", -- 1471 - 0x5bf  :  180 - 0xb4
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00011111", -- 1474 - 0x5c2  :   31 - 0x1f
    "00010000", -- 1475 - 0x5c3  :   16 - 0x10
    "00010000", -- 1476 - 0x5c4  :   16 - 0x10
    "00011111", -- 1477 - 0x5c5  :   31 - 0x1f
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "01111111", -- 1480 - 0x5c8  :  127 - 0x7f -- plane 1
    "10111111", -- 1481 - 0x5c9  :  191 - 0xbf
    "11111111", -- 1482 - 0x5ca  :  255 - 0xff
    "10110010", -- 1483 - 0x5cb  :  178 - 0xb2
    "10110001", -- 1484 - 0x5cc  :  177 - 0xb1
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "10111111", -- 1486 - 0x5ce  :  191 - 0xbf
    "01111111", -- 1487 - 0x5cf  :  127 - 0x7f
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "11111000", -- 1490 - 0x5d2  :  248 - 0xf8
    "00001000", -- 1491 - 0x5d3  :    8 - 0x8
    "00001000", -- 1492 - 0x5d4  :    8 - 0x8
    "11111000", -- 1493 - 0x5d5  :  248 - 0xf8
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "11111110", -- 1496 - 0x5d8  :  254 - 0xfe -- plane 1
    "11111101", -- 1497 - 0x5d9  :  253 - 0xfd
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11001101", -- 1499 - 0x5db  :  205 - 0xcd
    "01101101", -- 1500 - 0x5dc  :  109 - 0x6d
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111101", -- 1502 - 0x5de  :  253 - 0xfd
    "11111110", -- 1503 - 0x5df  :  254 - 0xfe
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0x5e
    "00000001", -- 1505 - 0x5e1  :    1 - 0x1
    "00000010", -- 1506 - 0x5e2  :    2 - 0x2
    "00000010", -- 1507 - 0x5e3  :    2 - 0x2
    "11110001", -- 1508 - 0x5e4  :  241 - 0xf1
    "00001000", -- 1509 - 0x5e5  :    8 - 0x8
    "00000100", -- 1510 - 0x5e6  :    4 - 0x4
    "00000011", -- 1511 - 0x5e7  :    3 - 0x3
    "11111111", -- 1512 - 0x5e8  :  255 - 0xff -- plane 1
    "11111111", -- 1513 - 0x5e9  :  255 - 0xff
    "10101110", -- 1514 - 0x5ea  :  174 - 0xae
    "11111110", -- 1515 - 0x5eb  :  254 - 0xfe
    "11111111", -- 1516 - 0x5ec  :  255 - 0xff
    "00001111", -- 1517 - 0x5ed  :   15 - 0xf
    "00000111", -- 1518 - 0x5ee  :    7 - 0x7
    "00000011", -- 1519 - 0x5ef  :    3 - 0x3
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0x5f
    "10000000", -- 1521 - 0x5f1  :  128 - 0x80
    "01000000", -- 1522 - 0x5f2  :   64 - 0x40
    "01000000", -- 1523 - 0x5f3  :   64 - 0x40
    "10001111", -- 1524 - 0x5f4  :  143 - 0x8f
    "00010000", -- 1525 - 0x5f5  :   16 - 0x10
    "00100000", -- 1526 - 0x5f6  :   32 - 0x20
    "11000000", -- 1527 - 0x5f7  :  192 - 0xc0
    "11111111", -- 1528 - 0x5f8  :  255 - 0xff -- plane 1
    "11111111", -- 1529 - 0x5f9  :  255 - 0xff
    "01110101", -- 1530 - 0x5fa  :  117 - 0x75
    "01111111", -- 1531 - 0x5fb  :  127 - 0x7f
    "11111111", -- 1532 - 0x5fc  :  255 - 0xff
    "11110000", -- 1533 - 0x5fd  :  240 - 0xf0
    "11100000", -- 1534 - 0x5fe  :  224 - 0xe0
    "11000000", -- 1535 - 0x5ff  :  192 - 0xc0
    "00000011", -- 1536 - 0x600  :    3 - 0x3 -- Background 0x60
    "00000100", -- 1537 - 0x601  :    4 - 0x4
    "00001000", -- 1538 - 0x602  :    8 - 0x8
    "11110001", -- 1539 - 0x603  :  241 - 0xf1
    "00000010", -- 1540 - 0x604  :    2 - 0x2
    "00000010", -- 1541 - 0x605  :    2 - 0x2
    "00000001", -- 1542 - 0x606  :    1 - 0x1
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000011", -- 1544 - 0x608  :    3 - 0x3 -- plane 1
    "00000111", -- 1545 - 0x609  :    7 - 0x7
    "00001111", -- 1546 - 0x60a  :   15 - 0xf
    "11111111", -- 1547 - 0x60b  :  255 - 0xff
    "11111110", -- 1548 - 0x60c  :  254 - 0xfe
    "10101110", -- 1549 - 0x60d  :  174 - 0xae
    "11111111", -- 1550 - 0x60e  :  255 - 0xff
    "11111111", -- 1551 - 0x60f  :  255 - 0xff
    "11000000", -- 1552 - 0x610  :  192 - 0xc0 -- Background 0x61
    "00100000", -- 1553 - 0x611  :   32 - 0x20
    "00010000", -- 1554 - 0x612  :   16 - 0x10
    "10001111", -- 1555 - 0x613  :  143 - 0x8f
    "01000000", -- 1556 - 0x614  :   64 - 0x40
    "01000000", -- 1557 - 0x615  :   64 - 0x40
    "10000000", -- 1558 - 0x616  :  128 - 0x80
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "11000000", -- 1560 - 0x618  :  192 - 0xc0 -- plane 1
    "11100000", -- 1561 - 0x619  :  224 - 0xe0
    "11110000", -- 1562 - 0x61a  :  240 - 0xf0
    "11111111", -- 1563 - 0x61b  :  255 - 0xff
    "01111111", -- 1564 - 0x61c  :  127 - 0x7f
    "01110101", -- 1565 - 0x61d  :  117 - 0x75
    "11111111", -- 1566 - 0x61e  :  255 - 0xff
    "11111111", -- 1567 - 0x61f  :  255 - 0xff
    "11111111", -- 1568 - 0x620  :  255 - 0xff -- Background 0x62
    "11111111", -- 1569 - 0x621  :  255 - 0xff
    "11000011", -- 1570 - 0x622  :  195 - 0xc3
    "10000001", -- 1571 - 0x623  :  129 - 0x81
    "10000001", -- 1572 - 0x624  :  129 - 0x81
    "11000011", -- 1573 - 0x625  :  195 - 0xc3
    "11111111", -- 1574 - 0x626  :  255 - 0xff
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "11111111", -- 1576 - 0x628  :  255 - 0xff -- plane 1
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "11000011", -- 1578 - 0x62a  :  195 - 0xc3
    "10000001", -- 1579 - 0x62b  :  129 - 0x81
    "10000001", -- 1580 - 0x62c  :  129 - 0x81
    "11000011", -- 1581 - 0x62d  :  195 - 0xc3
    "11111111", -- 1582 - 0x62e  :  255 - 0xff
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "11111111", -- 1584 - 0x630  :  255 - 0xff -- Background 0x63
    "10011001", -- 1585 - 0x631  :  153 - 0x99
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "10000001", -- 1589 - 0x635  :  129 - 0x81
    "10000001", -- 1590 - 0x636  :  129 - 0x81
    "10000001", -- 1591 - 0x637  :  129 - 0x81
    "10000001", -- 1592 - 0x638  :  129 - 0x81 -- plane 1
    "01100110", -- 1593 - 0x639  :  102 - 0x66
    "01111110", -- 1594 - 0x63a  :  126 - 0x7e
    "01111110", -- 1595 - 0x63b  :  126 - 0x7e
    "01111110", -- 1596 - 0x63c  :  126 - 0x7e
    "11111111", -- 1597 - 0x63d  :  255 - 0xff
    "11111111", -- 1598 - 0x63e  :  255 - 0xff
    "01111110", -- 1599 - 0x63f  :  126 - 0x7e
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "01100000", -- 1604 - 0x644  :   96 - 0x60
    "01100000", -- 1605 - 0x645  :   96 - 0x60
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- plane 1
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Background 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "01101100", -- 1620 - 0x654  :  108 - 0x6c
    "01101100", -- 1621 - 0x655  :  108 - 0x6c
    "00001000", -- 1622 - 0x656  :    8 - 0x8
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- plane 1
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00111100", -- 1632 - 0x660  :   60 - 0x3c -- Background 0x66
    "00011000", -- 1633 - 0x661  :   24 - 0x18
    "00011000", -- 1634 - 0x662  :   24 - 0x18
    "00011000", -- 1635 - 0x663  :   24 - 0x18
    "00011000", -- 1636 - 0x664  :   24 - 0x18
    "00011000", -- 1637 - 0x665  :   24 - 0x18
    "00111100", -- 1638 - 0x666  :   60 - 0x3c
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- plane 1
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11111111", -- 1648 - 0x670  :  255 - 0xff -- Background 0x67
    "01100110", -- 1649 - 0x671  :  102 - 0x66
    "01100110", -- 1650 - 0x672  :  102 - 0x66
    "01100110", -- 1651 - 0x673  :  102 - 0x66
    "01100110", -- 1652 - 0x674  :  102 - 0x66
    "01100110", -- 1653 - 0x675  :  102 - 0x66
    "01100110", -- 1654 - 0x676  :  102 - 0x66
    "11111111", -- 1655 - 0x677  :  255 - 0xff
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- plane 1
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000011", -- 1664 - 0x680  :    3 - 0x3 -- Background 0x68
    "00000001", -- 1665 - 0x681  :    1 - 0x1
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000011", -- 1672 - 0x688  :    3 - 0x3 -- plane 1
    "00000001", -- 1673 - 0x689  :    1 - 0x1
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "10000011", -- 1680 - 0x690  :  131 - 0x83 -- Background 0x69
    "11010001", -- 1681 - 0x691  :  209 - 0xd1
    "11100001", -- 1682 - 0x692  :  225 - 0xe1
    "11010001", -- 1683 - 0x693  :  209 - 0xd1
    "00000010", -- 1684 - 0x694  :    2 - 0x2
    "10000100", -- 1685 - 0x695  :  132 - 0x84
    "11110000", -- 1686 - 0x696  :  240 - 0xf0
    "11001110", -- 1687 - 0x697  :  206 - 0xce
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- plane 1
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111111", -- 1692 - 0x69c  :  255 - 0xff
    "11111111", -- 1693 - 0x69d  :  255 - 0xff
    "11111111", -- 1694 - 0x69e  :  255 - 0xff
    "11111111", -- 1695 - 0x69f  :  255 - 0xff
    "11000000", -- 1696 - 0x6a0  :  192 - 0xc0 -- Background 0x6a
    "10000000", -- 1697 - 0x6a1  :  128 - 0x80
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "11000000", -- 1704 - 0x6a8  :  192 - 0xc0 -- plane 1
    "10000000", -- 1705 - 0x6a9  :  128 - 0x80
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "11000001", -- 1712 - 0x6b0  :  193 - 0xc1 -- Background 0x6b
    "10001011", -- 1713 - 0x6b1  :  139 - 0x8b
    "10000111", -- 1714 - 0x6b2  :  135 - 0x87
    "10001011", -- 1715 - 0x6b3  :  139 - 0x8b
    "01000000", -- 1716 - 0x6b4  :   64 - 0x40
    "00100001", -- 1717 - 0x6b5  :   33 - 0x21
    "00001111", -- 1718 - 0x6b6  :   15 - 0xf
    "11010011", -- 1719 - 0x6b7  :  211 - 0xd3
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- plane 1
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111111", -- 1723 - 0x6bb  :  255 - 0xff
    "11111111", -- 1724 - 0x6bc  :  255 - 0xff
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Background 0x6c
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "00011111", -- 1731 - 0x6c3  :   31 - 0x1f
    "00001111", -- 1732 - 0x6c4  :   15 - 0xf
    "00011110", -- 1733 - 0x6c5  :   30 - 0x1e
    "00111111", -- 1734 - 0x6c6  :   63 - 0x3f
    "01111111", -- 1735 - 0x6c7  :  127 - 0x7f
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- plane 1
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "00011111", -- 1739 - 0x6cb  :   31 - 0x1f
    "00011111", -- 1740 - 0x6cc  :   31 - 0x1f
    "00111111", -- 1741 - 0x6cd  :   63 - 0x3f
    "01111111", -- 1742 - 0x6ce  :  127 - 0x7f
    "11111111", -- 1743 - 0x6cf  :  255 - 0xff
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Background 0x6d
    "11111111", -- 1745 - 0x6d1  :  255 - 0xff
    "11111111", -- 1746 - 0x6d2  :  255 - 0xff
    "11111000", -- 1747 - 0x6d3  :  248 - 0xf8
    "11110000", -- 1748 - 0x6d4  :  240 - 0xf0
    "01111000", -- 1749 - 0x6d5  :  120 - 0x78
    "11111100", -- 1750 - 0x6d6  :  252 - 0xfc
    "11111110", -- 1751 - 0x6d7  :  254 - 0xfe
    "11111111", -- 1752 - 0x6d8  :  255 - 0xff -- plane 1
    "11111111", -- 1753 - 0x6d9  :  255 - 0xff
    "11111111", -- 1754 - 0x6da  :  255 - 0xff
    "11111000", -- 1755 - 0x6db  :  248 - 0xf8
    "11111000", -- 1756 - 0x6dc  :  248 - 0xf8
    "11111100", -- 1757 - 0x6dd  :  252 - 0xfc
    "11111110", -- 1758 - 0x6de  :  254 - 0xfe
    "11111111", -- 1759 - 0x6df  :  255 - 0xff
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00111100", -- 1765 - 0x6e5  :   60 - 0x3c
    "01000010", -- 1766 - 0x6e6  :   66 - 0x42
    "10000001", -- 1767 - 0x6e7  :  129 - 0x81
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00111100", -- 1773 - 0x6ed  :   60 - 0x3c
    "01000010", -- 1774 - 0x6ee  :   66 - 0x42
    "10000001", -- 1775 - 0x6ef  :  129 - 0x81
    "10000001", -- 1776 - 0x6f0  :  129 - 0x81 -- Background 0x6f
    "10111101", -- 1777 - 0x6f1  :  189 - 0xbd
    "01111110", -- 1778 - 0x6f2  :  126 - 0x7e
    "11111111", -- 1779 - 0x6f3  :  255 - 0xff
    "11100111", -- 1780 - 0x6f4  :  231 - 0xe7
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "10000001", -- 1784 - 0x6f8  :  129 - 0x81 -- plane 1
    "10111101", -- 1785 - 0x6f9  :  189 - 0xbd
    "01111110", -- 1786 - 0x6fa  :  126 - 0x7e
    "10100101", -- 1787 - 0x6fb  :  165 - 0xa5
    "11011011", -- 1788 - 0x6fc  :  219 - 0xdb
    "11100111", -- 1789 - 0x6fd  :  231 - 0xe7
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111111", -- 1791 - 0x6ff  :  255 - 0xff
    "00000001", -- 1792 - 0x700  :    1 - 0x1 -- Background 0x70
    "00000111", -- 1793 - 0x701  :    7 - 0x7
    "00011111", -- 1794 - 0x702  :   31 - 0x1f
    "00111111", -- 1795 - 0x703  :   63 - 0x3f
    "01111111", -- 1796 - 0x704  :  127 - 0x7f
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11011101", -- 1799 - 0x707  :  221 - 0xdd
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- plane 1
    "00000101", -- 1801 - 0x709  :    5 - 0x5
    "00011001", -- 1802 - 0x70a  :   25 - 0x19
    "00110011", -- 1803 - 0x70b  :   51 - 0x33
    "01100011", -- 1804 - 0x70c  :   99 - 0x63
    "11000111", -- 1805 - 0x70d  :  199 - 0xc7
    "11000111", -- 1806 - 0x70e  :  199 - 0xc7
    "11000100", -- 1807 - 0x70f  :  196 - 0xc4
    "10001001", -- 1808 - 0x710  :  137 - 0x89 -- Background 0x71
    "00000001", -- 1809 - 0x711  :    1 - 0x1
    "00000001", -- 1810 - 0x712  :    1 - 0x1
    "00000001", -- 1811 - 0x713  :    1 - 0x1
    "00000001", -- 1812 - 0x714  :    1 - 0x1
    "00000001", -- 1813 - 0x715  :    1 - 0x1
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "10000000", -- 1816 - 0x718  :  128 - 0x80 -- plane 1
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000001", -- 1819 - 0x71b  :    1 - 0x1
    "00000001", -- 1820 - 0x71c  :    1 - 0x1
    "00000001", -- 1821 - 0x71d  :    1 - 0x1
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "10000000", -- 1824 - 0x720  :  128 - 0x80 -- Background 0x72
    "11100000", -- 1825 - 0x721  :  224 - 0xe0
    "11111000", -- 1826 - 0x722  :  248 - 0xf8
    "11111100", -- 1827 - 0x723  :  252 - 0xfc
    "11111110", -- 1828 - 0x724  :  254 - 0xfe
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "00111011", -- 1831 - 0x727  :   59 - 0x3b
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- plane 1
    "10100000", -- 1833 - 0x729  :  160 - 0xa0
    "10011000", -- 1834 - 0x72a  :  152 - 0x98
    "11001100", -- 1835 - 0x72b  :  204 - 0xcc
    "11000110", -- 1836 - 0x72c  :  198 - 0xc6
    "11100011", -- 1837 - 0x72d  :  227 - 0xe3
    "11100011", -- 1838 - 0x72e  :  227 - 0xe3
    "00100011", -- 1839 - 0x72f  :   35 - 0x23
    "00010001", -- 1840 - 0x730  :   17 - 0x11 -- Background 0x73
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "01000000", -- 1845 - 0x735  :   64 - 0x40
    "10000000", -- 1846 - 0x736  :  128 - 0x80
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000001", -- 1848 - 0x738  :    1 - 0x1 -- plane 1
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "01000000", -- 1853 - 0x73d  :   64 - 0x40
    "10000000", -- 1854 - 0x73e  :  128 - 0x80
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000001", -- 1856 - 0x740  :    1 - 0x1 -- Background 0x74
    "00000001", -- 1857 - 0x741  :    1 - 0x1
    "00000001", -- 1858 - 0x742  :    1 - 0x1
    "00000001", -- 1859 - 0x743  :    1 - 0x1
    "00000001", -- 1860 - 0x744  :    1 - 0x1
    "00000001", -- 1861 - 0x745  :    1 - 0x1
    "00000001", -- 1862 - 0x746  :    1 - 0x1
    "00000001", -- 1863 - 0x747  :    1 - 0x1
    "00000001", -- 1864 - 0x748  :    1 - 0x1 -- plane 1
    "00000001", -- 1865 - 0x749  :    1 - 0x1
    "00000001", -- 1866 - 0x74a  :    1 - 0x1
    "00000001", -- 1867 - 0x74b  :    1 - 0x1
    "00000001", -- 1868 - 0x74c  :    1 - 0x1
    "00000001", -- 1869 - 0x74d  :    1 - 0x1
    "00000001", -- 1870 - 0x74e  :    1 - 0x1
    "00000001", -- 1871 - 0x74f  :    1 - 0x1
    "10000000", -- 1872 - 0x750  :  128 - 0x80 -- Background 0x75
    "10000000", -- 1873 - 0x751  :  128 - 0x80
    "10000000", -- 1874 - 0x752  :  128 - 0x80
    "10000000", -- 1875 - 0x753  :  128 - 0x80
    "10000000", -- 1876 - 0x754  :  128 - 0x80
    "10000000", -- 1877 - 0x755  :  128 - 0x80
    "10000000", -- 1878 - 0x756  :  128 - 0x80
    "10000000", -- 1879 - 0x757  :  128 - 0x80
    "10000000", -- 1880 - 0x758  :  128 - 0x80 -- plane 1
    "10000000", -- 1881 - 0x759  :  128 - 0x80
    "10000000", -- 1882 - 0x75a  :  128 - 0x80
    "10000000", -- 1883 - 0x75b  :  128 - 0x80
    "10000000", -- 1884 - 0x75c  :  128 - 0x80
    "10000000", -- 1885 - 0x75d  :  128 - 0x80
    "10000000", -- 1886 - 0x75e  :  128 - 0x80
    "10000000", -- 1887 - 0x75f  :  128 - 0x80
    "00000001", -- 1888 - 0x760  :    1 - 0x1 -- Background 0x76
    "00000011", -- 1889 - 0x761  :    3 - 0x3
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000011", -- 1892 - 0x764  :    3 - 0x3
    "00011001", -- 1893 - 0x765  :   25 - 0x19
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000001", -- 1896 - 0x768  :    1 - 0x1 -- plane 1
    "00000011", -- 1897 - 0x769  :    3 - 0x3
    "00000011", -- 1898 - 0x76a  :    3 - 0x3
    "00000111", -- 1899 - 0x76b  :    7 - 0x7
    "00000100", -- 1900 - 0x76c  :    4 - 0x4
    "00011100", -- 1901 - 0x76d  :   28 - 0x1c
    "00111111", -- 1902 - 0x76e  :   63 - 0x3f
    "01111111", -- 1903 - 0x76f  :  127 - 0x7f
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "01111100", -- 1906 - 0x772  :  124 - 0x7c
    "00000010", -- 1907 - 0x773  :    2 - 0x2
    "00000001", -- 1908 - 0x774  :    1 - 0x1
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "01111111", -- 1912 - 0x778  :  127 - 0x7f -- plane 1
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111111", -- 1914 - 0x77a  :  255 - 0xff
    "01111111", -- 1915 - 0x77b  :  127 - 0x7f
    "01111111", -- 1916 - 0x77c  :  127 - 0x7f
    "00011111", -- 1917 - 0x77d  :   31 - 0x1f
    "00000011", -- 1918 - 0x77e  :    3 - 0x3
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000001", -- 1922 - 0x782  :    1 - 0x1
    "00000001", -- 1923 - 0x783  :    1 - 0x1
    "00000011", -- 1924 - 0x784  :    3 - 0x3
    "00000111", -- 1925 - 0x785  :    7 - 0x7
    "00000111", -- 1926 - 0x786  :    7 - 0x7
    "00001111", -- 1927 - 0x787  :   15 - 0xf
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- plane 1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000001", -- 1930 - 0x78a  :    1 - 0x1
    "00000001", -- 1931 - 0x78b  :    1 - 0x1
    "00000011", -- 1932 - 0x78c  :    3 - 0x3
    "00000111", -- 1933 - 0x78d  :    7 - 0x7
    "00000111", -- 1934 - 0x78e  :    7 - 0x7
    "00001111", -- 1935 - 0x78f  :   15 - 0xf
    "00001111", -- 1936 - 0x790  :   15 - 0xf -- Background 0x79
    "00000111", -- 1937 - 0x791  :    7 - 0x7
    "00001111", -- 1938 - 0x792  :   15 - 0xf
    "00000111", -- 1939 - 0x793  :    7 - 0x7
    "00000001", -- 1940 - 0x794  :    1 - 0x1
    "00010000", -- 1941 - 0x795  :   16 - 0x10
    "00100000", -- 1942 - 0x796  :   32 - 0x20
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- plane 1
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "00111111", -- 1946 - 0x79a  :   63 - 0x3f
    "00111111", -- 1947 - 0x79b  :   63 - 0x3f
    "01111111", -- 1948 - 0x79c  :  127 - 0x7f
    "11111110", -- 1949 - 0x79d  :  254 - 0xfe
    "11111100", -- 1950 - 0x79e  :  252 - 0xfc
    "00110000", -- 1951 - 0x79f  :   48 - 0x30
    "11111000", -- 1952 - 0x7a0  :  248 - 0xf8 -- Background 0x7a
    "11111110", -- 1953 - 0x7a1  :  254 - 0xfe
    "01111111", -- 1954 - 0x7a2  :  127 - 0x7f
    "00011111", -- 1955 - 0x7a3  :   31 - 0x1f
    "00001111", -- 1956 - 0x7a4  :   15 - 0xf
    "00011001", -- 1957 - 0x7a5  :   25 - 0x19
    "00110000", -- 1958 - 0x7a6  :   48 - 0x30
    "01110000", -- 1959 - 0x7a7  :  112 - 0x70
    "11111000", -- 1960 - 0x7a8  :  248 - 0xf8 -- plane 1
    "11111110", -- 1961 - 0x7a9  :  254 - 0xfe
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111011", -- 1968 - 0x7b0  :  251 - 0xfb -- Background 0x7b
    "01110011", -- 1969 - 0x7b1  :  115 - 0x73
    "00100111", -- 1970 - 0x7b2  :   39 - 0x27
    "00001111", -- 1971 - 0x7b3  :   15 - 0xf
    "00011111", -- 1972 - 0x7b4  :   31 - 0x1f
    "00011111", -- 1973 - 0x7b5  :   31 - 0x1f
    "00111111", -- 1974 - 0x7b6  :   63 - 0x3f
    "01111111", -- 1975 - 0x7b7  :  127 - 0x7f
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff -- plane 1
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "01111111", -- 1983 - 0x7bf  :  127 - 0x7f
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Background 0x7c
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111110", -- 1988 - 0x7c4  :  254 - 0xfe
    "11111101", -- 1989 - 0x7c5  :  253 - 0xfd
    "11111000", -- 1990 - 0x7c6  :  248 - 0xf8
    "11110110", -- 1991 - 0x7c7  :  246 - 0xf6
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- plane 1
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11101111", -- 2000 - 0x7d0  :  239 - 0xef -- Background 0x7d
    "11001111", -- 2001 - 0x7d1  :  207 - 0xcf
    "10011111", -- 2002 - 0x7d2  :  159 - 0x9f
    "00011111", -- 2003 - 0x7d3  :   31 - 0x1f
    "00001111", -- 2004 - 0x7d4  :   15 - 0xf
    "00101101", -- 2005 - 0x7d5  :   45 - 0x2d
    "01010000", -- 2006 - 0x7d6  :   80 - 0x50
    "01000000", -- 2007 - 0x7d7  :   64 - 0x40
    "11101111", -- 2008 - 0x7d8  :  239 - 0xef -- plane 1
    "11001111", -- 2009 - 0x7d9  :  207 - 0xcf
    "10011111", -- 2010 - 0x7da  :  159 - 0x9f
    "00011111", -- 2011 - 0x7db  :   31 - 0x1f
    "00001111", -- 2012 - 0x7dc  :   15 - 0xf
    "01111111", -- 2013 - 0x7dd  :  127 - 0x7f
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "11100000", -- 2020 - 0x7e4  :  224 - 0xe0
    "11111110", -- 2021 - 0x7e5  :  254 - 0xfe
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11110011", -- 2023 - 0x7e7  :  243 - 0xf3
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "11110000", -- 2027 - 0x7eb  :  240 - 0xf0
    "11111110", -- 2028 - 0x7ec  :  254 - 0xfe
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111011", -- 2032 - 0x7f0  :  251 - 0xfb -- Background 0x7f
    "11111011", -- 2033 - 0x7f1  :  251 - 0xfb
    "11111011", -- 2034 - 0x7f2  :  251 - 0xfb
    "11111011", -- 2035 - 0x7f3  :  251 - 0xfb
    "11111011", -- 2036 - 0x7f4  :  251 - 0xfb
    "11110011", -- 2037 - 0x7f5  :  243 - 0xf3
    "11110111", -- 2038 - 0x7f6  :  247 - 0xf7
    "11100111", -- 2039 - 0x7f7  :  231 - 0xe7
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- plane 1
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111", -- 2047 - 0x7ff  :  255 - 0xff
    "11001111", -- 2048 - 0x800  :  207 - 0xcf -- Background 0x80
    "10011111", -- 2049 - 0x801  :  159 - 0x9f
    "00111111", -- 2050 - 0x802  :   63 - 0x3f
    "00111111", -- 2051 - 0x803  :   63 - 0x3f
    "00111111", -- 2052 - 0x804  :   63 - 0x3f
    "00001111", -- 2053 - 0x805  :   15 - 0xf
    "00000011", -- 2054 - 0x806  :    3 - 0x3
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "11111111", -- 2056 - 0x808  :  255 - 0xff -- plane 1
    "11111111", -- 2057 - 0x809  :  255 - 0xff
    "11111111", -- 2058 - 0x80a  :  255 - 0xff
    "11111111", -- 2059 - 0x80b  :  255 - 0xff
    "11111111", -- 2060 - 0x80c  :  255 - 0xff
    "11111111", -- 2061 - 0x80d  :  255 - 0xff
    "11111111", -- 2062 - 0x80e  :  255 - 0xff
    "11111111", -- 2063 - 0x80f  :  255 - 0xff
    "11000000", -- 2064 - 0x810  :  192 - 0xc0 -- Background 0x81
    "11110000", -- 2065 - 0x811  :  240 - 0xf0
    "11111100", -- 2066 - 0x812  :  252 - 0xfc
    "11110000", -- 2067 - 0x813  :  240 - 0xf0
    "11110000", -- 2068 - 0x814  :  240 - 0xf0
    "10011000", -- 2069 - 0x815  :  152 - 0x98
    "00001000", -- 2070 - 0x816  :    8 - 0x8
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "11111111", -- 2072 - 0x818  :  255 - 0xff -- plane 1
    "11111111", -- 2073 - 0x819  :  255 - 0xff
    "11111111", -- 2074 - 0x81a  :  255 - 0xff
    "11110000", -- 2075 - 0x81b  :  240 - 0xf0
    "11110000", -- 2076 - 0x81c  :  240 - 0xf0
    "11111000", -- 2077 - 0x81d  :  248 - 0xf8
    "11111000", -- 2078 - 0x81e  :  248 - 0xf8
    "11111000", -- 2079 - 0x81f  :  248 - 0xf8
    "00000000", -- 2080 - 0x820  :    0 - 0x0 -- Background 0x82
    "00000000", -- 2081 - 0x821  :    0 - 0x0
    "00000000", -- 2082 - 0x822  :    0 - 0x0
    "00000000", -- 2083 - 0x823  :    0 - 0x0
    "00000000", -- 2084 - 0x824  :    0 - 0x0
    "00000000", -- 2085 - 0x825  :    0 - 0x0
    "10000000", -- 2086 - 0x826  :  128 - 0x80
    "11000000", -- 2087 - 0x827  :  192 - 0xc0
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- plane 1
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "00000000", -- 2092 - 0x82c  :    0 - 0x0
    "10000000", -- 2093 - 0x82d  :  128 - 0x80
    "11000000", -- 2094 - 0x82e  :  192 - 0xc0
    "11100000", -- 2095 - 0x82f  :  224 - 0xe0
    "11100000", -- 2096 - 0x830  :  224 - 0xe0 -- Background 0x83
    "11100000", -- 2097 - 0x831  :  224 - 0xe0
    "11110000", -- 2098 - 0x832  :  240 - 0xf0
    "11110000", -- 2099 - 0x833  :  240 - 0xf0
    "11110000", -- 2100 - 0x834  :  240 - 0xf0
    "11110000", -- 2101 - 0x835  :  240 - 0xf0
    "11111000", -- 2102 - 0x836  :  248 - 0xf8
    "11111000", -- 2103 - 0x837  :  248 - 0xf8
    "11110000", -- 2104 - 0x838  :  240 - 0xf0 -- plane 1
    "11110000", -- 2105 - 0x839  :  240 - 0xf0
    "11111000", -- 2106 - 0x83a  :  248 - 0xf8
    "11111000", -- 2107 - 0x83b  :  248 - 0xf8
    "11111000", -- 2108 - 0x83c  :  248 - 0xf8
    "11111100", -- 2109 - 0x83d  :  252 - 0xfc
    "11111100", -- 2110 - 0x83e  :  252 - 0xfc
    "11111110", -- 2111 - 0x83f  :  254 - 0xfe
    "11111110", -- 2112 - 0x840  :  254 - 0xfe -- Background 0x84
    "11111111", -- 2113 - 0x841  :  255 - 0xff
    "11111111", -- 2114 - 0x842  :  255 - 0xff
    "11111111", -- 2115 - 0x843  :  255 - 0xff
    "11111111", -- 2116 - 0x844  :  255 - 0xff
    "11111111", -- 2117 - 0x845  :  255 - 0xff
    "11111111", -- 2118 - 0x846  :  255 - 0xff
    "11111111", -- 2119 - 0x847  :  255 - 0xff
    "11111111", -- 2120 - 0x848  :  255 - 0xff -- plane 1
    "11111111", -- 2121 - 0x849  :  255 - 0xff
    "11111111", -- 2122 - 0x84a  :  255 - 0xff
    "11111111", -- 2123 - 0x84b  :  255 - 0xff
    "11111111", -- 2124 - 0x84c  :  255 - 0xff
    "11111111", -- 2125 - 0x84d  :  255 - 0xff
    "11111111", -- 2126 - 0x84e  :  255 - 0xff
    "11111111", -- 2127 - 0x84f  :  255 - 0xff
    "00111111", -- 2128 - 0x850  :   63 - 0x3f -- Background 0x85
    "00011111", -- 2129 - 0x851  :   31 - 0x1f
    "00011111", -- 2130 - 0x852  :   31 - 0x1f
    "00001111", -- 2131 - 0x853  :   15 - 0xf
    "00000111", -- 2132 - 0x854  :    7 - 0x7
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "11111111", -- 2136 - 0x858  :  255 - 0xff -- plane 1
    "11111111", -- 2137 - 0x859  :  255 - 0xff
    "11111111", -- 2138 - 0x85a  :  255 - 0xff
    "00001111", -- 2139 - 0x85b  :   15 - 0xf
    "00000111", -- 2140 - 0x85c  :    7 - 0x7
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Background 0x86
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "11000000", -- 2146 - 0x862  :  192 - 0xc0
    "11100000", -- 2147 - 0x863  :  224 - 0xe0
    "11110000", -- 2148 - 0x864  :  240 - 0xf0
    "11110000", -- 2149 - 0x865  :  240 - 0xf0
    "11110000", -- 2150 - 0x866  :  240 - 0xf0
    "11111000", -- 2151 - 0x867  :  248 - 0xf8
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- plane 1
    "10000000", -- 2153 - 0x869  :  128 - 0x80
    "11000000", -- 2154 - 0x86a  :  192 - 0xc0
    "11100000", -- 2155 - 0x86b  :  224 - 0xe0
    "11110000", -- 2156 - 0x86c  :  240 - 0xf0
    "11110000", -- 2157 - 0x86d  :  240 - 0xf0
    "11110000", -- 2158 - 0x86e  :  240 - 0xf0
    "11111100", -- 2159 - 0x86f  :  252 - 0xfc
    "11111001", -- 2160 - 0x870  :  249 - 0xf9 -- Background 0x87
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "00001110", -- 2165 - 0x875  :   14 - 0xe
    "00000010", -- 2166 - 0x876  :    2 - 0x2
    "00010100", -- 2167 - 0x877  :   20 - 0x14
    "11111111", -- 2168 - 0x878  :  255 - 0xff -- plane 1
    "11111111", -- 2169 - 0x879  :  255 - 0xff
    "11111111", -- 2170 - 0x87a  :  255 - 0xff
    "11111111", -- 2171 - 0x87b  :  255 - 0xff
    "11111111", -- 2172 - 0x87c  :  255 - 0xff
    "00001111", -- 2173 - 0x87d  :   15 - 0xf
    "00011111", -- 2174 - 0x87e  :   31 - 0x1f
    "00111111", -- 2175 - 0x87f  :   63 - 0x3f
    "10000000", -- 2176 - 0x880  :  128 - 0x80 -- Background 0x88
    "10100000", -- 2177 - 0x881  :  160 - 0xa0
    "00100000", -- 2178 - 0x882  :   32 - 0x20
    "00100000", -- 2179 - 0x883  :   32 - 0x20
    "10100000", -- 2180 - 0x884  :  160 - 0xa0
    "10000000", -- 2181 - 0x885  :  128 - 0x80
    "00000000", -- 2182 - 0x886  :    0 - 0x0
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "11000000", -- 2184 - 0x888  :  192 - 0xc0 -- plane 1
    "11100000", -- 2185 - 0x889  :  224 - 0xe0
    "11100000", -- 2186 - 0x88a  :  224 - 0xe0
    "11100000", -- 2187 - 0x88b  :  224 - 0xe0
    "11100000", -- 2188 - 0x88c  :  224 - 0xe0
    "11000000", -- 2189 - 0x88d  :  192 - 0xc0
    "11000000", -- 2190 - 0x88e  :  192 - 0xc0
    "10000000", -- 2191 - 0x88f  :  128 - 0x80
    "00000001", -- 2192 - 0x890  :    1 - 0x1 -- Background 0x89
    "00000101", -- 2193 - 0x891  :    5 - 0x5
    "00000100", -- 2194 - 0x892  :    4 - 0x4
    "00000100", -- 2195 - 0x893  :    4 - 0x4
    "00000101", -- 2196 - 0x894  :    5 - 0x5
    "00000001", -- 2197 - 0x895  :    1 - 0x1
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000011", -- 2200 - 0x898  :    3 - 0x3 -- plane 1
    "00000111", -- 2201 - 0x899  :    7 - 0x7
    "00000111", -- 2202 - 0x89a  :    7 - 0x7
    "00000111", -- 2203 - 0x89b  :    7 - 0x7
    "00000111", -- 2204 - 0x89c  :    7 - 0x7
    "00000011", -- 2205 - 0x89d  :    3 - 0x3
    "00000011", -- 2206 - 0x89e  :    3 - 0x3
    "00000001", -- 2207 - 0x89f  :    1 - 0x1
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000011", -- 2210 - 0x8a2  :    3 - 0x3
    "00000111", -- 2211 - 0x8a3  :    7 - 0x7
    "00001111", -- 2212 - 0x8a4  :   15 - 0xf
    "00001111", -- 2213 - 0x8a5  :   15 - 0xf
    "00001111", -- 2214 - 0x8a6  :   15 - 0xf
    "00001111", -- 2215 - 0x8a7  :   15 - 0xf
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- plane 1
    "00000001", -- 2217 - 0x8a9  :    1 - 0x1
    "00000011", -- 2218 - 0x8aa  :    3 - 0x3
    "00000111", -- 2219 - 0x8ab  :    7 - 0x7
    "00001111", -- 2220 - 0x8ac  :   15 - 0xf
    "00001111", -- 2221 - 0x8ad  :   15 - 0xf
    "00001111", -- 2222 - 0x8ae  :   15 - 0xf
    "00111111", -- 2223 - 0x8af  :   63 - 0x3f
    "10011111", -- 2224 - 0x8b0  :  159 - 0x9f -- Background 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11111111", -- 2226 - 0x8b2  :  255 - 0xff
    "11111111", -- 2227 - 0x8b3  :  255 - 0xff
    "11111111", -- 2228 - 0x8b4  :  255 - 0xff
    "01110000", -- 2229 - 0x8b5  :  112 - 0x70
    "01000000", -- 2230 - 0x8b6  :   64 - 0x40
    "00101000", -- 2231 - 0x8b7  :   40 - 0x28
    "11111111", -- 2232 - 0x8b8  :  255 - 0xff -- plane 1
    "11111111", -- 2233 - 0x8b9  :  255 - 0xff
    "11111111", -- 2234 - 0x8ba  :  255 - 0xff
    "11111111", -- 2235 - 0x8bb  :  255 - 0xff
    "11111111", -- 2236 - 0x8bc  :  255 - 0xff
    "11110000", -- 2237 - 0x8bd  :  240 - 0xf0
    "11111000", -- 2238 - 0x8be  :  248 - 0xf8
    "11111100", -- 2239 - 0x8bf  :  252 - 0xfc
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000000", -- 2244 - 0x8c4  :    0 - 0x0
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "00000001", -- 2246 - 0x8c6  :    1 - 0x1
    "00000011", -- 2247 - 0x8c7  :    3 - 0x3
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000001", -- 2253 - 0x8cd  :    1 - 0x1
    "00000011", -- 2254 - 0x8ce  :    3 - 0x3
    "00000111", -- 2255 - 0x8cf  :    7 - 0x7
    "00000111", -- 2256 - 0x8d0  :    7 - 0x7 -- Background 0x8d
    "00000111", -- 2257 - 0x8d1  :    7 - 0x7
    "00001111", -- 2258 - 0x8d2  :   15 - 0xf
    "00001111", -- 2259 - 0x8d3  :   15 - 0xf
    "00001111", -- 2260 - 0x8d4  :   15 - 0xf
    "00001111", -- 2261 - 0x8d5  :   15 - 0xf
    "00011111", -- 2262 - 0x8d6  :   31 - 0x1f
    "00011111", -- 2263 - 0x8d7  :   31 - 0x1f
    "00001111", -- 2264 - 0x8d8  :   15 - 0xf -- plane 1
    "00001111", -- 2265 - 0x8d9  :   15 - 0xf
    "00011111", -- 2266 - 0x8da  :   31 - 0x1f
    "00011111", -- 2267 - 0x8db  :   31 - 0x1f
    "00011111", -- 2268 - 0x8dc  :   31 - 0x1f
    "00111111", -- 2269 - 0x8dd  :   63 - 0x3f
    "00111111", -- 2270 - 0x8de  :   63 - 0x3f
    "01111111", -- 2271 - 0x8df  :  127 - 0x7f
    "01111111", -- 2272 - 0x8e0  :  127 - 0x7f -- Background 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11111111", -- 2274 - 0x8e2  :  255 - 0xff
    "11111111", -- 2275 - 0x8e3  :  255 - 0xff
    "11111111", -- 2276 - 0x8e4  :  255 - 0xff
    "11111111", -- 2277 - 0x8e5  :  255 - 0xff
    "11111111", -- 2278 - 0x8e6  :  255 - 0xff
    "11111111", -- 2279 - 0x8e7  :  255 - 0xff
    "11111111", -- 2280 - 0x8e8  :  255 - 0xff -- plane 1
    "11111111", -- 2281 - 0x8e9  :  255 - 0xff
    "11111111", -- 2282 - 0x8ea  :  255 - 0xff
    "11111111", -- 2283 - 0x8eb  :  255 - 0xff
    "11111111", -- 2284 - 0x8ec  :  255 - 0xff
    "11111111", -- 2285 - 0x8ed  :  255 - 0xff
    "11111111", -- 2286 - 0x8ee  :  255 - 0xff
    "11111111", -- 2287 - 0x8ef  :  255 - 0xff
    "11111100", -- 2288 - 0x8f0  :  252 - 0xfc -- Background 0x8f
    "11111000", -- 2289 - 0x8f1  :  248 - 0xf8
    "11111000", -- 2290 - 0x8f2  :  248 - 0xf8
    "11110000", -- 2291 - 0x8f3  :  240 - 0xf0
    "11100000", -- 2292 - 0x8f4  :  224 - 0xe0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "11111111", -- 2296 - 0x8f8  :  255 - 0xff -- plane 1
    "11111111", -- 2297 - 0x8f9  :  255 - 0xff
    "11111111", -- 2298 - 0x8fa  :  255 - 0xff
    "11110000", -- 2299 - 0x8fb  :  240 - 0xf0
    "11100000", -- 2300 - 0x8fc  :  224 - 0xe0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000111", -- 2308 - 0x904  :    7 - 0x7
    "01111111", -- 2309 - 0x905  :  127 - 0x7f
    "11111111", -- 2310 - 0x906  :  255 - 0xff
    "11001111", -- 2311 - 0x907  :  207 - 0xcf
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- plane 1
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00001111", -- 2315 - 0x90b  :   15 - 0xf
    "01111111", -- 2316 - 0x90c  :  127 - 0x7f
    "11111111", -- 2317 - 0x90d  :  255 - 0xff
    "11111111", -- 2318 - 0x90e  :  255 - 0xff
    "11111111", -- 2319 - 0x90f  :  255 - 0xff
    "11011111", -- 2320 - 0x910  :  223 - 0xdf -- Background 0x91
    "11011111", -- 2321 - 0x911  :  223 - 0xdf
    "11011111", -- 2322 - 0x912  :  223 - 0xdf
    "11011111", -- 2323 - 0x913  :  223 - 0xdf
    "11011111", -- 2324 - 0x914  :  223 - 0xdf
    "11001111", -- 2325 - 0x915  :  207 - 0xcf
    "11101111", -- 2326 - 0x916  :  239 - 0xef
    "11100111", -- 2327 - 0x917  :  231 - 0xe7
    "11111111", -- 2328 - 0x918  :  255 - 0xff -- plane 1
    "11111111", -- 2329 - 0x919  :  255 - 0xff
    "11111111", -- 2330 - 0x91a  :  255 - 0xff
    "11111111", -- 2331 - 0x91b  :  255 - 0xff
    "11111111", -- 2332 - 0x91c  :  255 - 0xff
    "11111111", -- 2333 - 0x91d  :  255 - 0xff
    "11111111", -- 2334 - 0x91e  :  255 - 0xff
    "11111111", -- 2335 - 0x91f  :  255 - 0xff
    "11110011", -- 2336 - 0x920  :  243 - 0xf3 -- Background 0x92
    "11111001", -- 2337 - 0x921  :  249 - 0xf9
    "11111100", -- 2338 - 0x922  :  252 - 0xfc
    "11111100", -- 2339 - 0x923  :  252 - 0xfc
    "11111100", -- 2340 - 0x924  :  252 - 0xfc
    "11110000", -- 2341 - 0x925  :  240 - 0xf0
    "11000000", -- 2342 - 0x926  :  192 - 0xc0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "11111111", -- 2344 - 0x928  :  255 - 0xff -- plane 1
    "11111111", -- 2345 - 0x929  :  255 - 0xff
    "11111111", -- 2346 - 0x92a  :  255 - 0xff
    "11111111", -- 2347 - 0x92b  :  255 - 0xff
    "11111111", -- 2348 - 0x92c  :  255 - 0xff
    "11111111", -- 2349 - 0x92d  :  255 - 0xff
    "11111111", -- 2350 - 0x92e  :  255 - 0xff
    "11111111", -- 2351 - 0x92f  :  255 - 0xff
    "00000011", -- 2352 - 0x930  :    3 - 0x3 -- Background 0x93
    "00001111", -- 2353 - 0x931  :   15 - 0xf
    "00111111", -- 2354 - 0x932  :   63 - 0x3f
    "00001111", -- 2355 - 0x933  :   15 - 0xf
    "00001111", -- 2356 - 0x934  :   15 - 0xf
    "00011001", -- 2357 - 0x935  :   25 - 0x19
    "00010000", -- 2358 - 0x936  :   16 - 0x10
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "11111111", -- 2360 - 0x938  :  255 - 0xff -- plane 1
    "11111111", -- 2361 - 0x939  :  255 - 0xff
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "00001111", -- 2363 - 0x93b  :   15 - 0xf
    "00001111", -- 2364 - 0x93c  :   15 - 0xf
    "00011111", -- 2365 - 0x93d  :   31 - 0x1f
    "00011111", -- 2366 - 0x93e  :   31 - 0x1f
    "00011111", -- 2367 - 0x93f  :   31 - 0x1f
    "00011111", -- 2368 - 0x940  :   31 - 0x1f -- Background 0x94
    "01111111", -- 2369 - 0x941  :  127 - 0x7f
    "11111110", -- 2370 - 0x942  :  254 - 0xfe
    "11111000", -- 2371 - 0x943  :  248 - 0xf8
    "11110000", -- 2372 - 0x944  :  240 - 0xf0
    "10011000", -- 2373 - 0x945  :  152 - 0x98
    "00001100", -- 2374 - 0x946  :   12 - 0xc
    "00001110", -- 2375 - 0x947  :   14 - 0xe
    "00011111", -- 2376 - 0x948  :   31 - 0x1f -- plane 1
    "01111111", -- 2377 - 0x949  :  127 - 0x7f
    "11111111", -- 2378 - 0x94a  :  255 - 0xff
    "11111111", -- 2379 - 0x94b  :  255 - 0xff
    "11111111", -- 2380 - 0x94c  :  255 - 0xff
    "11111111", -- 2381 - 0x94d  :  255 - 0xff
    "11111111", -- 2382 - 0x94e  :  255 - 0xff
    "11111111", -- 2383 - 0x94f  :  255 - 0xff
    "11011111", -- 2384 - 0x950  :  223 - 0xdf -- Background 0x95
    "11001110", -- 2385 - 0x951  :  206 - 0xce
    "11100100", -- 2386 - 0x952  :  228 - 0xe4
    "11110000", -- 2387 - 0x953  :  240 - 0xf0
    "11111000", -- 2388 - 0x954  :  248 - 0xf8
    "11111000", -- 2389 - 0x955  :  248 - 0xf8
    "11111100", -- 2390 - 0x956  :  252 - 0xfc
    "11111110", -- 2391 - 0x957  :  254 - 0xfe
    "11111111", -- 2392 - 0x958  :  255 - 0xff -- plane 1
    "11111111", -- 2393 - 0x959  :  255 - 0xff
    "11111111", -- 2394 - 0x95a  :  255 - 0xff
    "11111111", -- 2395 - 0x95b  :  255 - 0xff
    "11111111", -- 2396 - 0x95c  :  255 - 0xff
    "11111111", -- 2397 - 0x95d  :  255 - 0xff
    "11111111", -- 2398 - 0x95e  :  255 - 0xff
    "11111110", -- 2399 - 0x95f  :  254 - 0xfe
    "11111111", -- 2400 - 0x960  :  255 - 0xff -- Background 0x96
    "11111111", -- 2401 - 0x961  :  255 - 0xff
    "11111111", -- 2402 - 0x962  :  255 - 0xff
    "11111111", -- 2403 - 0x963  :  255 - 0xff
    "01111111", -- 2404 - 0x964  :  127 - 0x7f
    "10111111", -- 2405 - 0x965  :  191 - 0xbf
    "00011111", -- 2406 - 0x966  :   31 - 0x1f
    "01101111", -- 2407 - 0x967  :  111 - 0x6f
    "11111111", -- 2408 - 0x968  :  255 - 0xff -- plane 1
    "11111111", -- 2409 - 0x969  :  255 - 0xff
    "11111111", -- 2410 - 0x96a  :  255 - 0xff
    "11111111", -- 2411 - 0x96b  :  255 - 0xff
    "11111111", -- 2412 - 0x96c  :  255 - 0xff
    "11111111", -- 2413 - 0x96d  :  255 - 0xff
    "11111111", -- 2414 - 0x96e  :  255 - 0xff
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "11110111", -- 2416 - 0x970  :  247 - 0xf7 -- Background 0x97
    "11110011", -- 2417 - 0x971  :  243 - 0xf3
    "11111001", -- 2418 - 0x972  :  249 - 0xf9
    "11111000", -- 2419 - 0x973  :  248 - 0xf8
    "11110000", -- 2420 - 0x974  :  240 - 0xf0
    "10110100", -- 2421 - 0x975  :  180 - 0xb4
    "00001010", -- 2422 - 0x976  :   10 - 0xa
    "00000010", -- 2423 - 0x977  :    2 - 0x2
    "11110111", -- 2424 - 0x978  :  247 - 0xf7 -- plane 1
    "11110011", -- 2425 - 0x979  :  243 - 0xf3
    "11111001", -- 2426 - 0x97a  :  249 - 0xf9
    "11111000", -- 2427 - 0x97b  :  248 - 0xf8
    "11110000", -- 2428 - 0x97c  :  240 - 0xf0
    "11111110", -- 2429 - 0x97d  :  254 - 0xfe
    "11111111", -- 2430 - 0x97e  :  255 - 0xff
    "11111111", -- 2431 - 0x97f  :  255 - 0xff
    "10000000", -- 2432 - 0x980  :  128 - 0x80 -- Background 0x98
    "11000000", -- 2433 - 0x981  :  192 - 0xc0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "11000000", -- 2436 - 0x984  :  192 - 0xc0
    "10011000", -- 2437 - 0x985  :  152 - 0x98
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "10000000", -- 2440 - 0x988  :  128 - 0x80 -- plane 1
    "11000000", -- 2441 - 0x989  :  192 - 0xc0
    "11000000", -- 2442 - 0x98a  :  192 - 0xc0
    "11100000", -- 2443 - 0x98b  :  224 - 0xe0
    "00100000", -- 2444 - 0x98c  :   32 - 0x20
    "00111000", -- 2445 - 0x98d  :   56 - 0x38
    "11111100", -- 2446 - 0x98e  :  252 - 0xfc
    "11111110", -- 2447 - 0x98f  :  254 - 0xfe
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Background 0x99
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00111110", -- 2450 - 0x992  :   62 - 0x3e
    "01000000", -- 2451 - 0x993  :   64 - 0x40
    "10000000", -- 2452 - 0x994  :  128 - 0x80
    "00000000", -- 2453 - 0x995  :    0 - 0x0
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "11111110", -- 2456 - 0x998  :  254 - 0xfe -- plane 1
    "11111111", -- 2457 - 0x999  :  255 - 0xff
    "11111111", -- 2458 - 0x99a  :  255 - 0xff
    "11111110", -- 2459 - 0x99b  :  254 - 0xfe
    "11111100", -- 2460 - 0x99c  :  252 - 0xfc
    "11111000", -- 2461 - 0x99d  :  248 - 0xf8
    "11000000", -- 2462 - 0x99e  :  192 - 0xc0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "10000000", -- 2466 - 0x9a2  :  128 - 0x80
    "10000000", -- 2467 - 0x9a3  :  128 - 0x80
    "11000000", -- 2468 - 0x9a4  :  192 - 0xc0
    "11100000", -- 2469 - 0x9a5  :  224 - 0xe0
    "11100000", -- 2470 - 0x9a6  :  224 - 0xe0
    "11110000", -- 2471 - 0x9a7  :  240 - 0xf0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "10000000", -- 2474 - 0x9aa  :  128 - 0x80
    "10000000", -- 2475 - 0x9ab  :  128 - 0x80
    "11000000", -- 2476 - 0x9ac  :  192 - 0xc0
    "11100000", -- 2477 - 0x9ad  :  224 - 0xe0
    "11100000", -- 2478 - 0x9ae  :  224 - 0xe0
    "11110000", -- 2479 - 0x9af  :  240 - 0xf0
    "11110000", -- 2480 - 0x9b0  :  240 - 0xf0 -- Background 0x9b
    "11100000", -- 2481 - 0x9b1  :  224 - 0xe0
    "11110000", -- 2482 - 0x9b2  :  240 - 0xf0
    "11100000", -- 2483 - 0x9b3  :  224 - 0xe0
    "10000000", -- 2484 - 0x9b4  :  128 - 0x80
    "00001000", -- 2485 - 0x9b5  :    8 - 0x8
    "00000100", -- 2486 - 0x9b6  :    4 - 0x4
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "11111111", -- 2488 - 0x9b8  :  255 - 0xff -- plane 1
    "11111111", -- 2489 - 0x9b9  :  255 - 0xff
    "11111100", -- 2490 - 0x9ba  :  252 - 0xfc
    "11111100", -- 2491 - 0x9bb  :  252 - 0xfc
    "11111110", -- 2492 - 0x9bc  :  254 - 0xfe
    "01111110", -- 2493 - 0x9bd  :  126 - 0x7e
    "00111111", -- 2494 - 0x9be  :   63 - 0x3f
    "00001100", -- 2495 - 0x9bf  :   12 - 0xc
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000001", -- 2498 - 0x9c2  :    1 - 0x1
    "00000011", -- 2499 - 0x9c3  :    3 - 0x3
    "00000011", -- 2500 - 0x9c4  :    3 - 0x3
    "00000011", -- 2501 - 0x9c5  :    3 - 0x3
    "00000111", -- 2502 - 0x9c6  :    7 - 0x7
    "00000111", -- 2503 - 0x9c7  :    7 - 0x7
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- plane 1
    "00000001", -- 2505 - 0x9c9  :    1 - 0x1
    "00000011", -- 2506 - 0x9ca  :    3 - 0x3
    "00000111", -- 2507 - 0x9cb  :    7 - 0x7
    "00000111", -- 2508 - 0x9cc  :    7 - 0x7
    "00000111", -- 2509 - 0x9cd  :    7 - 0x7
    "00001111", -- 2510 - 0x9ce  :   15 - 0xf
    "00001111", -- 2511 - 0x9cf  :   15 - 0xf
    "00000111", -- 2512 - 0x9d0  :    7 - 0x7 -- Background 0x9d
    "00000011", -- 2513 - 0x9d1  :    3 - 0x3
    "00000011", -- 2514 - 0x9d2  :    3 - 0x3
    "00000011", -- 2515 - 0x9d3  :    3 - 0x3
    "00000011", -- 2516 - 0x9d4  :    3 - 0x3
    "00000011", -- 2517 - 0x9d5  :    3 - 0x3
    "00000011", -- 2518 - 0x9d6  :    3 - 0x3
    "00000001", -- 2519 - 0x9d7  :    1 - 0x1
    "00001111", -- 2520 - 0x9d8  :   15 - 0xf -- plane 1
    "00001111", -- 2521 - 0x9d9  :   15 - 0xf
    "00000111", -- 2522 - 0x9da  :    7 - 0x7
    "00000111", -- 2523 - 0x9db  :    7 - 0x7
    "00000111", -- 2524 - 0x9dc  :    7 - 0x7
    "00000011", -- 2525 - 0x9dd  :    3 - 0x3
    "00000011", -- 2526 - 0x9de  :    3 - 0x3
    "00000001", -- 2527 - 0x9df  :    1 - 0x1
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x9e
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000001", -- 2533 - 0x9e5  :    1 - 0x1
    "00000010", -- 2534 - 0x9e6  :    2 - 0x2
    "00000100", -- 2535 - 0x9e7  :    4 - 0x4
    "00000001", -- 2536 - 0x9e8  :    1 - 0x1 -- plane 1
    "00000001", -- 2537 - 0x9e9  :    1 - 0x1
    "00000001", -- 2538 - 0x9ea  :    1 - 0x1
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000011", -- 2541 - 0x9ed  :    3 - 0x3
    "00000111", -- 2542 - 0x9ee  :    7 - 0x7
    "00001111", -- 2543 - 0x9ef  :   15 - 0xf
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00011100", -- 2550 - 0x9f6  :   28 - 0x1c
    "00111011", -- 2551 - 0x9f7  :   59 - 0x3b
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- plane 1
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000001", -- 2556 - 0x9fc  :    1 - 0x1
    "00000011", -- 2557 - 0x9fd  :    3 - 0x3
    "00111111", -- 2558 - 0x9fe  :   63 - 0x3f
    "01111111", -- 2559 - 0x9ff  :  127 - 0x7f
    "01111110", -- 2560 - 0xa00  :  126 - 0x7e -- Background 0xa0
    "11111110", -- 2561 - 0xa01  :  254 - 0xfe
    "11111111", -- 2562 - 0xa02  :  255 - 0xff
    "11111111", -- 2563 - 0xa03  :  255 - 0xff
    "11111111", -- 2564 - 0xa04  :  255 - 0xff
    "11111111", -- 2565 - 0xa05  :  255 - 0xff
    "11111101", -- 2566 - 0xa06  :  253 - 0xfd
    "11111001", -- 2567 - 0xa07  :  249 - 0xf9
    "11111111", -- 2568 - 0xa08  :  255 - 0xff -- plane 1
    "11111111", -- 2569 - 0xa09  :  255 - 0xff
    "11111111", -- 2570 - 0xa0a  :  255 - 0xff
    "11111111", -- 2571 - 0xa0b  :  255 - 0xff
    "11111111", -- 2572 - 0xa0c  :  255 - 0xff
    "11111111", -- 2573 - 0xa0d  :  255 - 0xff
    "11111101", -- 2574 - 0xa0e  :  253 - 0xfd
    "11111001", -- 2575 - 0xa0f  :  249 - 0xf9
    "11110011", -- 2576 - 0xa10  :  243 - 0xf3 -- Background 0xa1
    "11110111", -- 2577 - 0xa11  :  247 - 0xf7
    "11110110", -- 2578 - 0xa12  :  246 - 0xf6
    "11101110", -- 2579 - 0xa13  :  238 - 0xee
    "11111101", -- 2580 - 0xa14  :  253 - 0xfd
    "11111100", -- 2581 - 0xa15  :  252 - 0xfc
    "11111000", -- 2582 - 0xa16  :  248 - 0xf8
    "11100001", -- 2583 - 0xa17  :  225 - 0xe1
    "11110011", -- 2584 - 0xa18  :  243 - 0xf3 -- plane 1
    "11111111", -- 2585 - 0xa19  :  255 - 0xff
    "11111111", -- 2586 - 0xa1a  :  255 - 0xff
    "11111111", -- 2587 - 0xa1b  :  255 - 0xff
    "11111111", -- 2588 - 0xa1c  :  255 - 0xff
    "11111111", -- 2589 - 0xa1d  :  255 - 0xff
    "11111111", -- 2590 - 0xa1e  :  255 - 0xff
    "11111111", -- 2591 - 0xa1f  :  255 - 0xff
    "11010011", -- 2592 - 0xa20  :  211 - 0xd3 -- Background 0xa2
    "11001011", -- 2593 - 0xa21  :  203 - 0xcb
    "11000011", -- 2594 - 0xa22  :  195 - 0xc3
    "11100001", -- 2595 - 0xa23  :  225 - 0xe1
    "11111001", -- 2596 - 0xa24  :  249 - 0xf9
    "00111001", -- 2597 - 0xa25  :   57 - 0x39
    "01000010", -- 2598 - 0xa26  :   66 - 0x42
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "11111111", -- 2600 - 0xa28  :  255 - 0xff -- plane 1
    "11111111", -- 2601 - 0xa29  :  255 - 0xff
    "11111111", -- 2602 - 0xa2a  :  255 - 0xff
    "11111111", -- 2603 - 0xa2b  :  255 - 0xff
    "11111111", -- 2604 - 0xa2c  :  255 - 0xff
    "11111111", -- 2605 - 0xa2d  :  255 - 0xff
    "11111111", -- 2606 - 0xa2e  :  255 - 0xff
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "00000111", -- 2608 - 0xa30  :    7 - 0x7 -- Background 0xa3
    "00001111", -- 2609 - 0xa31  :   15 - 0xf
    "00011001", -- 2610 - 0xa32  :   25 - 0x19
    "00110000", -- 2611 - 0xa33  :   48 - 0x30
    "01100011", -- 2612 - 0xa34  :   99 - 0x63
    "01110010", -- 2613 - 0xa35  :  114 - 0x72
    "01110000", -- 2614 - 0xa36  :  112 - 0x70
    "00000001", -- 2615 - 0xa37  :    1 - 0x1
    "00000111", -- 2616 - 0xa38  :    7 - 0x7 -- plane 1
    "00001111", -- 2617 - 0xa39  :   15 - 0xf
    "00011111", -- 2618 - 0xa3a  :   31 - 0x1f
    "00111111", -- 2619 - 0xa3b  :   63 - 0x3f
    "11111100", -- 2620 - 0xa3c  :  252 - 0xfc
    "11111100", -- 2621 - 0xa3d  :  252 - 0xfc
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0xa4
    "00011111", -- 2625 - 0xa41  :   31 - 0x1f
    "00100000", -- 2626 - 0xa42  :   32 - 0x20
    "11000000", -- 2627 - 0xa43  :  192 - 0xc0
    "11000000", -- 2628 - 0xa44  :  192 - 0xc0
    "11110000", -- 2629 - 0xa45  :  240 - 0xf0
    "11111111", -- 2630 - 0xa46  :  255 - 0xff
    "11111111", -- 2631 - 0xa47  :  255 - 0xff
    "11111111", -- 2632 - 0xa48  :  255 - 0xff -- plane 1
    "11111111", -- 2633 - 0xa49  :  255 - 0xff
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11111111", -- 2635 - 0xa4b  :  255 - 0xff
    "11111111", -- 2636 - 0xa4c  :  255 - 0xff
    "11111111", -- 2637 - 0xa4d  :  255 - 0xff
    "11111111", -- 2638 - 0xa4e  :  255 - 0xff
    "11111111", -- 2639 - 0xa4f  :  255 - 0xff
    "10101011", -- 2640 - 0xa50  :  171 - 0xab -- Background 0xa5
    "11000001", -- 2641 - 0xa51  :  193 - 0xc1
    "10000001", -- 2642 - 0xa52  :  129 - 0x81
    "10010001", -- 2643 - 0xa53  :  145 - 0x91
    "10000010", -- 2644 - 0xa54  :  130 - 0x82
    "11111100", -- 2645 - 0xa55  :  252 - 0xfc
    "11100000", -- 2646 - 0xa56  :  224 - 0xe0
    "11001110", -- 2647 - 0xa57  :  206 - 0xce
    "11111111", -- 2648 - 0xa58  :  255 - 0xff -- plane 1
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "11111111", -- 2652 - 0xa5c  :  255 - 0xff
    "11111111", -- 2653 - 0xa5d  :  255 - 0xff
    "11111111", -- 2654 - 0xa5e  :  255 - 0xff
    "11111111", -- 2655 - 0xa5f  :  255 - 0xff
    "11100101", -- 2656 - 0xa60  :  229 - 0xe5 -- Background 0xa6
    "11011010", -- 2657 - 0xa61  :  218 - 0xda
    "11110000", -- 2658 - 0xa62  :  240 - 0xf0
    "11100000", -- 2659 - 0xa63  :  224 - 0xe0
    "11000000", -- 2660 - 0xa64  :  192 - 0xc0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "11111111", -- 2664 - 0xa68  :  255 - 0xff -- plane 1
    "11111111", -- 2665 - 0xa69  :  255 - 0xff
    "11110000", -- 2666 - 0xa6a  :  240 - 0xf0
    "11100000", -- 2667 - 0xa6b  :  224 - 0xe0
    "11000000", -- 2668 - 0xa6c  :  192 - 0xc0
    "10000000", -- 2669 - 0xa6d  :  128 - 0x80
    "10000000", -- 2670 - 0xa6e  :  128 - 0x80
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "11110000", -- 2672 - 0xa70  :  240 - 0xf0 -- Background 0xa7
    "11111000", -- 2673 - 0xa71  :  248 - 0xf8
    "11001100", -- 2674 - 0xa72  :  204 - 0xcc
    "10000110", -- 2675 - 0xa73  :  134 - 0x86
    "01100010", -- 2676 - 0xa74  :   98 - 0x62
    "00100110", -- 2677 - 0xa75  :   38 - 0x26
    "00000110", -- 2678 - 0xa76  :    6 - 0x6
    "11000000", -- 2679 - 0xa77  :  192 - 0xc0
    "11110000", -- 2680 - 0xa78  :  240 - 0xf0 -- plane 1
    "11111000", -- 2681 - 0xa79  :  248 - 0xf8
    "11111100", -- 2682 - 0xa7a  :  252 - 0xfc
    "11111110", -- 2683 - 0xa7b  :  254 - 0xfe
    "10011111", -- 2684 - 0xa7c  :  159 - 0x9f
    "10011111", -- 2685 - 0xa7d  :  159 - 0x9f
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Background 0xa8
    "11111100", -- 2689 - 0xa81  :  252 - 0xfc
    "00000110", -- 2690 - 0xa82  :    6 - 0x6
    "00000011", -- 2691 - 0xa83  :    3 - 0x3
    "00000001", -- 2692 - 0xa84  :    1 - 0x1
    "00000111", -- 2693 - 0xa85  :    7 - 0x7
    "11111111", -- 2694 - 0xa86  :  255 - 0xff
    "11111111", -- 2695 - 0xa87  :  255 - 0xff
    "11111111", -- 2696 - 0xa88  :  255 - 0xff -- plane 1
    "11111111", -- 2697 - 0xa89  :  255 - 0xff
    "11111111", -- 2698 - 0xa8a  :  255 - 0xff
    "11111111", -- 2699 - 0xa8b  :  255 - 0xff
    "11111111", -- 2700 - 0xa8c  :  255 - 0xff
    "11111111", -- 2701 - 0xa8d  :  255 - 0xff
    "11111111", -- 2702 - 0xa8e  :  255 - 0xff
    "11111111", -- 2703 - 0xa8f  :  255 - 0xff
    "11010101", -- 2704 - 0xa90  :  213 - 0xd5 -- Background 0xa9
    "10000011", -- 2705 - 0xa91  :  131 - 0x83
    "10000001", -- 2706 - 0xa92  :  129 - 0x81
    "10001001", -- 2707 - 0xa93  :  137 - 0x89
    "01000001", -- 2708 - 0xa94  :   65 - 0x41
    "00111111", -- 2709 - 0xa95  :   63 - 0x3f
    "00000111", -- 2710 - 0xa96  :    7 - 0x7
    "11010011", -- 2711 - 0xa97  :  211 - 0xd3
    "11111111", -- 2712 - 0xa98  :  255 - 0xff -- plane 1
    "11111111", -- 2713 - 0xa99  :  255 - 0xff
    "11111111", -- 2714 - 0xa9a  :  255 - 0xff
    "11111111", -- 2715 - 0xa9b  :  255 - 0xff
    "11111111", -- 2716 - 0xa9c  :  255 - 0xff
    "11111111", -- 2717 - 0xa9d  :  255 - 0xff
    "11111111", -- 2718 - 0xa9e  :  255 - 0xff
    "11111111", -- 2719 - 0xa9f  :  255 - 0xff
    "01101111", -- 2720 - 0xaa0  :  111 - 0x6f -- Background 0xaa
    "11011011", -- 2721 - 0xaa1  :  219 - 0xdb
    "00001111", -- 2722 - 0xaa2  :   15 - 0xf
    "00000111", -- 2723 - 0xaa3  :    7 - 0x7
    "00000011", -- 2724 - 0xaa4  :    3 - 0x3
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "11111111", -- 2728 - 0xaa8  :  255 - 0xff -- plane 1
    "11111111", -- 2729 - 0xaa9  :  255 - 0xff
    "00001111", -- 2730 - 0xaaa  :   15 - 0xf
    "00000111", -- 2731 - 0xaab  :    7 - 0x7
    "00000011", -- 2732 - 0xaac  :    3 - 0x3
    "00000001", -- 2733 - 0xaad  :    1 - 0x1
    "00000001", -- 2734 - 0xaae  :    1 - 0x1
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "00000000", -- 2736 - 0xab0  :    0 - 0x0 -- Background 0xab
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00111000", -- 2742 - 0xab6  :   56 - 0x38
    "11011100", -- 2743 - 0xab7  :  220 - 0xdc
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- plane 1
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "10000000", -- 2748 - 0xabc  :  128 - 0x80
    "11000000", -- 2749 - 0xabd  :  192 - 0xc0
    "11111100", -- 2750 - 0xabe  :  252 - 0xfc
    "11111110", -- 2751 - 0xabf  :  254 - 0xfe
    "01111110", -- 2752 - 0xac0  :  126 - 0x7e -- Background 0xac
    "01111111", -- 2753 - 0xac1  :  127 - 0x7f
    "01111111", -- 2754 - 0xac2  :  127 - 0x7f
    "11111111", -- 2755 - 0xac3  :  255 - 0xff
    "11111111", -- 2756 - 0xac4  :  255 - 0xff
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "10111111", -- 2758 - 0xac6  :  191 - 0xbf
    "10011111", -- 2759 - 0xac7  :  159 - 0x9f
    "11111111", -- 2760 - 0xac8  :  255 - 0xff -- plane 1
    "11111111", -- 2761 - 0xac9  :  255 - 0xff
    "11111111", -- 2762 - 0xaca  :  255 - 0xff
    "11111111", -- 2763 - 0xacb  :  255 - 0xff
    "11111111", -- 2764 - 0xacc  :  255 - 0xff
    "11111111", -- 2765 - 0xacd  :  255 - 0xff
    "10111111", -- 2766 - 0xace  :  191 - 0xbf
    "10011111", -- 2767 - 0xacf  :  159 - 0x9f
    "11001111", -- 2768 - 0xad0  :  207 - 0xcf -- Background 0xad
    "11101111", -- 2769 - 0xad1  :  239 - 0xef
    "01101111", -- 2770 - 0xad2  :  111 - 0x6f
    "01110111", -- 2771 - 0xad3  :  119 - 0x77
    "10111111", -- 2772 - 0xad4  :  191 - 0xbf
    "00111111", -- 2773 - 0xad5  :   63 - 0x3f
    "00011111", -- 2774 - 0xad6  :   31 - 0x1f
    "10000111", -- 2775 - 0xad7  :  135 - 0x87
    "11001111", -- 2776 - 0xad8  :  207 - 0xcf -- plane 1
    "11111111", -- 2777 - 0xad9  :  255 - 0xff
    "11111111", -- 2778 - 0xada  :  255 - 0xff
    "11111111", -- 2779 - 0xadb  :  255 - 0xff
    "11111111", -- 2780 - 0xadc  :  255 - 0xff
    "11111111", -- 2781 - 0xadd  :  255 - 0xff
    "11111111", -- 2782 - 0xade  :  255 - 0xff
    "11111111", -- 2783 - 0xadf  :  255 - 0xff
    "11001011", -- 2784 - 0xae0  :  203 - 0xcb -- Background 0xae
    "11010011", -- 2785 - 0xae1  :  211 - 0xd3
    "11000011", -- 2786 - 0xae2  :  195 - 0xc3
    "10000111", -- 2787 - 0xae3  :  135 - 0x87
    "10011111", -- 2788 - 0xae4  :  159 - 0x9f
    "10011100", -- 2789 - 0xae5  :  156 - 0x9c
    "01000010", -- 2790 - 0xae6  :   66 - 0x42
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "11111111", -- 2792 - 0xae8  :  255 - 0xff -- plane 1
    "11111111", -- 2793 - 0xae9  :  255 - 0xff
    "11111111", -- 2794 - 0xaea  :  255 - 0xff
    "11111111", -- 2795 - 0xaeb  :  255 - 0xff
    "11111111", -- 2796 - 0xaec  :  255 - 0xff
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "11111111", -- 2798 - 0xaee  :  255 - 0xff
    "11111111", -- 2799 - 0xaef  :  255 - 0xff
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "10000000", -- 2802 - 0xaf2  :  128 - 0x80
    "11000000", -- 2803 - 0xaf3  :  192 - 0xc0
    "11000000", -- 2804 - 0xaf4  :  192 - 0xc0
    "11000000", -- 2805 - 0xaf5  :  192 - 0xc0
    "11100000", -- 2806 - 0xaf6  :  224 - 0xe0
    "11100000", -- 2807 - 0xaf7  :  224 - 0xe0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- plane 1
    "10000000", -- 2809 - 0xaf9  :  128 - 0x80
    "11000000", -- 2810 - 0xafa  :  192 - 0xc0
    "11100000", -- 2811 - 0xafb  :  224 - 0xe0
    "11100000", -- 2812 - 0xafc  :  224 - 0xe0
    "11100000", -- 2813 - 0xafd  :  224 - 0xe0
    "11110000", -- 2814 - 0xafe  :  240 - 0xf0
    "11110000", -- 2815 - 0xaff  :  240 - 0xf0
    "11100000", -- 2816 - 0xb00  :  224 - 0xe0 -- Background 0xb0
    "11000000", -- 2817 - 0xb01  :  192 - 0xc0
    "11000000", -- 2818 - 0xb02  :  192 - 0xc0
    "11000000", -- 2819 - 0xb03  :  192 - 0xc0
    "11000000", -- 2820 - 0xb04  :  192 - 0xc0
    "11000000", -- 2821 - 0xb05  :  192 - 0xc0
    "11000000", -- 2822 - 0xb06  :  192 - 0xc0
    "10000000", -- 2823 - 0xb07  :  128 - 0x80
    "11110000", -- 2824 - 0xb08  :  240 - 0xf0 -- plane 1
    "11110000", -- 2825 - 0xb09  :  240 - 0xf0
    "11100000", -- 2826 - 0xb0a  :  224 - 0xe0
    "11100000", -- 2827 - 0xb0b  :  224 - 0xe0
    "11100000", -- 2828 - 0xb0c  :  224 - 0xe0
    "11000000", -- 2829 - 0xb0d  :  192 - 0xc0
    "11000000", -- 2830 - 0xb0e  :  192 - 0xc0
    "10000000", -- 2831 - 0xb0f  :  128 - 0x80
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 2833 - 0xb11  :    0 - 0x0
    "00000000", -- 2834 - 0xb12  :    0 - 0x0
    "00000000", -- 2835 - 0xb13  :    0 - 0x0
    "00000000", -- 2836 - 0xb14  :    0 - 0x0
    "10000000", -- 2837 - 0xb15  :  128 - 0x80
    "01000000", -- 2838 - 0xb16  :   64 - 0x40
    "00100000", -- 2839 - 0xb17  :   32 - 0x20
    "10000000", -- 2840 - 0xb18  :  128 - 0x80 -- plane 1
    "10000000", -- 2841 - 0xb19  :  128 - 0x80
    "10000000", -- 2842 - 0xb1a  :  128 - 0x80
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "11000000", -- 2845 - 0xb1d  :  192 - 0xc0
    "11100000", -- 2846 - 0xb1e  :  224 - 0xe0
    "11110000", -- 2847 - 0xb1f  :  240 - 0xf0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000001", -- 2851 - 0xb23  :    1 - 0x1
    "00000011", -- 2852 - 0xb24  :    3 - 0x3
    "00000111", -- 2853 - 0xb25  :    7 - 0x7
    "00000111", -- 2854 - 0xb26  :    7 - 0x7
    "00000111", -- 2855 - 0xb27  :    7 - 0x7
    "00000000", -- 2856 - 0xb28  :    0 - 0x0 -- plane 1
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000001", -- 2858 - 0xb2a  :    1 - 0x1
    "00000011", -- 2859 - 0xb2b  :    3 - 0x3
    "00000111", -- 2860 - 0xb2c  :    7 - 0x7
    "00000111", -- 2861 - 0xb2d  :    7 - 0x7
    "00000111", -- 2862 - 0xb2e  :    7 - 0x7
    "00000111", -- 2863 - 0xb2f  :    7 - 0x7
    "00000011", -- 2864 - 0xb30  :    3 - 0x3 -- Background 0xb3
    "00000001", -- 2865 - 0xb31  :    1 - 0x1
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "00000000", -- 2867 - 0xb33  :    0 - 0x0
    "00000000", -- 2868 - 0xb34  :    0 - 0x0
    "00000000", -- 2869 - 0xb35  :    0 - 0x0
    "00000001", -- 2870 - 0xb36  :    1 - 0x1
    "00000001", -- 2871 - 0xb37  :    1 - 0x1
    "00000011", -- 2872 - 0xb38  :    3 - 0x3 -- plane 1
    "00000001", -- 2873 - 0xb39  :    1 - 0x1
    "00000000", -- 2874 - 0xb3a  :    0 - 0x0
    "00000000", -- 2875 - 0xb3b  :    0 - 0x0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000001", -- 2877 - 0xb3d  :    1 - 0x1
    "00000011", -- 2878 - 0xb3e  :    3 - 0x3
    "00000011", -- 2879 - 0xb3f  :    3 - 0x3
    "00000001", -- 2880 - 0xb40  :    1 - 0x1 -- Background 0xb4
    "00000001", -- 2881 - 0xb41  :    1 - 0x1
    "00000111", -- 2882 - 0xb42  :    7 - 0x7
    "00000011", -- 2883 - 0xb43  :    3 - 0x3
    "00000100", -- 2884 - 0xb44  :    4 - 0x4
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000011", -- 2888 - 0xb48  :    3 - 0x3 -- plane 1
    "00000011", -- 2889 - 0xb49  :    3 - 0x3
    "00000111", -- 2890 - 0xb4a  :    7 - 0x7
    "00011111", -- 2891 - 0xb4b  :   31 - 0x1f
    "00111111", -- 2892 - 0xb4c  :   63 - 0x3f
    "00111111", -- 2893 - 0xb4d  :   63 - 0x3f
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000111", -- 2903 - 0xb57  :    7 - 0x7
    "00000000", -- 2904 - 0xb58  :    0 - 0x0 -- plane 1
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "00000000", -- 2906 - 0xb5a  :    0 - 0x0
    "00000000", -- 2907 - 0xb5b  :    0 - 0x0
    "00000001", -- 2908 - 0xb5c  :    1 - 0x1
    "00000011", -- 2909 - 0xb5d  :    3 - 0x3
    "00000011", -- 2910 - 0xb5e  :    3 - 0x3
    "00001111", -- 2911 - 0xb5f  :   15 - 0xf
    "00001110", -- 2912 - 0xb60  :   14 - 0xe -- Background 0xb6
    "00111110", -- 2913 - 0xb61  :   62 - 0x3e
    "01111111", -- 2914 - 0xb62  :  127 - 0x7f
    "11111111", -- 2915 - 0xb63  :  255 - 0xff
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11101111", -- 2917 - 0xb65  :  239 - 0xef
    "11110111", -- 2918 - 0xb66  :  247 - 0xf7
    "11111000", -- 2919 - 0xb67  :  248 - 0xf8
    "00111111", -- 2920 - 0xb68  :   63 - 0x3f -- plane 1
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "11111111", -- 2922 - 0xb6a  :  255 - 0xff
    "11111111", -- 2923 - 0xb6b  :  255 - 0xff
    "11111111", -- 2924 - 0xb6c  :  255 - 0xff
    "11111111", -- 2925 - 0xb6d  :  255 - 0xff
    "11111111", -- 2926 - 0xb6e  :  255 - 0xff
    "11111111", -- 2927 - 0xb6f  :  255 - 0xff
    "11111111", -- 2928 - 0xb70  :  255 - 0xff -- Background 0xb7
    "11111111", -- 2929 - 0xb71  :  255 - 0xff
    "11111111", -- 2930 - 0xb72  :  255 - 0xff
    "00011111", -- 2931 - 0xb73  :   31 - 0x1f
    "00011111", -- 2932 - 0xb74  :   31 - 0x1f
    "01111111", -- 2933 - 0xb75  :  127 - 0x7f
    "11111111", -- 2934 - 0xb76  :  255 - 0xff
    "11111110", -- 2935 - 0xb77  :  254 - 0xfe
    "11111111", -- 2936 - 0xb78  :  255 - 0xff -- plane 1
    "11111111", -- 2937 - 0xb79  :  255 - 0xff
    "11111111", -- 2938 - 0xb7a  :  255 - 0xff
    "00011111", -- 2939 - 0xb7b  :   31 - 0x1f
    "01111111", -- 2940 - 0xb7c  :  127 - 0x7f
    "11111111", -- 2941 - 0xb7d  :  255 - 0xff
    "11111111", -- 2942 - 0xb7e  :  255 - 0xff
    "11111111", -- 2943 - 0xb7f  :  255 - 0xff
    "11111111", -- 2944 - 0xb80  :  255 - 0xff -- Background 0xb8
    "11111111", -- 2945 - 0xb81  :  255 - 0xff
    "11111111", -- 2946 - 0xb82  :  255 - 0xff
    "11111100", -- 2947 - 0xb83  :  252 - 0xfc
    "11111000", -- 2948 - 0xb84  :  248 - 0xf8
    "10000000", -- 2949 - 0xb85  :  128 - 0x80
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "11111111", -- 2952 - 0xb88  :  255 - 0xff -- plane 1
    "11111111", -- 2953 - 0xb89  :  255 - 0xff
    "11111111", -- 2954 - 0xb8a  :  255 - 0xff
    "11111100", -- 2955 - 0xb8b  :  252 - 0xfc
    "11111000", -- 2956 - 0xb8c  :  248 - 0xf8
    "11111000", -- 2957 - 0xb8d  :  248 - 0xf8
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00110000", -- 2960 - 0xb90  :   48 - 0x30 -- Background 0xb9
    "01111111", -- 2961 - 0xb91  :  127 - 0x7f
    "01111111", -- 2962 - 0xb92  :  127 - 0x7f
    "00111111", -- 2963 - 0xb93  :   63 - 0x3f
    "10000111", -- 2964 - 0xb94  :  135 - 0x87
    "11110000", -- 2965 - 0xb95  :  240 - 0xf0
    "11111111", -- 2966 - 0xb96  :  255 - 0xff
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "11001111", -- 2968 - 0xb98  :  207 - 0xcf -- plane 1
    "10001000", -- 2969 - 0xb99  :  136 - 0x88
    "11011101", -- 2970 - 0xb9a  :  221 - 0xdd
    "11001000", -- 2971 - 0xb9b  :  200 - 0xc8
    "11111000", -- 2972 - 0xb9c  :  248 - 0xf8
    "11111111", -- 2973 - 0xb9d  :  255 - 0xff
    "11111111", -- 2974 - 0xb9e  :  255 - 0xff
    "11111111", -- 2975 - 0xb9f  :  255 - 0xff
    "11100101", -- 2976 - 0xba0  :  229 - 0xe5 -- Background 0xba
    "11011010", -- 2977 - 0xba1  :  218 - 0xda
    "11000000", -- 2978 - 0xba2  :  192 - 0xc0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00000000", -- 2980 - 0xba4  :    0 - 0x0
    "00000000", -- 2981 - 0xba5  :    0 - 0x0
    "00000000", -- 2982 - 0xba6  :    0 - 0x0
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "11111111", -- 2984 - 0xba8  :  255 - 0xff -- plane 1
    "11111111", -- 2985 - 0xba9  :  255 - 0xff
    "11000000", -- 2986 - 0xbaa  :  192 - 0xc0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000110", -- 2992 - 0xbb0  :    6 - 0x6 -- Background 0xbb
    "11111111", -- 2993 - 0xbb1  :  255 - 0xff
    "11111111", -- 2994 - 0xbb2  :  255 - 0xff
    "11111110", -- 2995 - 0xbb3  :  254 - 0xfe
    "11110001", -- 2996 - 0xbb4  :  241 - 0xf1
    "00000111", -- 2997 - 0xbb5  :    7 - 0x7
    "11111111", -- 2998 - 0xbb6  :  255 - 0xff
    "11111111", -- 2999 - 0xbb7  :  255 - 0xff
    "11111001", -- 3000 - 0xbb8  :  249 - 0xf9 -- plane 1
    "10001000", -- 3001 - 0xbb9  :  136 - 0x88
    "11011101", -- 3002 - 0xbba  :  221 - 0xdd
    "10001001", -- 3003 - 0xbbb  :  137 - 0x89
    "00001111", -- 3004 - 0xbbc  :   15 - 0xf
    "11111111", -- 3005 - 0xbbd  :  255 - 0xff
    "11111111", -- 3006 - 0xbbe  :  255 - 0xff
    "11111111", -- 3007 - 0xbbf  :  255 - 0xff
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0xbc
    "00000001", -- 3009 - 0xbc1  :    1 - 0x1
    "00000010", -- 3010 - 0xbc2  :    2 - 0x2
    "00000111", -- 3011 - 0xbc3  :    7 - 0x7
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00100000", -- 3014 - 0xbc6  :   32 - 0x20
    "11111111", -- 3015 - 0xbc7  :  255 - 0xff
    "00000011", -- 3016 - 0xbc8  :    3 - 0x3 -- plane 1
    "00000111", -- 3017 - 0xbc9  :    7 - 0x7
    "00001111", -- 3018 - 0xbca  :   15 - 0xf
    "00000111", -- 3019 - 0xbcb  :    7 - 0x7
    "10000111", -- 3020 - 0xbcc  :  135 - 0x87
    "11000011", -- 3021 - 0xbcd  :  195 - 0xc3
    "11100000", -- 3022 - 0xbce  :  224 - 0xe0
    "11111111", -- 3023 - 0xbcf  :  255 - 0xff
    "01111111", -- 3024 - 0xbd0  :  127 - 0x7f -- Background 0xbd
    "01111111", -- 3025 - 0xbd1  :  127 - 0x7f
    "01111111", -- 3026 - 0xbd2  :  127 - 0x7f
    "11111111", -- 3027 - 0xbd3  :  255 - 0xff
    "11111111", -- 3028 - 0xbd4  :  255 - 0xff
    "11111111", -- 3029 - 0xbd5  :  255 - 0xff
    "11111111", -- 3030 - 0xbd6  :  255 - 0xff
    "11111110", -- 3031 - 0xbd7  :  254 - 0xfe
    "11111111", -- 3032 - 0xbd8  :  255 - 0xff -- plane 1
    "11111111", -- 3033 - 0xbd9  :  255 - 0xff
    "11111111", -- 3034 - 0xbda  :  255 - 0xff
    "11111111", -- 3035 - 0xbdb  :  255 - 0xff
    "11111111", -- 3036 - 0xbdc  :  255 - 0xff
    "11111111", -- 3037 - 0xbdd  :  255 - 0xff
    "11111111", -- 3038 - 0xbde  :  255 - 0xff
    "11111110", -- 3039 - 0xbdf  :  254 - 0xfe
    "11111100", -- 3040 - 0xbe0  :  252 - 0xfc -- Background 0xbe
    "10111000", -- 3041 - 0xbe1  :  184 - 0xb8
    "01111000", -- 3042 - 0xbe2  :  120 - 0x78
    "01111000", -- 3043 - 0xbe3  :  120 - 0x78
    "10110000", -- 3044 - 0xbe4  :  176 - 0xb0
    "01111000", -- 3045 - 0xbe5  :  120 - 0x78
    "11111100", -- 3046 - 0xbe6  :  252 - 0xfc
    "11111110", -- 3047 - 0xbe7  :  254 - 0xfe
    "11111100", -- 3048 - 0xbe8  :  252 - 0xfc -- plane 1
    "11111000", -- 3049 - 0xbe9  :  248 - 0xf8
    "11111000", -- 3050 - 0xbea  :  248 - 0xf8
    "11111000", -- 3051 - 0xbeb  :  248 - 0xf8
    "11111000", -- 3052 - 0xbec  :  248 - 0xf8
    "11111100", -- 3053 - 0xbed  :  252 - 0xfc
    "11111110", -- 3054 - 0xbee  :  254 - 0xfe
    "11111111", -- 3055 - 0xbef  :  255 - 0xff
    "11111111", -- 3056 - 0xbf0  :  255 - 0xff -- Background 0xbf
    "11111111", -- 3057 - 0xbf1  :  255 - 0xff
    "11111111", -- 3058 - 0xbf2  :  255 - 0xff
    "11111111", -- 3059 - 0xbf3  :  255 - 0xff
    "11111111", -- 3060 - 0xbf4  :  255 - 0xff
    "10011100", -- 3061 - 0xbf5  :  156 - 0x9c
    "01000010", -- 3062 - 0xbf6  :   66 - 0x42
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "11111111", -- 3064 - 0xbf8  :  255 - 0xff -- plane 1
    "11111111", -- 3065 - 0xbf9  :  255 - 0xff
    "11111111", -- 3066 - 0xbfa  :  255 - 0xff
    "11111111", -- 3067 - 0xbfb  :  255 - 0xff
    "11111111", -- 3068 - 0xbfc  :  255 - 0xff
    "11111111", -- 3069 - 0xbfd  :  255 - 0xff
    "11111111", -- 3070 - 0xbfe  :  255 - 0xff
    "11111111", -- 3071 - 0xbff  :  255 - 0xff
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00100000", -- 3074 - 0xc02  :   32 - 0x20
    "01000000", -- 3075 - 0xc03  :   64 - 0x40
    "10001010", -- 3076 - 0xc04  :  138 - 0x8a
    "00011110", -- 3077 - 0xc05  :   30 - 0x1e
    "01111110", -- 3078 - 0xc06  :  126 - 0x7e
    "10111110", -- 3079 - 0xc07  :  190 - 0xbe
    "11000000", -- 3080 - 0xc08  :  192 - 0xc0 -- plane 1
    "11110000", -- 3081 - 0xc09  :  240 - 0xf0
    "11111100", -- 3082 - 0xc0a  :  252 - 0xfc
    "11111100", -- 3083 - 0xc0b  :  252 - 0xfc
    "11111110", -- 3084 - 0xc0c  :  254 - 0xfe
    "11111110", -- 3085 - 0xc0d  :  254 - 0xfe
    "11111110", -- 3086 - 0xc0e  :  254 - 0xfe
    "11111110", -- 3087 - 0xc0f  :  254 - 0xfe
    "11011111", -- 3088 - 0xc10  :  223 - 0xdf -- Background 0xc1
    "11111111", -- 3089 - 0xc11  :  255 - 0xff
    "11111110", -- 3090 - 0xc12  :  254 - 0xfe
    "11111100", -- 3091 - 0xc13  :  252 - 0xfc
    "11110000", -- 3092 - 0xc14  :  240 - 0xf0
    "11100000", -- 3093 - 0xc15  :  224 - 0xe0
    "10000000", -- 3094 - 0xc16  :  128 - 0x80
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "11111111", -- 3096 - 0xc18  :  255 - 0xff -- plane 1
    "11111111", -- 3097 - 0xc19  :  255 - 0xff
    "11111110", -- 3098 - 0xc1a  :  254 - 0xfe
    "11111100", -- 3099 - 0xc1b  :  252 - 0xfc
    "11110000", -- 3100 - 0xc1c  :  240 - 0xf0
    "11100000", -- 3101 - 0xc1d  :  224 - 0xe0
    "10000000", -- 3102 - 0xc1e  :  128 - 0x80
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000100", -- 3106 - 0xc22  :    4 - 0x4
    "00000010", -- 3107 - 0xc23  :    2 - 0x2
    "01010001", -- 3108 - 0xc24  :   81 - 0x51
    "01111000", -- 3109 - 0xc25  :  120 - 0x78
    "01111110", -- 3110 - 0xc26  :  126 - 0x7e
    "11111101", -- 3111 - 0xc27  :  253 - 0xfd
    "00000011", -- 3112 - 0xc28  :    3 - 0x3 -- plane 1
    "00001111", -- 3113 - 0xc29  :   15 - 0xf
    "00111111", -- 3114 - 0xc2a  :   63 - 0x3f
    "00111111", -- 3115 - 0xc2b  :   63 - 0x3f
    "01111111", -- 3116 - 0xc2c  :  127 - 0x7f
    "01111111", -- 3117 - 0xc2d  :  127 - 0x7f
    "01111110", -- 3118 - 0xc2e  :  126 - 0x7e
    "11111111", -- 3119 - 0xc2f  :  255 - 0xff
    "11111011", -- 3120 - 0xc30  :  251 - 0xfb -- Background 0xc3
    "11111111", -- 3121 - 0xc31  :  255 - 0xff
    "01111111", -- 3122 - 0xc32  :  127 - 0x7f
    "00111111", -- 3123 - 0xc33  :   63 - 0x3f
    "00001111", -- 3124 - 0xc34  :   15 - 0xf
    "00000111", -- 3125 - 0xc35  :    7 - 0x7
    "00000001", -- 3126 - 0xc36  :    1 - 0x1
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "11111111", -- 3128 - 0xc38  :  255 - 0xff -- plane 1
    "11111111", -- 3129 - 0xc39  :  255 - 0xff
    "01111111", -- 3130 - 0xc3a  :  127 - 0x7f
    "00111111", -- 3131 - 0xc3b  :   63 - 0x3f
    "00001111", -- 3132 - 0xc3c  :   15 - 0xf
    "00000111", -- 3133 - 0xc3d  :    7 - 0x7
    "00000001", -- 3134 - 0xc3e  :    1 - 0x1
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0xc4
    "10000000", -- 3137 - 0xc41  :  128 - 0x80
    "01000000", -- 3138 - 0xc42  :   64 - 0x40
    "11100000", -- 3139 - 0xc43  :  224 - 0xe0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "00000100", -- 3142 - 0xc46  :    4 - 0x4
    "11111111", -- 3143 - 0xc47  :  255 - 0xff
    "11000000", -- 3144 - 0xc48  :  192 - 0xc0 -- plane 1
    "11100000", -- 3145 - 0xc49  :  224 - 0xe0
    "11110000", -- 3146 - 0xc4a  :  240 - 0xf0
    "11100000", -- 3147 - 0xc4b  :  224 - 0xe0
    "11100001", -- 3148 - 0xc4c  :  225 - 0xe1
    "11000011", -- 3149 - 0xc4d  :  195 - 0xc3
    "00000111", -- 3150 - 0xc4e  :    7 - 0x7
    "11111111", -- 3151 - 0xc4f  :  255 - 0xff
    "11111110", -- 3152 - 0xc50  :  254 - 0xfe -- Background 0xc5
    "11111110", -- 3153 - 0xc51  :  254 - 0xfe
    "11111110", -- 3154 - 0xc52  :  254 - 0xfe
    "11111111", -- 3155 - 0xc53  :  255 - 0xff
    "11111111", -- 3156 - 0xc54  :  255 - 0xff
    "11111111", -- 3157 - 0xc55  :  255 - 0xff
    "11111111", -- 3158 - 0xc56  :  255 - 0xff
    "01111111", -- 3159 - 0xc57  :  127 - 0x7f
    "11111111", -- 3160 - 0xc58  :  255 - 0xff -- plane 1
    "11111111", -- 3161 - 0xc59  :  255 - 0xff
    "11111111", -- 3162 - 0xc5a  :  255 - 0xff
    "11111111", -- 3163 - 0xc5b  :  255 - 0xff
    "11111111", -- 3164 - 0xc5c  :  255 - 0xff
    "11111111", -- 3165 - 0xc5d  :  255 - 0xff
    "11111111", -- 3166 - 0xc5e  :  255 - 0xff
    "01111111", -- 3167 - 0xc5f  :  127 - 0x7f
    "00111111", -- 3168 - 0xc60  :   63 - 0x3f -- Background 0xc6
    "00011101", -- 3169 - 0xc61  :   29 - 0x1d
    "00011110", -- 3170 - 0xc62  :   30 - 0x1e
    "00011110", -- 3171 - 0xc63  :   30 - 0x1e
    "00001101", -- 3172 - 0xc64  :   13 - 0xd
    "00011110", -- 3173 - 0xc65  :   30 - 0x1e
    "00111111", -- 3174 - 0xc66  :   63 - 0x3f
    "01111111", -- 3175 - 0xc67  :  127 - 0x7f
    "00111111", -- 3176 - 0xc68  :   63 - 0x3f -- plane 1
    "00011111", -- 3177 - 0xc69  :   31 - 0x1f
    "00011111", -- 3178 - 0xc6a  :   31 - 0x1f
    "00011111", -- 3179 - 0xc6b  :   31 - 0x1f
    "00011111", -- 3180 - 0xc6c  :   31 - 0x1f
    "00111111", -- 3181 - 0xc6d  :   63 - 0x3f
    "01111111", -- 3182 - 0xc6e  :  127 - 0x7f
    "11111111", -- 3183 - 0xc6f  :  255 - 0xff
    "11111111", -- 3184 - 0xc70  :  255 - 0xff -- Background 0xc7
    "11111111", -- 3185 - 0xc71  :  255 - 0xff
    "11111111", -- 3186 - 0xc72  :  255 - 0xff
    "11111111", -- 3187 - 0xc73  :  255 - 0xff
    "11111111", -- 3188 - 0xc74  :  255 - 0xff
    "00111001", -- 3189 - 0xc75  :   57 - 0x39
    "01000010", -- 3190 - 0xc76  :   66 - 0x42
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "11111111", -- 3192 - 0xc78  :  255 - 0xff -- plane 1
    "11111111", -- 3193 - 0xc79  :  255 - 0xff
    "11111111", -- 3194 - 0xc7a  :  255 - 0xff
    "11111111", -- 3195 - 0xc7b  :  255 - 0xff
    "11111111", -- 3196 - 0xc7c  :  255 - 0xff
    "11111111", -- 3197 - 0xc7d  :  255 - 0xff
    "11111111", -- 3198 - 0xc7e  :  255 - 0xff
    "11111111", -- 3199 - 0xc7f  :  255 - 0xff
    "01101111", -- 3200 - 0xc80  :  111 - 0x6f -- Background 0xc8
    "11011011", -- 3201 - 0xc81  :  219 - 0xdb
    "00000011", -- 3202 - 0xc82  :    3 - 0x3
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "11111111", -- 3208 - 0xc88  :  255 - 0xff -- plane 1
    "11111111", -- 3209 - 0xc89  :  255 - 0xff
    "00000011", -- 3210 - 0xc8a  :    3 - 0x3
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 3217 - 0xc91  :    0 - 0x0
    "00000000", -- 3218 - 0xc92  :    0 - 0x0
    "00000000", -- 3219 - 0xc93  :    0 - 0x0
    "00000000", -- 3220 - 0xc94  :    0 - 0x0
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "11100000", -- 3223 - 0xc97  :  224 - 0xe0
    "00000000", -- 3224 - 0xc98  :    0 - 0x0 -- plane 1
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00000000", -- 3226 - 0xc9a  :    0 - 0x0
    "00000000", -- 3227 - 0xc9b  :    0 - 0x0
    "10000000", -- 3228 - 0xc9c  :  128 - 0x80
    "11000000", -- 3229 - 0xc9d  :  192 - 0xc0
    "11000000", -- 3230 - 0xc9e  :  192 - 0xc0
    "11110000", -- 3231 - 0xc9f  :  240 - 0xf0
    "01110000", -- 3232 - 0xca0  :  112 - 0x70 -- Background 0xca
    "01111100", -- 3233 - 0xca1  :  124 - 0x7c
    "01111110", -- 3234 - 0xca2  :  126 - 0x7e
    "11111111", -- 3235 - 0xca3  :  255 - 0xff
    "11111111", -- 3236 - 0xca4  :  255 - 0xff
    "11110111", -- 3237 - 0xca5  :  247 - 0xf7
    "11101111", -- 3238 - 0xca6  :  239 - 0xef
    "00011111", -- 3239 - 0xca7  :   31 - 0x1f
    "11111100", -- 3240 - 0xca8  :  252 - 0xfc -- plane 1
    "11111110", -- 3241 - 0xca9  :  254 - 0xfe
    "11111111", -- 3242 - 0xcaa  :  255 - 0xff
    "11111111", -- 3243 - 0xcab  :  255 - 0xff
    "11111111", -- 3244 - 0xcac  :  255 - 0xff
    "11111111", -- 3245 - 0xcad  :  255 - 0xff
    "11111111", -- 3246 - 0xcae  :  255 - 0xff
    "11111111", -- 3247 - 0xcaf  :  255 - 0xff
    "11111111", -- 3248 - 0xcb0  :  255 - 0xff -- Background 0xcb
    "11111111", -- 3249 - 0xcb1  :  255 - 0xff
    "11111111", -- 3250 - 0xcb2  :  255 - 0xff
    "11111000", -- 3251 - 0xcb3  :  248 - 0xf8
    "11111000", -- 3252 - 0xcb4  :  248 - 0xf8
    "11111110", -- 3253 - 0xcb5  :  254 - 0xfe
    "11111111", -- 3254 - 0xcb6  :  255 - 0xff
    "11111111", -- 3255 - 0xcb7  :  255 - 0xff
    "11111111", -- 3256 - 0xcb8  :  255 - 0xff -- plane 1
    "11111111", -- 3257 - 0xcb9  :  255 - 0xff
    "11111111", -- 3258 - 0xcba  :  255 - 0xff
    "11111000", -- 3259 - 0xcbb  :  248 - 0xf8
    "11111110", -- 3260 - 0xcbc  :  254 - 0xfe
    "11111111", -- 3261 - 0xcbd  :  255 - 0xff
    "11111111", -- 3262 - 0xcbe  :  255 - 0xff
    "11111111", -- 3263 - 0xcbf  :  255 - 0xff
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff -- Background 0xcc
    "11111111", -- 3265 - 0xcc1  :  255 - 0xff
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "00111111", -- 3267 - 0xcc3  :   63 - 0x3f
    "00011110", -- 3268 - 0xcc4  :   30 - 0x1e
    "00000001", -- 3269 - 0xcc5  :    1 - 0x1
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "11111111", -- 3272 - 0xcc8  :  255 - 0xff -- plane 1
    "11111111", -- 3273 - 0xcc9  :  255 - 0xff
    "11111111", -- 3274 - 0xcca  :  255 - 0xff
    "00111111", -- 3275 - 0xccb  :   63 - 0x3f
    "00011111", -- 3276 - 0xccc  :   31 - 0x1f
    "00011111", -- 3277 - 0xccd  :   31 - 0x1f
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "10000000", -- 3283 - 0xcd3  :  128 - 0x80
    "11000000", -- 3284 - 0xcd4  :  192 - 0xc0
    "11100000", -- 3285 - 0xcd5  :  224 - 0xe0
    "11100000", -- 3286 - 0xcd6  :  224 - 0xe0
    "11100000", -- 3287 - 0xcd7  :  224 - 0xe0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "10000000", -- 3290 - 0xcda  :  128 - 0x80
    "11000000", -- 3291 - 0xcdb  :  192 - 0xc0
    "11100000", -- 3292 - 0xcdc  :  224 - 0xe0
    "11100000", -- 3293 - 0xcdd  :  224 - 0xe0
    "11100000", -- 3294 - 0xcde  :  224 - 0xe0
    "11100000", -- 3295 - 0xcdf  :  224 - 0xe0
    "11000000", -- 3296 - 0xce0  :  192 - 0xc0 -- Background 0xce
    "10000000", -- 3297 - 0xce1  :  128 - 0x80
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "10000000", -- 3302 - 0xce6  :  128 - 0x80
    "10000000", -- 3303 - 0xce7  :  128 - 0x80
    "11000000", -- 3304 - 0xce8  :  192 - 0xc0 -- plane 1
    "10000000", -- 3305 - 0xce9  :  128 - 0x80
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "10000000", -- 3309 - 0xced  :  128 - 0x80
    "11000000", -- 3310 - 0xcee  :  192 - 0xc0
    "11000000", -- 3311 - 0xcef  :  192 - 0xc0
    "10000000", -- 3312 - 0xcf0  :  128 - 0x80 -- Background 0xcf
    "10000000", -- 3313 - 0xcf1  :  128 - 0x80
    "11100000", -- 3314 - 0xcf2  :  224 - 0xe0
    "11000000", -- 3315 - 0xcf3  :  192 - 0xc0
    "00100000", -- 3316 - 0xcf4  :   32 - 0x20
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "11000000", -- 3320 - 0xcf8  :  192 - 0xc0 -- plane 1
    "11000000", -- 3321 - 0xcf9  :  192 - 0xc0
    "11100000", -- 3322 - 0xcfa  :  224 - 0xe0
    "11111000", -- 3323 - 0xcfb  :  248 - 0xf8
    "11111100", -- 3324 - 0xcfc  :  252 - 0xfc
    "11111100", -- 3325 - 0xcfd  :  252 - 0xfc
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00011111", -- 3328 - 0xd00  :   31 - 0x1f -- Background 0xd0
    "00000110", -- 3329 - 0xd01  :    6 - 0x6
    "00000110", -- 3330 - 0xd02  :    6 - 0x6
    "00000110", -- 3331 - 0xd03  :    6 - 0x6
    "00000110", -- 3332 - 0xd04  :    6 - 0x6
    "00000110", -- 3333 - 0xd05  :    6 - 0x6
    "00000110", -- 3334 - 0xd06  :    6 - 0x6
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- plane 1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00111001", -- 3344 - 0xd10  :   57 - 0x39 -- Background 0xd1
    "01100101", -- 3345 - 0xd11  :  101 - 0x65
    "01100101", -- 3346 - 0xd12  :  101 - 0x65
    "01100101", -- 3347 - 0xd13  :  101 - 0x65
    "01100101", -- 3348 - 0xd14  :  101 - 0x65
    "01100101", -- 3349 - 0xd15  :  101 - 0x65
    "00111001", -- 3350 - 0xd16  :   57 - 0x39
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0 -- plane 1
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "11100000", -- 3360 - 0xd20  :  224 - 0xe0 -- Background 0xd2
    "10110000", -- 3361 - 0xd21  :  176 - 0xb0
    "10110000", -- 3362 - 0xd22  :  176 - 0xb0
    "10110110", -- 3363 - 0xd23  :  182 - 0xb6
    "11100110", -- 3364 - 0xd24  :  230 - 0xe6
    "10000000", -- 3365 - 0xd25  :  128 - 0x80
    "10000000", -- 3366 - 0xd26  :  128 - 0x80
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- plane 1
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000000", -- 3372 - 0xd2c  :    0 - 0x0
    "00000000", -- 3373 - 0xd2d  :    0 - 0x0
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00111100", -- 3376 - 0xd30  :   60 - 0x3c -- Background 0xd3
    "01000010", -- 3377 - 0xd31  :   66 - 0x42
    "10011001", -- 3378 - 0xd32  :  153 - 0x99
    "10100001", -- 3379 - 0xd33  :  161 - 0xa1
    "10100001", -- 3380 - 0xd34  :  161 - 0xa1
    "10011001", -- 3381 - 0xd35  :  153 - 0x99
    "01000010", -- 3382 - 0xd36  :   66 - 0x42
    "00111100", -- 3383 - 0xd37  :   60 - 0x3c
    "00000000", -- 3384 - 0xd38  :    0 - 0x0 -- plane 1
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "00000000", -- 3386 - 0xd3a  :    0 - 0x0
    "00000000", -- 3387 - 0xd3b  :    0 - 0x0
    "00000000", -- 3388 - 0xd3c  :    0 - 0x0
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00000011", -- 3395 - 0xd43  :    3 - 0x3
    "00000110", -- 3396 - 0xd44  :    6 - 0x6
    "00000000", -- 3397 - 0xd45  :    0 - 0x0
    "00000001", -- 3398 - 0xd46  :    1 - 0x1
    "00000111", -- 3399 - 0xd47  :    7 - 0x7
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- plane 1
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000011", -- 3404 - 0xd4c  :    3 - 0x3
    "00000111", -- 3405 - 0xd4d  :    7 - 0x7
    "00000011", -- 3406 - 0xd4e  :    3 - 0x3
    "00000111", -- 3407 - 0xd4f  :    7 - 0x7
    "00001111", -- 3408 - 0xd50  :   15 - 0xf -- Background 0xd5
    "00011111", -- 3409 - 0xd51  :   31 - 0x1f
    "00111111", -- 3410 - 0xd52  :   63 - 0x3f
    "01111111", -- 3411 - 0xd53  :  127 - 0x7f
    "01111111", -- 3412 - 0xd54  :  127 - 0x7f
    "01111111", -- 3413 - 0xd55  :  127 - 0x7f
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "01111111", -- 3415 - 0xd57  :  127 - 0x7f
    "00011111", -- 3416 - 0xd58  :   31 - 0x1f -- plane 1
    "00111111", -- 3417 - 0xd59  :   63 - 0x3f
    "01111111", -- 3418 - 0xd5a  :  127 - 0x7f
    "11111111", -- 3419 - 0xd5b  :  255 - 0xff
    "11111111", -- 3420 - 0xd5c  :  255 - 0xff
    "11111111", -- 3421 - 0xd5d  :  255 - 0xff
    "11111111", -- 3422 - 0xd5e  :  255 - 0xff
    "01111111", -- 3423 - 0xd5f  :  127 - 0x7f
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "10000000", -- 3427 - 0xd63  :  128 - 0x80
    "00000000", -- 3428 - 0xd64  :    0 - 0x0
    "00000000", -- 3429 - 0xd65  :    0 - 0x0
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "10100000", -- 3431 - 0xd67  :  160 - 0xa0
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- plane 1
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "11000000", -- 3435 - 0xd6b  :  192 - 0xc0
    "11100000", -- 3436 - 0xd6c  :  224 - 0xe0
    "11110000", -- 3437 - 0xd6d  :  240 - 0xf0
    "11110000", -- 3438 - 0xd6e  :  240 - 0xf0
    "11111000", -- 3439 - 0xd6f  :  248 - 0xf8
    "11100000", -- 3440 - 0xd70  :  224 - 0xe0 -- Background 0xd7
    "11110000", -- 3441 - 0xd71  :  240 - 0xf0
    "11100000", -- 3442 - 0xd72  :  224 - 0xe0
    "11011101", -- 3443 - 0xd73  :  221 - 0xdd
    "11111010", -- 3444 - 0xd74  :  250 - 0xfa
    "11101011", -- 3445 - 0xd75  :  235 - 0xeb
    "10000000", -- 3446 - 0xd76  :  128 - 0x80
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "11111100", -- 3448 - 0xd78  :  252 - 0xfc -- plane 1
    "11111000", -- 3449 - 0xd79  :  248 - 0xf8
    "11110000", -- 3450 - 0xd7a  :  240 - 0xf0
    "11111111", -- 3451 - 0xd7b  :  255 - 0xff
    "11111111", -- 3452 - 0xd7c  :  255 - 0xff
    "11111111", -- 3453 - 0xd7d  :  255 - 0xff
    "11111111", -- 3454 - 0xd7e  :  255 - 0xff
    "11111111", -- 3455 - 0xd7f  :  255 - 0xff
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000011", -- 3459 - 0xd83  :    3 - 0x3
    "00000110", -- 3460 - 0xd84  :    6 - 0x6
    "00000000", -- 3461 - 0xd85  :    0 - 0x0
    "00000001", -- 3462 - 0xd86  :    1 - 0x1
    "00000001", -- 3463 - 0xd87  :    1 - 0x1
    "00000000", -- 3464 - 0xd88  :    0 - 0x0 -- plane 1
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "00000000", -- 3467 - 0xd8b  :    0 - 0x0
    "00000011", -- 3468 - 0xd8c  :    3 - 0x3
    "00000111", -- 3469 - 0xd8d  :    7 - 0x7
    "00001111", -- 3470 - 0xd8e  :   15 - 0xf
    "00011111", -- 3471 - 0xd8f  :   31 - 0x1f
    "00001011", -- 3472 - 0xd90  :   11 - 0xb -- Background 0xd9
    "00000111", -- 3473 - 0xd91  :    7 - 0x7
    "00000011", -- 3474 - 0xd92  :    3 - 0x3
    "01011101", -- 3475 - 0xd93  :   93 - 0x5d
    "10101111", -- 3476 - 0xd94  :  175 - 0xaf
    "01010011", -- 3477 - 0xd95  :   83 - 0x53
    "00000000", -- 3478 - 0xd96  :    0 - 0x0
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "00111111", -- 3480 - 0xd98  :   63 - 0x3f -- plane 1
    "00011111", -- 3481 - 0xd99  :   31 - 0x1f
    "00000111", -- 3482 - 0xd9a  :    7 - 0x7
    "11111111", -- 3483 - 0xd9b  :  255 - 0xff
    "11111111", -- 3484 - 0xd9c  :  255 - 0xff
    "11111111", -- 3485 - 0xd9d  :  255 - 0xff
    "11111111", -- 3486 - 0xd9e  :  255 - 0xff
    "11111111", -- 3487 - 0xd9f  :  255 - 0xff
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000000", -- 3490 - 0xda2  :    0 - 0x0
    "10000000", -- 3491 - 0xda3  :  128 - 0x80
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "01100000", -- 3494 - 0xda6  :   96 - 0x60
    "11110000", -- 3495 - 0xda7  :  240 - 0xf0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0 -- plane 1
    "00000000", -- 3497 - 0xda9  :    0 - 0x0
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "11000000", -- 3499 - 0xdab  :  192 - 0xc0
    "11000000", -- 3500 - 0xdac  :  192 - 0xc0
    "11000000", -- 3501 - 0xdad  :  192 - 0xc0
    "11100000", -- 3502 - 0xdae  :  224 - 0xe0
    "11111000", -- 3503 - 0xdaf  :  248 - 0xf8
    "11111000", -- 3504 - 0xdb0  :  248 - 0xf8 -- Background 0xdb
    "11111100", -- 3505 - 0xdb1  :  252 - 0xfc
    "11111100", -- 3506 - 0xdb2  :  252 - 0xfc
    "11111110", -- 3507 - 0xdb3  :  254 - 0xfe
    "11111110", -- 3508 - 0xdb4  :  254 - 0xfe
    "11111111", -- 3509 - 0xdb5  :  255 - 0xff
    "11111111", -- 3510 - 0xdb6  :  255 - 0xff
    "01111110", -- 3511 - 0xdb7  :  126 - 0x7e
    "11111100", -- 3512 - 0xdb8  :  252 - 0xfc -- plane 1
    "11111110", -- 3513 - 0xdb9  :  254 - 0xfe
    "11111110", -- 3514 - 0xdba  :  254 - 0xfe
    "11111111", -- 3515 - 0xdbb  :  255 - 0xff
    "11111111", -- 3516 - 0xdbc  :  255 - 0xff
    "11111111", -- 3517 - 0xdbd  :  255 - 0xff
    "11111111", -- 3518 - 0xdbe  :  255 - 0xff
    "11111110", -- 3519 - 0xdbf  :  254 - 0xfe
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00000000", -- 3523 - 0xdc3  :    0 - 0x0
    "00000000", -- 3524 - 0xdc4  :    0 - 0x0
    "00000000", -- 3525 - 0xdc5  :    0 - 0x0
    "00100001", -- 3526 - 0xdc6  :   33 - 0x21
    "00111111", -- 3527 - 0xdc7  :   63 - 0x3f
    "00110110", -- 3528 - 0xdc8  :   54 - 0x36 -- plane 1
    "00110110", -- 3529 - 0xdc9  :   54 - 0x36
    "01111110", -- 3530 - 0xdca  :  126 - 0x7e
    "01111111", -- 3531 - 0xdcb  :  127 - 0x7f
    "01111111", -- 3532 - 0xdcc  :  127 - 0x7f
    "01111111", -- 3533 - 0xdcd  :  127 - 0x7f
    "00111111", -- 3534 - 0xdce  :   63 - 0x3f
    "00111111", -- 3535 - 0xdcf  :   63 - 0x3f
    "00111111", -- 3536 - 0xdd0  :   63 - 0x3f -- Background 0xdd
    "00011111", -- 3537 - 0xdd1  :   31 - 0x1f
    "00011111", -- 3538 - 0xdd2  :   31 - 0x1f
    "00001111", -- 3539 - 0xdd3  :   15 - 0xf
    "00000111", -- 3540 - 0xdd4  :    7 - 0x7
    "00000011", -- 3541 - 0xdd5  :    3 - 0x3
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00111111", -- 3544 - 0xdd8  :   63 - 0x3f -- plane 1
    "00011111", -- 3545 - 0xdd9  :   31 - 0x1f
    "00011111", -- 3546 - 0xdda  :   31 - 0x1f
    "00001111", -- 3547 - 0xddb  :   15 - 0xf
    "00000111", -- 3548 - 0xddc  :    7 - 0x7
    "00000011", -- 3549 - 0xddd  :    3 - 0x3
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00111110", -- 3552 - 0xde0  :   62 - 0x3e -- Background 0xde
    "00011110", -- 3553 - 0xde1  :   30 - 0x1e
    "00011110", -- 3554 - 0xde2  :   30 - 0x1e
    "00001110", -- 3555 - 0xde3  :   14 - 0xe
    "00001111", -- 3556 - 0xde4  :   15 - 0xf
    "00011111", -- 3557 - 0xde5  :   31 - 0x1f
    "10011111", -- 3558 - 0xde6  :  159 - 0x9f
    "10011111", -- 3559 - 0xde7  :  159 - 0x9f
    "00111111", -- 3560 - 0xde8  :   63 - 0x3f -- plane 1
    "00011111", -- 3561 - 0xde9  :   31 - 0x1f
    "11011111", -- 3562 - 0xdea  :  223 - 0xdf
    "11001111", -- 3563 - 0xdeb  :  207 - 0xcf
    "11001111", -- 3564 - 0xdec  :  207 - 0xcf
    "10011111", -- 3565 - 0xded  :  159 - 0x9f
    "11011111", -- 3566 - 0xdee  :  223 - 0xdf
    "11111111", -- 3567 - 0xdef  :  255 - 0xff
    "11011111", -- 3568 - 0xdf0  :  223 - 0xdf -- Background 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "11111111", -- 3570 - 0xdf2  :  255 - 0xff
    "11111111", -- 3571 - 0xdf3  :  255 - 0xff
    "11111111", -- 3572 - 0xdf4  :  255 - 0xff
    "11011111", -- 3573 - 0xdf5  :  223 - 0xdf
    "11100111", -- 3574 - 0xdf6  :  231 - 0xe7
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "11111111", -- 3576 - 0xdf8  :  255 - 0xff -- plane 1
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11111111", -- 3580 - 0xdfc  :  255 - 0xff
    "11111111", -- 3581 - 0xdfd  :  255 - 0xff
    "11111111", -- 3582 - 0xdfe  :  255 - 0xff
    "00001111", -- 3583 - 0xdff  :   15 - 0xf
    "00100000", -- 3584 - 0xe00  :   32 - 0x20 -- Background 0xe0
    "00001111", -- 3585 - 0xe01  :   15 - 0xf
    "00110000", -- 3586 - 0xe02  :   48 - 0x30
    "01000000", -- 3587 - 0xe03  :   64 - 0x40
    "10011000", -- 3588 - 0xe04  :  152 - 0x98
    "00111110", -- 3589 - 0xe05  :   62 - 0x3e
    "00011111", -- 3590 - 0xe06  :   31 - 0x1f
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "11111111", -- 3592 - 0xe08  :  255 - 0xff -- plane 1
    "11111111", -- 3593 - 0xe09  :  255 - 0xff
    "11111111", -- 3594 - 0xe0a  :  255 - 0xff
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "11111111", -- 3596 - 0xe0c  :  255 - 0xff
    "11111111", -- 3597 - 0xe0d  :  255 - 0xff
    "11111111", -- 3598 - 0xe0e  :  255 - 0xff
    "11111111", -- 3599 - 0xe0f  :  255 - 0xff
    "10000001", -- 3600 - 0xe10  :  129 - 0x81 -- Background 0xe1
    "00110110", -- 3601 - 0xe11  :   54 - 0x36
    "00101110", -- 3602 - 0xe12  :   46 - 0x2e
    "10101111", -- 3603 - 0xe13  :  175 - 0xaf
    "10101110", -- 3604 - 0xe14  :  174 - 0xae
    "11010001", -- 3605 - 0xe15  :  209 - 0xd1
    "11101111", -- 3606 - 0xe16  :  239 - 0xef
    "10000111", -- 3607 - 0xe17  :  135 - 0x87
    "11111111", -- 3608 - 0xe18  :  255 - 0xff -- plane 1
    "11111001", -- 3609 - 0xe19  :  249 - 0xf9
    "11110000", -- 3610 - 0xe1a  :  240 - 0xf0
    "11110000", -- 3611 - 0xe1b  :  240 - 0xf0
    "10110001", -- 3612 - 0xe1c  :  177 - 0xb1
    "11011111", -- 3613 - 0xe1d  :  223 - 0xdf
    "11101111", -- 3614 - 0xe1e  :  239 - 0xef
    "10000111", -- 3615 - 0xe1f  :  135 - 0x87
    "00000010", -- 3616 - 0xe20  :    2 - 0x2 -- Background 0xe2
    "11111000", -- 3617 - 0xe21  :  248 - 0xf8
    "00000110", -- 3618 - 0xe22  :    6 - 0x6
    "00000001", -- 3619 - 0xe23  :    1 - 0x1
    "00001100", -- 3620 - 0xe24  :   12 - 0xc
    "00111110", -- 3621 - 0xe25  :   62 - 0x3e
    "11111100", -- 3622 - 0xe26  :  252 - 0xfc
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "11111111", -- 3624 - 0xe28  :  255 - 0xff -- plane 1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "11111111", -- 3631 - 0xe2f  :  255 - 0xff
    "11000000", -- 3632 - 0xe30  :  192 - 0xc0 -- Background 0xe3
    "00110110", -- 3633 - 0xe31  :   54 - 0x36
    "00111110", -- 3634 - 0xe32  :   62 - 0x3e
    "01111010", -- 3635 - 0xe33  :  122 - 0x7a
    "10110110", -- 3636 - 0xe34  :  182 - 0xb6
    "11001101", -- 3637 - 0xe35  :  205 - 0xcd
    "11111011", -- 3638 - 0xe36  :  251 - 0xfb
    "11110000", -- 3639 - 0xe37  :  240 - 0xf0
    "11111111", -- 3640 - 0xe38  :  255 - 0xff -- plane 1
    "11001111", -- 3641 - 0xe39  :  207 - 0xcf
    "10000111", -- 3642 - 0xe3a  :  135 - 0x87
    "10000111", -- 3643 - 0xe3b  :  135 - 0x87
    "11001110", -- 3644 - 0xe3c  :  206 - 0xce
    "11111101", -- 3645 - 0xe3d  :  253 - 0xfd
    "11111011", -- 3646 - 0xe3e  :  251 - 0xfb
    "11110000", -- 3647 - 0xe3f  :  240 - 0xf0
    "00111110", -- 3648 - 0xe40  :   62 - 0x3e -- Background 0xe4
    "00111100", -- 3649 - 0xe41  :   60 - 0x3c
    "00111100", -- 3650 - 0xe42  :   60 - 0x3c
    "00111000", -- 3651 - 0xe43  :   56 - 0x38
    "11111000", -- 3652 - 0xe44  :  248 - 0xf8
    "01111100", -- 3653 - 0xe45  :  124 - 0x7c
    "01111110", -- 3654 - 0xe46  :  126 - 0x7e
    "01111000", -- 3655 - 0xe47  :  120 - 0x78
    "11111110", -- 3656 - 0xe48  :  254 - 0xfe -- plane 1
    "11111100", -- 3657 - 0xe49  :  252 - 0xfc
    "11111100", -- 3658 - 0xe4a  :  252 - 0xfc
    "11111000", -- 3659 - 0xe4b  :  248 - 0xf8
    "11111011", -- 3660 - 0xe4c  :  251 - 0xfb
    "11111101", -- 3661 - 0xe4d  :  253 - 0xfd
    "11111110", -- 3662 - 0xe4e  :  254 - 0xfe
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "11111000", -- 3664 - 0xe50  :  248 - 0xf8 -- Background 0xe5
    "01111111", -- 3665 - 0xe51  :  127 - 0x7f
    "01111111", -- 3666 - 0xe52  :  127 - 0x7f
    "11111110", -- 3667 - 0xe53  :  254 - 0xfe
    "11111111", -- 3668 - 0xe54  :  255 - 0xff
    "11111111", -- 3669 - 0xe55  :  255 - 0xff
    "11110011", -- 3670 - 0xe56  :  243 - 0xf3
    "10000001", -- 3671 - 0xe57  :  129 - 0x81
    "11111111", -- 3672 - 0xe58  :  255 - 0xff -- plane 1
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "11111111", -- 3674 - 0xe5a  :  255 - 0xff
    "11111111", -- 3675 - 0xe5b  :  255 - 0xff
    "11111111", -- 3676 - 0xe5c  :  255 - 0xff
    "11111111", -- 3677 - 0xe5d  :  255 - 0xff
    "11111111", -- 3678 - 0xe5e  :  255 - 0xff
    "11111001", -- 3679 - 0xe5f  :  249 - 0xf9
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00010000", -- 3683 - 0xe63  :   16 - 0x10
    "01000000", -- 3684 - 0xe64  :   64 - 0x40
    "00100000", -- 3685 - 0xe65  :   32 - 0x20
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- plane 1
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "01111000", -- 3691 - 0xe6b  :  120 - 0x78
    "11111100", -- 3692 - 0xe6c  :  252 - 0xfc
    "11111100", -- 3693 - 0xe6d  :  252 - 0xfc
    "11111100", -- 3694 - 0xe6e  :  252 - 0xfc
    "11111100", -- 3695 - 0xe6f  :  252 - 0xfc
    "00000110", -- 3696 - 0xe70  :    6 - 0x6 -- Background 0xe7
    "00001110", -- 3697 - 0xe71  :   14 - 0xe
    "01111110", -- 3698 - 0xe72  :  126 - 0x7e
    "11111110", -- 3699 - 0xe73  :  254 - 0xfe
    "11111110", -- 3700 - 0xe74  :  254 - 0xfe
    "11111100", -- 3701 - 0xe75  :  252 - 0xfc
    "11111000", -- 3702 - 0xe76  :  248 - 0xf8
    "11110000", -- 3703 - 0xe77  :  240 - 0xf0
    "11111110", -- 3704 - 0xe78  :  254 - 0xfe -- plane 1
    "11111110", -- 3705 - 0xe79  :  254 - 0xfe
    "11111110", -- 3706 - 0xe7a  :  254 - 0xfe
    "11111110", -- 3707 - 0xe7b  :  254 - 0xfe
    "11111110", -- 3708 - 0xe7c  :  254 - 0xfe
    "11111100", -- 3709 - 0xe7d  :  252 - 0xfc
    "11111000", -- 3710 - 0xe7e  :  248 - 0xf8
    "11110000", -- 3711 - 0xe7f  :  240 - 0xf0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000001", -- 3719 - 0xe87  :    1 - 0x1
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- plane 1
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000010", -- 3728 - 0xe90  :    2 - 0x2 -- Background 0xe9
    "00000000", -- 3729 - 0xe91  :    0 - 0x0
    "00001000", -- 3730 - 0xe92  :    8 - 0x8
    "00000001", -- 3731 - 0xe93  :    1 - 0x1
    "00010011", -- 3732 - 0xe94  :   19 - 0x13
    "00000001", -- 3733 - 0xe95  :    1 - 0x1
    "00000000", -- 3734 - 0xe96  :    0 - 0x0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00000001", -- 3736 - 0xe98  :    1 - 0x1 -- plane 1
    "00001111", -- 3737 - 0xe99  :   15 - 0xf
    "00011111", -- 3738 - 0xe9a  :   31 - 0x1f
    "00011111", -- 3739 - 0xe9b  :   31 - 0x1f
    "00111011", -- 3740 - 0xe9c  :   59 - 0x3b
    "00110011", -- 3741 - 0xe9d  :   51 - 0x33
    "00000001", -- 3742 - 0xe9e  :    1 - 0x1
    "00000001", -- 3743 - 0xe9f  :    1 - 0x1
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xea
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0 -- plane 1
    "00000000", -- 3753 - 0xea9  :    0 - 0x0
    "00000000", -- 3754 - 0xeaa  :    0 - 0x0
    "00110110", -- 3755 - 0xeab  :   54 - 0x36
    "01101100", -- 3756 - 0xeac  :  108 - 0x6c
    "11111101", -- 3757 - 0xead  :  253 - 0xfd
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xeb
    "01000011", -- 3761 - 0xeb1  :   67 - 0x43
    "01111111", -- 3762 - 0xeb2  :  127 - 0x7f
    "01111111", -- 3763 - 0xeb3  :  127 - 0x7f
    "01111111", -- 3764 - 0xeb4  :  127 - 0x7f
    "00111111", -- 3765 - 0xeb5  :   63 - 0x3f
    "00011111", -- 3766 - 0xeb6  :   31 - 0x1f
    "00000111", -- 3767 - 0xeb7  :    7 - 0x7
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff -- plane 1
    "01111111", -- 3769 - 0xeb9  :  127 - 0x7f
    "01111111", -- 3770 - 0xeba  :  127 - 0x7f
    "01111111", -- 3771 - 0xebb  :  127 - 0x7f
    "01111111", -- 3772 - 0xebc  :  127 - 0x7f
    "00111111", -- 3773 - 0xebd  :   63 - 0x3f
    "00011111", -- 3774 - 0xebe  :   31 - 0x1f
    "00000111", -- 3775 - 0xebf  :    7 - 0x7
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "11000000", -- 3782 - 0xec6  :  192 - 0xc0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "11100000", -- 3791 - 0xecf  :  224 - 0xe0
    "00010000", -- 3792 - 0xed0  :   16 - 0x10 -- Background 0xed
    "00111000", -- 3793 - 0xed1  :   56 - 0x38
    "10111111", -- 3794 - 0xed2  :  191 - 0xbf
    "11111111", -- 3795 - 0xed3  :  255 - 0xff
    "11111111", -- 3796 - 0xed4  :  255 - 0xff
    "11111111", -- 3797 - 0xed5  :  255 - 0xff
    "11111111", -- 3798 - 0xed6  :  255 - 0xff
    "11111111", -- 3799 - 0xed7  :  255 - 0xff
    "11111000", -- 3800 - 0xed8  :  248 - 0xf8 -- plane 1
    "11111111", -- 3801 - 0xed9  :  255 - 0xff
    "11111111", -- 3802 - 0xeda  :  255 - 0xff
    "11111111", -- 3803 - 0xedb  :  255 - 0xff
    "11111111", -- 3804 - 0xedc  :  255 - 0xff
    "11111111", -- 3805 - 0xedd  :  255 - 0xff
    "11111111", -- 3806 - 0xede  :  255 - 0xff
    "11111111", -- 3807 - 0xedf  :  255 - 0xff
    "01111110", -- 3808 - 0xee0  :  126 - 0x7e -- Background 0xee
    "00011110", -- 3809 - 0xee1  :   30 - 0x1e
    "00011110", -- 3810 - 0xee2  :   30 - 0x1e
    "00001110", -- 3811 - 0xee3  :   14 - 0xe
    "00001111", -- 3812 - 0xee4  :   15 - 0xf
    "00011110", -- 3813 - 0xee5  :   30 - 0x1e
    "00011110", -- 3814 - 0xee6  :   30 - 0x1e
    "00111110", -- 3815 - 0xee7  :   62 - 0x3e
    "11111111", -- 3816 - 0xee8  :  255 - 0xff -- plane 1
    "01111111", -- 3817 - 0xee9  :  127 - 0x7f
    "00011111", -- 3818 - 0xeea  :   31 - 0x1f
    "00001111", -- 3819 - 0xeeb  :   15 - 0xf
    "00001111", -- 3820 - 0xeec  :   15 - 0xf
    "10011111", -- 3821 - 0xeed  :  159 - 0x9f
    "10011111", -- 3822 - 0xeee  :  159 - 0x9f
    "10111111", -- 3823 - 0xeef  :  191 - 0xbf
    "01111111", -- 3824 - 0xef0  :  127 - 0x7f -- Background 0xef
    "01111111", -- 3825 - 0xef1  :  127 - 0x7f
    "10111111", -- 3826 - 0xef2  :  191 - 0xbf
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11111111", -- 3828 - 0xef4  :  255 - 0xff
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11100111", -- 3830 - 0xef6  :  231 - 0xe7
    "11000000", -- 3831 - 0xef7  :  192 - 0xc0
    "01111111", -- 3832 - 0xef8  :  127 - 0x7f -- plane 1
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "11111111", -- 3834 - 0xefa  :  255 - 0xff
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111111", -- 3836 - 0xefc  :  255 - 0xff
    "11111111", -- 3837 - 0xefd  :  255 - 0xff
    "11111111", -- 3838 - 0xefe  :  255 - 0xff
    "11001111", -- 3839 - 0xeff  :  207 - 0xcf
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00010000", -- 3842 - 0xf02  :   16 - 0x10
    "11111101", -- 3843 - 0xf03  :  253 - 0xfd
    "11111010", -- 3844 - 0xf04  :  250 - 0xfa
    "11101011", -- 3845 - 0xf05  :  235 - 0xeb
    "10000000", -- 3846 - 0xf06  :  128 - 0x80
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- plane 1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "11110000", -- 3850 - 0xf0a  :  240 - 0xf0
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "00100000", -- 3856 - 0xf10  :   32 - 0x20 -- Background 0xf1
    "00011111", -- 3857 - 0xf11  :   31 - 0x1f
    "01100000", -- 3858 - 0xf12  :   96 - 0x60
    "10001110", -- 3859 - 0xf13  :  142 - 0x8e
    "00111111", -- 3860 - 0xf14  :   63 - 0x3f
    "01111111", -- 3861 - 0xf15  :  127 - 0x7f
    "01111111", -- 3862 - 0xf16  :  127 - 0x7f
    "01111100", -- 3863 - 0xf17  :  124 - 0x7c
    "11111111", -- 3864 - 0xf18  :  255 - 0xff -- plane 1
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11110001", -- 3867 - 0xf1b  :  241 - 0xf1
    "11000100", -- 3868 - 0xf1c  :  196 - 0xc4
    "11101110", -- 3869 - 0xf1d  :  238 - 0xee
    "11000100", -- 3870 - 0xf1e  :  196 - 0xc4
    "10000011", -- 3871 - 0xf1f  :  131 - 0x83
    "00111001", -- 3872 - 0xf20  :   57 - 0x39 -- Background 0xf2
    "00110110", -- 3873 - 0xf21  :   54 - 0x36
    "00101110", -- 3874 - 0xf22  :   46 - 0x2e
    "10101111", -- 3875 - 0xf23  :  175 - 0xaf
    "10101110", -- 3876 - 0xf24  :  174 - 0xae
    "11010001", -- 3877 - 0xf25  :  209 - 0xd1
    "11101111", -- 3878 - 0xf26  :  239 - 0xef
    "10000111", -- 3879 - 0xf27  :  135 - 0x87
    "11000111", -- 3880 - 0xf28  :  199 - 0xc7 -- plane 1
    "11111001", -- 3881 - 0xf29  :  249 - 0xf9
    "11110000", -- 3882 - 0xf2a  :  240 - 0xf0
    "11110000", -- 3883 - 0xf2b  :  240 - 0xf0
    "10110001", -- 3884 - 0xf2c  :  177 - 0xb1
    "11011111", -- 3885 - 0xf2d  :  223 - 0xdf
    "11101111", -- 3886 - 0xf2e  :  239 - 0xef
    "10000111", -- 3887 - 0xf2f  :  135 - 0x87
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000100", -- 3890 - 0xf32  :    4 - 0x4
    "01011111", -- 3891 - 0xf33  :   95 - 0x5f
    "10101111", -- 3892 - 0xf34  :  175 - 0xaf
    "01010011", -- 3893 - 0xf35  :   83 - 0x53
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000000", -- 3896 - 0xf38  :    0 - 0x0 -- plane 1
    "00000000", -- 3897 - 0xf39  :    0 - 0x0
    "00000111", -- 3898 - 0xf3a  :    7 - 0x7
    "11111111", -- 3899 - 0xf3b  :  255 - 0xff
    "11111111", -- 3900 - 0xf3c  :  255 - 0xff
    "11111111", -- 3901 - 0xf3d  :  255 - 0xff
    "11111111", -- 3902 - 0xf3e  :  255 - 0xff
    "11111111", -- 3903 - 0xf3f  :  255 - 0xff
    "00000010", -- 3904 - 0xf40  :    2 - 0x2 -- Background 0xf4
    "11111100", -- 3905 - 0xf41  :  252 - 0xfc
    "00000011", -- 3906 - 0xf42  :    3 - 0x3
    "00111000", -- 3907 - 0xf43  :   56 - 0x38
    "11111110", -- 3908 - 0xf44  :  254 - 0xfe
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "00011110", -- 3911 - 0xf47  :   30 - 0x1e
    "11111111", -- 3912 - 0xf48  :  255 - 0xff -- plane 1
    "11111111", -- 3913 - 0xf49  :  255 - 0xff
    "11111111", -- 3914 - 0xf4a  :  255 - 0xff
    "11000111", -- 3915 - 0xf4b  :  199 - 0xc7
    "01000101", -- 3916 - 0xf4c  :   69 - 0x45
    "11101110", -- 3917 - 0xf4d  :  238 - 0xee
    "01000100", -- 3918 - 0xf4e  :   68 - 0x44
    "11100001", -- 3919 - 0xf4f  :  225 - 0xe1
    "11000000", -- 3920 - 0xf50  :  192 - 0xc0 -- Background 0xf5
    "00110110", -- 3921 - 0xf51  :   54 - 0x36
    "00111110", -- 3922 - 0xf52  :   62 - 0x3e
    "01111010", -- 3923 - 0xf53  :  122 - 0x7a
    "10110110", -- 3924 - 0xf54  :  182 - 0xb6
    "11001101", -- 3925 - 0xf55  :  205 - 0xcd
    "11111011", -- 3926 - 0xf56  :  251 - 0xfb
    "11110000", -- 3927 - 0xf57  :  240 - 0xf0
    "11111111", -- 3928 - 0xf58  :  255 - 0xff -- plane 1
    "11001111", -- 3929 - 0xf59  :  207 - 0xcf
    "10000111", -- 3930 - 0xf5a  :  135 - 0x87
    "10000111", -- 3931 - 0xf5b  :  135 - 0x87
    "11001110", -- 3932 - 0xf5c  :  206 - 0xce
    "11111101", -- 3933 - 0xf5d  :  253 - 0xfd
    "11111011", -- 3934 - 0xf5e  :  251 - 0xfb
    "11110000", -- 3935 - 0xf5f  :  240 - 0xf0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00001110", -- 3941 - 0xf65  :   14 - 0xe
    "00001000", -- 3942 - 0xf66  :    8 - 0x8
    "00001000", -- 3943 - 0xf67  :    8 - 0x8
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- plane 1
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000001", -- 3949 - 0xf6d  :    1 - 0x1
    "00000111", -- 3950 - 0xf6e  :    7 - 0x7
    "00001111", -- 3951 - 0xf6f  :   15 - 0xf
    "00011111", -- 3952 - 0xf70  :   31 - 0x1f -- Background 0xf7
    "00111111", -- 3953 - 0xf71  :   63 - 0x3f
    "11111111", -- 3954 - 0xf72  :  255 - 0xff
    "11111111", -- 3955 - 0xf73  :  255 - 0xff
    "11111111", -- 3956 - 0xf74  :  255 - 0xff
    "11111111", -- 3957 - 0xf75  :  255 - 0xff
    "11111111", -- 3958 - 0xf76  :  255 - 0xff
    "01111111", -- 3959 - 0xf77  :  127 - 0x7f
    "00111111", -- 3960 - 0xf78  :   63 - 0x3f -- plane 1
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "00111111", -- 3968 - 0xf80  :   63 - 0x3f -- Background 0xf8
    "00111110", -- 3969 - 0xf81  :   62 - 0x3e
    "00111100", -- 3970 - 0xf82  :   60 - 0x3c
    "10111000", -- 3971 - 0xf83  :  184 - 0xb8
    "01111000", -- 3972 - 0xf84  :  120 - 0x78
    "01111000", -- 3973 - 0xf85  :  120 - 0x78
    "01111110", -- 3974 - 0xf86  :  126 - 0x7e
    "01111110", -- 3975 - 0xf87  :  126 - 0x7e
    "11111111", -- 3976 - 0xf88  :  255 - 0xff -- plane 1
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111101", -- 3978 - 0xf8a  :  253 - 0xfd
    "11111000", -- 3979 - 0xf8b  :  248 - 0xf8
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111110", -- 3982 - 0xf8e  :  254 - 0xfe
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111101", -- 3984 - 0xf90  :  253 - 0xfd -- Background 0xf9
    "01111001", -- 3985 - 0xf91  :  121 - 0x79
    "01111011", -- 3986 - 0xf92  :  123 - 0x7b
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11110011", -- 3990 - 0xf96  :  243 - 0xf3
    "10000000", -- 3991 - 0xf97  :  128 - 0x80
    "11111111", -- 3992 - 0xf98  :  255 - 0xff -- plane 1
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111000", -- 3999 - 0xf9f  :  248 - 0xf8
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- plane 1
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "11000000", -- 4014 - 0xfae  :  192 - 0xc0
    "11110000", -- 4015 - 0xfaf  :  240 - 0xf0
    "00010000", -- 4016 - 0xfb0  :   16 - 0x10 -- Background 0xfb
    "10000100", -- 4017 - 0xfb1  :  132 - 0x84
    "11100000", -- 4018 - 0xfb2  :  224 - 0xe0
    "11000000", -- 4019 - 0xfb3  :  192 - 0xc0
    "10000000", -- 4020 - 0xfb4  :  128 - 0x80
    "10000000", -- 4021 - 0xfb5  :  128 - 0x80
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "11111100", -- 4024 - 0xfb8  :  252 - 0xfc -- plane 1
    "11111110", -- 4025 - 0xfb9  :  254 - 0xfe
    "11101100", -- 4026 - 0xfba  :  236 - 0xec
    "11100000", -- 4027 - 0xfbb  :  224 - 0xe0
    "11000000", -- 4028 - 0xfbc  :  192 - 0xc0
    "11000000", -- 4029 - 0xfbd  :  192 - 0xc0
    "10000000", -- 4030 - 0xfbe  :  128 - 0x80
    "10000000", -- 4031 - 0xfbf  :  128 - 0x80
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Background 0xfc
    "01001000", -- 4033 - 0xfc1  :   72 - 0x48
    "00100000", -- 4034 - 0xfc2  :   32 - 0x20
    "00000000", -- 4035 - 0xfc3  :    0 - 0x0
    "00000000", -- 4036 - 0xfc4  :    0 - 0x0
    "00000100", -- 4037 - 0xfc5  :    4 - 0x4
    "00001110", -- 4038 - 0xfc6  :   14 - 0xe
    "11111110", -- 4039 - 0xfc7  :  254 - 0xfe
    "01110000", -- 4040 - 0xfc8  :  112 - 0x70 -- plane 1
    "11111100", -- 4041 - 0xfc9  :  252 - 0xfc
    "11111100", -- 4042 - 0xfca  :  252 - 0xfc
    "11111100", -- 4043 - 0xfcb  :  252 - 0xfc
    "11111100", -- 4044 - 0xfcc  :  252 - 0xfc
    "11111100", -- 4045 - 0xfcd  :  252 - 0xfc
    "11111110", -- 4046 - 0xfce  :  254 - 0xfe
    "11111110", -- 4047 - 0xfcf  :  254 - 0xfe
    "11111110", -- 4048 - 0xfd0  :  254 - 0xfe -- Background 0xfd
    "11111100", -- 4049 - 0xfd1  :  252 - 0xfc
    "11111100", -- 4050 - 0xfd2  :  252 - 0xfc
    "11111000", -- 4051 - 0xfd3  :  248 - 0xf8
    "11110000", -- 4052 - 0xfd4  :  240 - 0xf0
    "11100000", -- 4053 - 0xfd5  :  224 - 0xe0
    "10000000", -- 4054 - 0xfd6  :  128 - 0x80
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "11111110", -- 4056 - 0xfd8  :  254 - 0xfe -- plane 1
    "11111100", -- 4057 - 0xfd9  :  252 - 0xfc
    "11111100", -- 4058 - 0xfda  :  252 - 0xfc
    "11111000", -- 4059 - 0xfdb  :  248 - 0xf8
    "11110000", -- 4060 - 0xfdc  :  240 - 0xf0
    "11100000", -- 4061 - 0xfdd  :  224 - 0xe0
    "10000000", -- 4062 - 0xfde  :  128 - 0x80
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00001111", -- 4064 - 0xfe0  :   15 - 0xf -- Background 0xfe
    "00000110", -- 4065 - 0xfe1  :    6 - 0x6
    "00000110", -- 4066 - 0xfe2  :    6 - 0x6
    "00000110", -- 4067 - 0xfe3  :    6 - 0x6
    "00000110", -- 4068 - 0xfe4  :    6 - 0x6
    "00000110", -- 4069 - 0xfe5  :    6 - 0x6
    "00001111", -- 4070 - 0xfe6  :   15 - 0xf
    "00000000", -- 4071 - 0xfe7  :    0 - 0x0
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- plane 1
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "00000000", -- 4075 - 0xfeb  :    0 - 0x0
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "11110000", -- 4080 - 0xff0  :  240 - 0xf0 -- Background 0xff
    "01100000", -- 4081 - 0xff1  :   96 - 0x60
    "01100000", -- 4082 - 0xff2  :   96 - 0x60
    "01100110", -- 4083 - 0xff3  :  102 - 0x66
    "01100110", -- 4084 - 0xff4  :  102 - 0x66
    "01100000", -- 4085 - 0xff5  :   96 - 0x60
    "11110000", -- 4086 - 0xff6  :  240 - 0xf0
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- plane 1
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
