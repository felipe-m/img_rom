---   Sprites Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG_SPR is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG_SPR;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG_SPR is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table both color planes
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000011", --    1 -  0x1  :    3 - 0x3
    "00000111", --    2 -  0x2  :    7 - 0x7
    "00000111", --    3 -  0x3  :    7 - 0x7
    "00001001", --    4 -  0x4  :    9 - 0x9
    "00001001", --    5 -  0x5  :    9 - 0x9
    "00011100", --    6 -  0x6  :   28 - 0x1c
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000011", --    9 -  0x9  :    3 - 0x3
    "00000111", --   10 -  0xa  :    7 - 0x7
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000110", --   12 -  0xc  :    6 - 0x6
    "00000110", --   13 -  0xd  :    6 - 0x6
    "00000011", --   14 -  0xe  :    3 - 0x3
    "00000011", --   15 -  0xf  :    3 - 0x3
    "00001111", --   16 - 0x10  :   15 - 0xf -- Sprite 0x1
    "00001111", --   17 - 0x11  :   15 - 0xf
    "00001111", --   18 - 0x12  :   15 - 0xf
    "11111111", --   19 - 0x13  :  255 - 0xff
    "11111111", --   20 - 0x14  :  255 - 0xff
    "11111100", --   21 - 0x15  :  252 - 0xfc
    "10000001", --   22 - 0x16  :  129 - 0x81
    "00000001", --   23 - 0x17  :    1 - 0x1
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00010000", --   25 - 0x19  :   16 - 0x10
    "00111100", --   26 - 0x1a  :   60 - 0x3c
    "00111111", --   27 - 0x1b  :   63 - 0x3f
    "00111111", --   28 - 0x1c  :   63 - 0x3f
    "00111100", --   29 - 0x1d  :   60 - 0x3c
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "11000000", --   33 - 0x21  :  192 - 0xc0
    "11111000", --   34 - 0x22  :  248 - 0xf8
    "10000000", --   35 - 0x23  :  128 - 0x80
    "00100000", --   36 - 0x24  :   32 - 0x20
    "10010000", --   37 - 0x25  :  144 - 0x90
    "00111100", --   38 - 0x26  :   60 - 0x3c
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "11000000", --   41 - 0x29  :  192 - 0xc0
    "11111000", --   42 - 0x2a  :  248 - 0xf8
    "01100000", --   43 - 0x2b  :   96 - 0x60
    "11011100", --   44 - 0x2c  :  220 - 0xdc
    "01101110", --   45 - 0x2d  :  110 - 0x6e
    "11000000", --   46 - 0x2e  :  192 - 0xc0
    "11111000", --   47 - 0x2f  :  248 - 0xf8
    "11000000", --   48 - 0x30  :  192 - 0xc0 -- Sprite 0x3
    "11000000", --   49 - 0x31  :  192 - 0xc0
    "11000000", --   50 - 0x32  :  192 - 0xc0
    "11110000", --   51 - 0x33  :  240 - 0xf0
    "11110000", --   52 - 0x34  :  240 - 0xf0
    "11100000", --   53 - 0x35  :  224 - 0xe0
    "11000000", --   54 - 0x36  :  192 - 0xc0
    "11100000", --   55 - 0x37  :  224 - 0xe0
    "01010000", --   56 - 0x38  :   80 - 0x50 -- plane 1
    "00111000", --   57 - 0x39  :   56 - 0x38
    "00110000", --   58 - 0x3a  :   48 - 0x30
    "11110000", --   59 - 0x3b  :  240 - 0xf0
    "11110000", --   60 - 0x3c  :  240 - 0xf0
    "11100000", --   61 - 0x3d  :  224 - 0xe0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000111", --   64 - 0x40  :    7 - 0x7 -- Sprite 0x4
    "00001111", --   65 - 0x41  :   15 - 0xf
    "00001111", --   66 - 0x42  :   15 - 0xf
    "00010010", --   67 - 0x43  :   18 - 0x12
    "00010011", --   68 - 0x44  :   19 - 0x13
    "00111000", --   69 - 0x45  :   56 - 0x38
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00001111", --   71 - 0x47  :   15 - 0xf
    "00000111", --   72 - 0x48  :    7 - 0x7 -- plane 1
    "00001111", --   73 - 0x49  :   15 - 0xf
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00001101", --   75 - 0x4b  :   13 - 0xd
    "00001100", --   76 - 0x4c  :   12 - 0xc
    "00000111", --   77 - 0x4d  :    7 - 0x7
    "00000111", --   78 - 0x4e  :    7 - 0x7
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00011111", --   80 - 0x50  :   31 - 0x1f -- Sprite 0x5
    "00011111", --   81 - 0x51  :   31 - 0x1f
    "00011111", --   82 - 0x52  :   31 - 0x1f
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00011001", --   84 - 0x54  :   25 - 0x19
    "00011110", --   85 - 0x55  :   30 - 0x1e
    "00011100", --   86 - 0x56  :   28 - 0x1c
    "00011110", --   87 - 0x57  :   30 - 0x1e
    "00000001", --   88 - 0x58  :    1 - 0x1 -- plane 1
    "00000011", --   89 - 0x59  :    3 - 0x3
    "00000001", --   90 - 0x5a  :    1 - 0x1
    "00010111", --   91 - 0x5b  :   23 - 0x17
    "00011111", --   92 - 0x5c  :   31 - 0x1f
    "00011110", --   93 - 0x5d  :   30 - 0x1e
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "10000000", --   96 - 0x60  :  128 - 0x80 -- Sprite 0x6
    "11110000", --   97 - 0x61  :  240 - 0xf0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "01000000", --   99 - 0x63  :   64 - 0x40
    "00100000", --  100 - 0x64  :   32 - 0x20
    "01111000", --  101 - 0x65  :  120 - 0x78
    "00000000", --  102 - 0x66  :    0 - 0x0
    "11000000", --  103 - 0x67  :  192 - 0xc0
    "10000000", --  104 - 0x68  :  128 - 0x80 -- plane 1
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11000000", --  106 - 0x6a  :  192 - 0xc0
    "10111000", --  107 - 0x6b  :  184 - 0xb8
    "11011100", --  108 - 0x6c  :  220 - 0xdc
    "10000000", --  109 - 0x6d  :  128 - 0x80
    "11110000", --  110 - 0x6e  :  240 - 0xf0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11100000", --  112 - 0x70  :  224 - 0xe0 -- Sprite 0x7
    "01100000", --  113 - 0x71  :   96 - 0x60
    "11110000", --  114 - 0x72  :  240 - 0xf0
    "11110000", --  115 - 0x73  :  240 - 0xf0
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11100000", --  117 - 0x75  :  224 - 0xe0
    "11100000", --  118 - 0x76  :  224 - 0xe0
    "11110000", --  119 - 0x77  :  240 - 0xf0
    "10000000", --  120 - 0x78  :  128 - 0x80 -- plane 1
    "11100000", --  121 - 0x79  :  224 - 0xe0
    "11110000", --  122 - 0x7a  :  240 - 0xf0
    "11110000", --  123 - 0x7b  :  240 - 0xf0
    "11110000", --  124 - 0x7c  :  240 - 0xf0
    "11100000", --  125 - 0x7d  :  224 - 0xe0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000111", --  128 - 0x80  :    7 - 0x7 -- Sprite 0x8
    "00001111", --  129 - 0x81  :   15 - 0xf
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00010010", --  131 - 0x83  :   18 - 0x12
    "00010011", --  132 - 0x84  :   19 - 0x13
    "00111000", --  133 - 0x85  :   56 - 0x38
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00000111", --  136 - 0x88  :    7 - 0x7 -- plane 1
    "00001111", --  137 - 0x89  :   15 - 0xf
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00001101", --  139 - 0x8b  :   13 - 0xd
    "00001100", --  140 - 0x8c  :   12 - 0xc
    "00000111", --  141 - 0x8d  :    7 - 0x7
    "00000111", --  142 - 0x8e  :    7 - 0x7
    "00000011", --  143 - 0x8f  :    3 - 0x3
    "00111111", --  144 - 0x90  :   63 - 0x3f -- Sprite 0x9
    "00001110", --  145 - 0x91  :   14 - 0xe
    "00001111", --  146 - 0x92  :   15 - 0xf
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00111111", --  148 - 0x94  :   63 - 0x3f
    "01111100", --  149 - 0x95  :  124 - 0x7c
    "01110000", --  150 - 0x96  :  112 - 0x70
    "00111000", --  151 - 0x97  :   56 - 0x38
    "11000011", --  152 - 0x98  :  195 - 0xc3 -- plane 1
    "11100011", --  153 - 0x99  :  227 - 0xe3
    "11001111", --  154 - 0x9a  :  207 - 0xcf
    "00011111", --  155 - 0x9b  :   31 - 0x1f
    "00111111", --  156 - 0x9c  :   63 - 0x3f
    "00001100", --  157 - 0x9d  :   12 - 0xc
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "10000000", --  160 - 0xa0  :  128 - 0x80 -- Sprite 0xa
    "11110000", --  161 - 0xa1  :  240 - 0xf0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "01000000", --  163 - 0xa3  :   64 - 0x40
    "00100000", --  164 - 0xa4  :   32 - 0x20
    "01111000", --  165 - 0xa5  :  120 - 0x78
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "11000000", --  167 - 0xa7  :  192 - 0xc0
    "10000000", --  168 - 0xa8  :  128 - 0x80 -- plane 1
    "11110000", --  169 - 0xa9  :  240 - 0xf0
    "11000000", --  170 - 0xaa  :  192 - 0xc0
    "10111000", --  171 - 0xab  :  184 - 0xb8
    "11011100", --  172 - 0xac  :  220 - 0xdc
    "10000000", --  173 - 0xad  :  128 - 0x80
    "11110000", --  174 - 0xae  :  240 - 0xf0
    "00000110", --  175 - 0xaf  :    6 - 0x6
    "11110000", --  176 - 0xb0  :  240 - 0xf0 -- Sprite 0xb
    "11111000", --  177 - 0xb1  :  248 - 0xf8
    "11100100", --  178 - 0xb2  :  228 - 0xe4
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11111100", --  180 - 0xb4  :  252 - 0xfc
    "01111100", --  181 - 0xb5  :  124 - 0x7c
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "10001110", --  184 - 0xb8  :  142 - 0x8e -- plane 1
    "11100110", --  185 - 0xb9  :  230 - 0xe6
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "11110000", --  187 - 0xbb  :  240 - 0xf0
    "11110000", --  188 - 0xbc  :  240 - 0xf0
    "01110000", --  189 - 0xbd  :  112 - 0x70
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00000010", --  193 - 0xc1  :    2 - 0x2
    "00000110", --  194 - 0xc2  :    6 - 0x6
    "00000111", --  195 - 0xc3  :    7 - 0x7
    "00001001", --  196 - 0xc4  :    9 - 0x9
    "00001001", --  197 - 0xc5  :    9 - 0x9
    "00011101", --  198 - 0xc6  :   29 - 0x1d
    "00000011", --  199 - 0xc7  :    3 - 0x3
    "00000001", --  200 - 0xc8  :    1 - 0x1 -- plane 1
    "00000011", --  201 - 0xc9  :    3 - 0x3
    "00000111", --  202 - 0xca  :    7 - 0x7
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000110", --  204 - 0xcc  :    6 - 0x6
    "00000110", --  205 - 0xcd  :    6 - 0x6
    "00000010", --  206 - 0xce  :    2 - 0x2
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00001111", --  208 - 0xd0  :   15 - 0xf -- Sprite 0xd
    "00001111", --  209 - 0xd1  :   15 - 0xf
    "00001111", --  210 - 0xd2  :   15 - 0xf
    "11111111", --  211 - 0xd3  :  255 - 0xff
    "11111111", --  212 - 0xd4  :  255 - 0xff
    "11111100", --  213 - 0xd5  :  252 - 0xfc
    "10000001", --  214 - 0xd6  :  129 - 0x81
    "00000001", --  215 - 0xd7  :    1 - 0x1
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- plane 1
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00001100", --  218 - 0xda  :   12 - 0xc
    "00111111", --  219 - 0xdb  :   63 - 0x3f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00111100", --  221 - 0xdd  :   60 - 0x3c
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00111000", --  226 - 0xe2  :   56 - 0x38
    "11000000", --  227 - 0xe3  :  192 - 0xc0
    "11100000", --  228 - 0xe4  :  224 - 0xe0
    "11010000", --  229 - 0xe5  :  208 - 0xd0
    "11111100", --  230 - 0xe6  :  252 - 0xfc
    "11000000", --  231 - 0xe7  :  192 - 0xc0
    "11000000", --  232 - 0xe8  :  192 - 0xc0 -- plane 1
    "11000000", --  233 - 0xe9  :  192 - 0xc0
    "11111000", --  234 - 0xea  :  248 - 0xf8
    "00100000", --  235 - 0xeb  :   32 - 0x20
    "00011100", --  236 - 0xec  :   28 - 0x1c
    "00101110", --  237 - 0xed  :   46 - 0x2e
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00111000", --  239 - 0xef  :   56 - 0x38
    "11100000", --  240 - 0xf0  :  224 - 0xe0 -- Sprite 0xf
    "11100000", --  241 - 0xf1  :  224 - 0xe0
    "10110000", --  242 - 0xf2  :  176 - 0xb0
    "11110000", --  243 - 0xf3  :  240 - 0xf0
    "11110000", --  244 - 0xf4  :  240 - 0xf0
    "11100000", --  245 - 0xf5  :  224 - 0xe0
    "11000000", --  246 - 0xf6  :  192 - 0xc0
    "11100000", --  247 - 0xf7  :  224 - 0xe0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- plane 1
    "01100000", --  249 - 0xf9  :   96 - 0x60
    "11110000", --  250 - 0xfa  :  240 - 0xf0
    "11110000", --  251 - 0xfb  :  240 - 0xf0
    "11110000", --  252 - 0xfc  :  240 - 0xf0
    "11100000", --  253 - 0xfd  :  224 - 0xe0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  257 - 0x101  :    3 - 0x3
    "00000111", --  258 - 0x102  :    7 - 0x7
    "00000111", --  259 - 0x103  :    7 - 0x7
    "00001001", --  260 - 0x104  :    9 - 0x9
    "00001001", --  261 - 0x105  :    9 - 0x9
    "00011100", --  262 - 0x106  :   28 - 0x1c
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- plane 1
    "00000011", --  265 - 0x109  :    3 - 0x3
    "00000111", --  266 - 0x10a  :    7 - 0x7
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000110", --  268 - 0x10c  :    6 - 0x6
    "00000110", --  269 - 0x10d  :    6 - 0x6
    "00000011", --  270 - 0x10e  :    3 - 0x3
    "00000011", --  271 - 0x10f  :    3 - 0x3
    "00001111", --  272 - 0x110  :   15 - 0xf -- Sprite 0x11
    "00001111", --  273 - 0x111  :   15 - 0xf
    "00001111", --  274 - 0x112  :   15 - 0xf
    "11111111", --  275 - 0x113  :  255 - 0xff
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111100", --  277 - 0x115  :  252 - 0xfc
    "10000001", --  278 - 0x116  :  129 - 0x81
    "00000001", --  279 - 0x117  :    1 - 0x1
    "00000000", --  280 - 0x118  :    0 - 0x0 -- plane 1
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00001100", --  282 - 0x11a  :   12 - 0xc
    "00111111", --  283 - 0x11b  :   63 - 0x3f
    "00111111", --  284 - 0x11c  :   63 - 0x3f
    "00111100", --  285 - 0x11d  :   60 - 0x3c
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x12
    "11000000", --  289 - 0x121  :  192 - 0xc0
    "11111000", --  290 - 0x122  :  248 - 0xf8
    "10000000", --  291 - 0x123  :  128 - 0x80
    "00100000", --  292 - 0x124  :   32 - 0x20
    "10010000", --  293 - 0x125  :  144 - 0x90
    "00111100", --  294 - 0x126  :   60 - 0x3c
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- plane 1
    "11000000", --  297 - 0x129  :  192 - 0xc0
    "11111000", --  298 - 0x12a  :  248 - 0xf8
    "01100000", --  299 - 0x12b  :   96 - 0x60
    "11011100", --  300 - 0x12c  :  220 - 0xdc
    "01101110", --  301 - 0x12d  :  110 - 0x6e
    "11000000", --  302 - 0x12e  :  192 - 0xc0
    "11111000", --  303 - 0x12f  :  248 - 0xf8
    "11100000", --  304 - 0x130  :  224 - 0xe0 -- Sprite 0x13
    "11110000", --  305 - 0x131  :  240 - 0xf0
    "11110000", --  306 - 0x132  :  240 - 0xf0
    "11110000", --  307 - 0x133  :  240 - 0xf0
    "11110000", --  308 - 0x134  :  240 - 0xf0
    "11100000", --  309 - 0x135  :  224 - 0xe0
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "11100000", --  311 - 0x137  :  224 - 0xe0
    "01000111", --  312 - 0x138  :   71 - 0x47 -- plane 1
    "00001111", --  313 - 0x139  :   15 - 0xf
    "00001110", --  314 - 0x13a  :   14 - 0xe
    "11110000", --  315 - 0x13b  :  240 - 0xf0
    "11110000", --  316 - 0x13c  :  240 - 0xf0
    "11100000", --  317 - 0x13d  :  224 - 0xe0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000100", --  320 - 0x140  :    4 - 0x4 -- Sprite 0x14
    "00001100", --  321 - 0x141  :   12 - 0xc
    "00001100", --  322 - 0x142  :   12 - 0xc
    "00010011", --  323 - 0x143  :   19 - 0x13
    "00010011", --  324 - 0x144  :   19 - 0x13
    "00111011", --  325 - 0x145  :   59 - 0x3b
    "00000111", --  326 - 0x146  :    7 - 0x7
    "00001111", --  327 - 0x147  :   15 - 0xf
    "00000111", --  328 - 0x148  :    7 - 0x7 -- plane 1
    "00001111", --  329 - 0x149  :   15 - 0xf
    "00000011", --  330 - 0x14a  :    3 - 0x3
    "00001100", --  331 - 0x14b  :   12 - 0xc
    "00001100", --  332 - 0x14c  :   12 - 0xc
    "00000100", --  333 - 0x14d  :    4 - 0x4
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00001111", --  336 - 0x150  :   15 - 0xf -- Sprite 0x15
    "00001111", --  337 - 0x151  :   15 - 0xf
    "00001111", --  338 - 0x152  :   15 - 0xf
    "00011111", --  339 - 0x153  :   31 - 0x1f
    "00011111", --  340 - 0x154  :   31 - 0x1f
    "00011110", --  341 - 0x155  :   30 - 0x1e
    "00011100", --  342 - 0x156  :   28 - 0x1c
    "00011110", --  343 - 0x157  :   30 - 0x1e
    "00000000", --  344 - 0x158  :    0 - 0x0 -- plane 1
    "00000001", --  345 - 0x159  :    1 - 0x1
    "00001111", --  346 - 0x15a  :   15 - 0xf
    "00011111", --  347 - 0x15b  :   31 - 0x1f
    "00011111", --  348 - 0x15c  :   31 - 0x1f
    "00011110", --  349 - 0x15d  :   30 - 0x1e
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x16
    "01110000", --  353 - 0x161  :  112 - 0x70
    "00000000", --  354 - 0x162  :    0 - 0x0
    "11000000", --  355 - 0x163  :  192 - 0xc0
    "10100000", --  356 - 0x164  :  160 - 0xa0
    "11111000", --  357 - 0x165  :  248 - 0xf8
    "10000000", --  358 - 0x166  :  128 - 0x80
    "11000000", --  359 - 0x167  :  192 - 0xc0
    "10000000", --  360 - 0x168  :  128 - 0x80 -- plane 1
    "11110000", --  361 - 0x169  :  240 - 0xf0
    "11000000", --  362 - 0x16a  :  192 - 0xc0
    "00111000", --  363 - 0x16b  :   56 - 0x38
    "01011100", --  364 - 0x16c  :   92 - 0x5c
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "01110000", --  366 - 0x16e  :  112 - 0x70
    "01000000", --  367 - 0x16f  :   64 - 0x40
    "11100000", --  368 - 0x170  :  224 - 0xe0 -- Sprite 0x17
    "01100000", --  369 - 0x171  :   96 - 0x60
    "11110000", --  370 - 0x172  :  240 - 0xf0
    "11110000", --  371 - 0x173  :  240 - 0xf0
    "11110000", --  372 - 0x174  :  240 - 0xf0
    "11100000", --  373 - 0x175  :  224 - 0xe0
    "11100000", --  374 - 0x176  :  224 - 0xe0
    "11110000", --  375 - 0x177  :  240 - 0xf0
    "11000000", --  376 - 0x178  :  192 - 0xc0 -- plane 1
    "11100000", --  377 - 0x179  :  224 - 0xe0
    "11110000", --  378 - 0x17a  :  240 - 0xf0
    "11110000", --  379 - 0x17b  :  240 - 0xf0
    "11110000", --  380 - 0x17c  :  240 - 0xf0
    "11100000", --  381 - 0x17d  :  224 - 0xe0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000111", --  384 - 0x180  :    7 - 0x7 -- Sprite 0x18
    "00001111", --  385 - 0x181  :   15 - 0xf
    "00001111", --  386 - 0x182  :   15 - 0xf
    "00010010", --  387 - 0x183  :   18 - 0x12
    "00010011", --  388 - 0x184  :   19 - 0x13
    "00111000", --  389 - 0x185  :   56 - 0x38
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00001111", --  391 - 0x187  :   15 - 0xf
    "00000111", --  392 - 0x188  :    7 - 0x7 -- plane 1
    "00001111", --  393 - 0x189  :   15 - 0xf
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00001101", --  395 - 0x18b  :   13 - 0xd
    "00001100", --  396 - 0x18c  :   12 - 0xc
    "00000111", --  397 - 0x18d  :    7 - 0x7
    "00000111", --  398 - 0x18e  :    7 - 0x7
    "00000001", --  399 - 0x18f  :    1 - 0x1
    "00011111", --  400 - 0x190  :   31 - 0x1f -- Sprite 0x19
    "00011111", --  401 - 0x191  :   31 - 0x1f
    "00011111", --  402 - 0x192  :   31 - 0x1f
    "00011111", --  403 - 0x193  :   31 - 0x1f
    "00011111", --  404 - 0x194  :   31 - 0x1f
    "00011110", --  405 - 0x195  :   30 - 0x1e
    "00011100", --  406 - 0x196  :   28 - 0x1c
    "00011110", --  407 - 0x197  :   30 - 0x1e
    "00000000", --  408 - 0x198  :    0 - 0x0 -- plane 1
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00010011", --  410 - 0x19a  :   19 - 0x13
    "00011111", --  411 - 0x19b  :   31 - 0x1f
    "00011111", --  412 - 0x19c  :   31 - 0x1f
    "00011110", --  413 - 0x19d  :   30 - 0x1e
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "10000000", --  416 - 0x1a0  :  128 - 0x80 -- Sprite 0x1a
    "11110000", --  417 - 0x1a1  :  240 - 0xf0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "01000000", --  419 - 0x1a3  :   64 - 0x40
    "00100000", --  420 - 0x1a4  :   32 - 0x20
    "01111000", --  421 - 0x1a5  :  120 - 0x78
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "11000000", --  423 - 0x1a7  :  192 - 0xc0
    "10000000", --  424 - 0x1a8  :  128 - 0x80 -- plane 1
    "11110000", --  425 - 0x1a9  :  240 - 0xf0
    "11000000", --  426 - 0x1aa  :  192 - 0xc0
    "10111000", --  427 - 0x1ab  :  184 - 0xb8
    "11011100", --  428 - 0x1ac  :  220 - 0xdc
    "10000000", --  429 - 0x1ad  :  128 - 0x80
    "11110000", --  430 - 0x1ae  :  240 - 0xf0
    "10000000", --  431 - 0x1af  :  128 - 0x80
    "11111000", --  432 - 0x1b0  :  248 - 0xf8 -- Sprite 0x1b
    "11111000", --  433 - 0x1b1  :  248 - 0xf8
    "11110000", --  434 - 0x1b2  :  240 - 0xf0
    "11110000", --  435 - 0x1b3  :  240 - 0xf0
    "11110000", --  436 - 0x1b4  :  240 - 0xf0
    "11100000", --  437 - 0x1b5  :  224 - 0xe0
    "11100000", --  438 - 0x1b6  :  224 - 0xe0
    "11110000", --  439 - 0x1b7  :  240 - 0xf0
    "00000111", --  440 - 0x1b8  :    7 - 0x7 -- plane 1
    "00000111", --  441 - 0x1b9  :    7 - 0x7
    "11111110", --  442 - 0x1ba  :  254 - 0xfe
    "11110000", --  443 - 0x1bb  :  240 - 0xf0
    "11110000", --  444 - 0x1bc  :  240 - 0xf0
    "11100000", --  445 - 0x1bd  :  224 - 0xe0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000100", --  448 - 0x1c0  :    4 - 0x4 -- Sprite 0x1c
    "00001100", --  449 - 0x1c1  :   12 - 0xc
    "00001100", --  450 - 0x1c2  :   12 - 0xc
    "00010011", --  451 - 0x1c3  :   19 - 0x13
    "00010011", --  452 - 0x1c4  :   19 - 0x13
    "00111111", --  453 - 0x1c5  :   63 - 0x3f
    "00000111", --  454 - 0x1c6  :    7 - 0x7
    "00001111", --  455 - 0x1c7  :   15 - 0xf
    "00000111", --  456 - 0x1c8  :    7 - 0x7 -- plane 1
    "00001111", --  457 - 0x1c9  :   15 - 0xf
    "00000011", --  458 - 0x1ca  :    3 - 0x3
    "00001100", --  459 - 0x1cb  :   12 - 0xc
    "00001100", --  460 - 0x1cc  :   12 - 0xc
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00001111", --  464 - 0x1d0  :   15 - 0xf -- Sprite 0x1d
    "00001111", --  465 - 0x1d1  :   15 - 0xf
    "00001111", --  466 - 0x1d2  :   15 - 0xf
    "00011111", --  467 - 0x1d3  :   31 - 0x1f
    "00111111", --  468 - 0x1d4  :   63 - 0x3f
    "01111100", --  469 - 0x1d5  :  124 - 0x7c
    "01110000", --  470 - 0x1d6  :  112 - 0x70
    "00111000", --  471 - 0x1d7  :   56 - 0x38
    "00000001", --  472 - 0x1d8  :    1 - 0x1 -- plane 1
    "00000001", --  473 - 0x1d9  :    1 - 0x1
    "00001111", --  474 - 0x1da  :   15 - 0xf
    "00011111", --  475 - 0x1db  :   31 - 0x1f
    "00111111", --  476 - 0x1dc  :   63 - 0x3f
    "00011100", --  477 - 0x1dd  :   28 - 0x1c
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x1e
    "01110000", --  481 - 0x1e1  :  112 - 0x70
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "11000000", --  483 - 0x1e3  :  192 - 0xc0
    "10100000", --  484 - 0x1e4  :  160 - 0xa0
    "11111000", --  485 - 0x1e5  :  248 - 0xf8
    "10000000", --  486 - 0x1e6  :  128 - 0x80
    "11000000", --  487 - 0x1e7  :  192 - 0xc0
    "10000000", --  488 - 0x1e8  :  128 - 0x80 -- plane 1
    "11110000", --  489 - 0x1e9  :  240 - 0xf0
    "11000000", --  490 - 0x1ea  :  192 - 0xc0
    "00111000", --  491 - 0x1eb  :   56 - 0x38
    "01011100", --  492 - 0x1ec  :   92 - 0x5c
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "01110000", --  494 - 0x1ee  :  112 - 0x70
    "01000000", --  495 - 0x1ef  :   64 - 0x40
    "11000000", --  496 - 0x1f0  :  192 - 0xc0 -- Sprite 0x1f
    "01100000", --  497 - 0x1f1  :   96 - 0x60
    "11100100", --  498 - 0x1f2  :  228 - 0xe4
    "11111100", --  499 - 0x1f3  :  252 - 0xfc
    "11111100", --  500 - 0x1f4  :  252 - 0xfc
    "01111100", --  501 - 0x1f5  :  124 - 0x7c
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11000000", --  504 - 0x1f8  :  192 - 0xc0 -- plane 1
    "11100000", --  505 - 0x1f9  :  224 - 0xe0
    "11100000", --  506 - 0x1fa  :  224 - 0xe0
    "11110000", --  507 - 0x1fb  :  240 - 0xf0
    "11110000", --  508 - 0x1fc  :  240 - 0xf0
    "01110000", --  509 - 0x1fd  :  112 - 0x70
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000111", --  512 - 0x200  :    7 - 0x7 -- Sprite 0x20
    "00001111", --  513 - 0x201  :   15 - 0xf
    "00001111", --  514 - 0x202  :   15 - 0xf
    "00010010", --  515 - 0x203  :   18 - 0x12
    "00010011", --  516 - 0x204  :   19 - 0x13
    "00111000", --  517 - 0x205  :   56 - 0x38
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000111", --  519 - 0x207  :    7 - 0x7
    "00000111", --  520 - 0x208  :    7 - 0x7 -- plane 1
    "00001111", --  521 - 0x209  :   15 - 0xf
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00001101", --  523 - 0x20b  :   13 - 0xd
    "00001100", --  524 - 0x20c  :   12 - 0xc
    "00000111", --  525 - 0x20d  :    7 - 0x7
    "00000111", --  526 - 0x20e  :    7 - 0x7
    "00000001", --  527 - 0x20f  :    1 - 0x1
    "00001111", --  528 - 0x210  :   15 - 0xf -- Sprite 0x21
    "00001111", --  529 - 0x211  :   15 - 0xf
    "00001111", --  530 - 0x212  :   15 - 0xf
    "00011111", --  531 - 0x213  :   31 - 0x1f
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "01111100", --  533 - 0x215  :  124 - 0x7c
    "01110000", --  534 - 0x216  :  112 - 0x70
    "00111000", --  535 - 0x217  :   56 - 0x38
    "00000000", --  536 - 0x218  :    0 - 0x0 -- plane 1
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00001001", --  538 - 0x21a  :    9 - 0x9
    "00011111", --  539 - 0x21b  :   31 - 0x1f
    "00111111", --  540 - 0x21c  :   63 - 0x3f
    "00011100", --  541 - 0x21d  :   28 - 0x1c
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "10000000", --  544 - 0x220  :  128 - 0x80 -- Sprite 0x22
    "11110000", --  545 - 0x221  :  240 - 0xf0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "01000000", --  547 - 0x223  :   64 - 0x40
    "00100000", --  548 - 0x224  :   32 - 0x20
    "01111000", --  549 - 0x225  :  120 - 0x78
    "00000000", --  550 - 0x226  :    0 - 0x0
    "11000000", --  551 - 0x227  :  192 - 0xc0
    "10000000", --  552 - 0x228  :  128 - 0x80 -- plane 1
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11000000", --  554 - 0x22a  :  192 - 0xc0
    "10111000", --  555 - 0x22b  :  184 - 0xb8
    "11011100", --  556 - 0x22c  :  220 - 0xdc
    "10000000", --  557 - 0x22d  :  128 - 0x80
    "11110000", --  558 - 0x22e  :  240 - 0xf0
    "10000000", --  559 - 0x22f  :  128 - 0x80
    "11111000", --  560 - 0x230  :  248 - 0xf8 -- Sprite 0x23
    "11111000", --  561 - 0x231  :  248 - 0xf8
    "11100000", --  562 - 0x232  :  224 - 0xe0
    "11111100", --  563 - 0x233  :  252 - 0xfc
    "11111100", --  564 - 0x234  :  252 - 0xfc
    "01111100", --  565 - 0x235  :  124 - 0x7c
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000111", --  568 - 0x238  :    7 - 0x7 -- plane 1
    "00000111", --  569 - 0x239  :    7 - 0x7
    "11101110", --  570 - 0x23a  :  238 - 0xee
    "11110000", --  571 - 0x23b  :  240 - 0xf0
    "11110000", --  572 - 0x23c  :  240 - 0xf0
    "01110000", --  573 - 0x23d  :  112 - 0x70
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x24
    "00000111", --  577 - 0x241  :    7 - 0x7
    "00000111", --  578 - 0x242  :    7 - 0x7
    "00001111", --  579 - 0x243  :   15 - 0xf
    "00001111", --  580 - 0x244  :   15 - 0xf
    "00111000", --  581 - 0x245  :   56 - 0x38
    "01111111", --  582 - 0x246  :  127 - 0x7f
    "01111111", --  583 - 0x247  :  127 - 0x7f
    "00000000", --  584 - 0x248  :    0 - 0x0 -- plane 1
    "00000111", --  585 - 0x249  :    7 - 0x7
    "00000011", --  586 - 0x24a  :    3 - 0x3
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000111", --  589 - 0x24d  :    7 - 0x7
    "00000100", --  590 - 0x24e  :    4 - 0x4
    "00000100", --  591 - 0x24f  :    4 - 0x4
    "00011111", --  592 - 0x250  :   31 - 0x1f -- Sprite 0x25
    "00011111", --  593 - 0x251  :   31 - 0x1f
    "00011111", --  594 - 0x252  :   31 - 0x1f
    "00011111", --  595 - 0x253  :   31 - 0x1f
    "00001111", --  596 - 0x254  :   15 - 0xf
    "00001111", --  597 - 0x255  :   15 - 0xf
    "00001111", --  598 - 0x256  :   15 - 0xf
    "00000111", --  599 - 0x257  :    7 - 0x7
    "00011110", --  600 - 0x258  :   30 - 0x1e -- plane 1
    "00011111", --  601 - 0x259  :   31 - 0x1f
    "00011111", --  602 - 0x25a  :   31 - 0x1f
    "00011111", --  603 - 0x25b  :   31 - 0x1f
    "00001111", --  604 - 0x25c  :   15 - 0xf
    "00001000", --  605 - 0x25d  :    8 - 0x8
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x26
    "11100000", --  609 - 0x261  :  224 - 0xe0
    "11111000", --  610 - 0x262  :  248 - 0xf8
    "11111100", --  611 - 0x263  :  252 - 0xfc
    "11111100", --  612 - 0x264  :  252 - 0xfc
    "00011100", --  613 - 0x265  :   28 - 0x1c
    "11111000", --  614 - 0x266  :  248 - 0xf8
    "11111000", --  615 - 0x267  :  248 - 0xf8
    "00111000", --  616 - 0x268  :   56 - 0x38 -- plane 1
    "11111000", --  617 - 0x269  :  248 - 0xf8
    "11000000", --  618 - 0x26a  :  192 - 0xc0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "11100000", --  621 - 0x26d  :  224 - 0xe0
    "00100000", --  622 - 0x26e  :   32 - 0x20
    "00100000", --  623 - 0x26f  :   32 - 0x20
    "11111000", --  624 - 0x270  :  248 - 0xf8 -- Sprite 0x27
    "11111100", --  625 - 0x271  :  252 - 0xfc
    "11111100", --  626 - 0x272  :  252 - 0xfc
    "11111000", --  627 - 0x273  :  248 - 0xf8
    "01111000", --  628 - 0x274  :  120 - 0x78
    "10000000", --  629 - 0x275  :  128 - 0x80
    "11000000", --  630 - 0x276  :  192 - 0xc0
    "11000000", --  631 - 0x277  :  192 - 0xc0
    "01111000", --  632 - 0x278  :  120 - 0x78 -- plane 1
    "11111100", --  633 - 0x279  :  252 - 0xfc
    "11111100", --  634 - 0x27a  :  252 - 0xfc
    "11111000", --  635 - 0x27b  :  248 - 0xf8
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "10000000", --  637 - 0x27d  :  128 - 0x80
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x28
    "00000011", --  641 - 0x281  :    3 - 0x3
    "00000111", --  642 - 0x282  :    7 - 0x7
    "00000111", --  643 - 0x283  :    7 - 0x7
    "00001001", --  644 - 0x284  :    9 - 0x9
    "00001001", --  645 - 0x285  :    9 - 0x9
    "00011100", --  646 - 0x286  :   28 - 0x1c
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00000011", --  649 - 0x289  :    3 - 0x3
    "00000111", --  650 - 0x28a  :    7 - 0x7
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000110", --  652 - 0x28c  :    6 - 0x6
    "00000110", --  653 - 0x28d  :    6 - 0x6
    "00000011", --  654 - 0x28e  :    3 - 0x3
    "01100011", --  655 - 0x28f  :   99 - 0x63
    "00011111", --  656 - 0x290  :   31 - 0x1f -- Sprite 0x29
    "00001111", --  657 - 0x291  :   15 - 0xf
    "00000111", --  658 - 0x292  :    7 - 0x7
    "00110111", --  659 - 0x293  :   55 - 0x37
    "01111111", --  660 - 0x294  :  127 - 0x7f
    "11011111", --  661 - 0x295  :  223 - 0xdf
    "00001111", --  662 - 0x296  :   15 - 0xf
    "00000110", --  663 - 0x297  :    6 - 0x6
    "11100000", --  664 - 0x298  :  224 - 0xe0 -- plane 1
    "00100001", --  665 - 0x299  :   33 - 0x21
    "00000001", --  666 - 0x29a  :    1 - 0x1
    "00000111", --  667 - 0x29b  :    7 - 0x7
    "00000111", --  668 - 0x29c  :    7 - 0x7
    "00011111", --  669 - 0x29d  :   31 - 0x1f
    "00001111", --  670 - 0x29e  :   15 - 0xf
    "00000110", --  671 - 0x29f  :    6 - 0x6
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x2a
    "11000000", --  673 - 0x2a1  :  192 - 0xc0
    "11111000", --  674 - 0x2a2  :  248 - 0xf8
    "10000000", --  675 - 0x2a3  :  128 - 0x80
    "00100000", --  676 - 0x2a4  :   32 - 0x20
    "10010000", --  677 - 0x2a5  :  144 - 0x90
    "00111100", --  678 - 0x2a6  :   60 - 0x3c
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- plane 1
    "11000000", --  681 - 0x2a9  :  192 - 0xc0
    "11111000", --  682 - 0x2aa  :  248 - 0xf8
    "01100000", --  683 - 0x2ab  :   96 - 0x60
    "11011100", --  684 - 0x2ac  :  220 - 0xdc
    "01101110", --  685 - 0x2ad  :  110 - 0x6e
    "11000000", --  686 - 0x2ae  :  192 - 0xc0
    "11111011", --  687 - 0x2af  :  251 - 0xfb
    "11100100", --  688 - 0x2b0  :  228 - 0xe4 -- Sprite 0x2b
    "11111110", --  689 - 0x2b1  :  254 - 0xfe
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "11110001", --  691 - 0x2b3  :  241 - 0xf1
    "11111111", --  692 - 0x2b4  :  255 - 0xff
    "11111111", --  693 - 0x2b5  :  255 - 0xff
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "10000011", --  696 - 0x2b8  :  131 - 0x83 -- plane 1
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "11110000", --  698 - 0x2ba  :  240 - 0xf0
    "11110000", --  699 - 0x2bb  :  240 - 0xf0
    "11111100", --  700 - 0x2bc  :  252 - 0xfc
    "11111100", --  701 - 0x2bd  :  252 - 0xfc
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000111", --  704 - 0x2c0  :    7 - 0x7 -- Sprite 0x2c
    "00001111", --  705 - 0x2c1  :   15 - 0xf
    "00001111", --  706 - 0x2c2  :   15 - 0xf
    "00010010", --  707 - 0x2c3  :   18 - 0x12
    "00010011", --  708 - 0x2c4  :   19 - 0x13
    "00111000", --  709 - 0x2c5  :   56 - 0x38
    "01110000", --  710 - 0x2c6  :  112 - 0x70
    "11111111", --  711 - 0x2c7  :  255 - 0xff
    "00000111", --  712 - 0x2c8  :    7 - 0x7 -- plane 1
    "00001111", --  713 - 0x2c9  :   15 - 0xf
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00001101", --  715 - 0x2cb  :   13 - 0xd
    "00001100", --  716 - 0x2cc  :   12 - 0xc
    "00000111", --  717 - 0x2cd  :    7 - 0x7
    "00001111", --  718 - 0x2ce  :   15 - 0xf
    "00000010", --  719 - 0x2cf  :    2 - 0x2
    "11011111", --  720 - 0x2d0  :  223 - 0xdf -- Sprite 0x2d
    "00011110", --  721 - 0x2d1  :   30 - 0x1e
    "00011111", --  722 - 0x2d2  :   31 - 0x1f
    "00011111", --  723 - 0x2d3  :   31 - 0x1f
    "00011111", --  724 - 0x2d4  :   31 - 0x1f
    "00001111", --  725 - 0x2d5  :   15 - 0xf
    "00000111", --  726 - 0x2d6  :    7 - 0x7
    "00000001", --  727 - 0x2d7  :    1 - 0x1
    "00000001", --  728 - 0x2d8  :    1 - 0x1 -- plane 1
    "11110011", --  729 - 0x2d9  :  243 - 0xf3
    "01011111", --  730 - 0x2da  :   95 - 0x5f
    "00011111", --  731 - 0x2db  :   31 - 0x1f
    "00011111", --  732 - 0x2dc  :   31 - 0x1f
    "01001111", --  733 - 0x2dd  :   79 - 0x4f
    "00110111", --  734 - 0x2de  :   55 - 0x37
    "11000000", --  735 - 0x2df  :  192 - 0xc0
    "10000000", --  736 - 0x2e0  :  128 - 0x80 -- Sprite 0x2e
    "11110000", --  737 - 0x2e1  :  240 - 0xf0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "01000000", --  739 - 0x2e3  :   64 - 0x40
    "00100000", --  740 - 0x2e4  :   32 - 0x20
    "01111000", --  741 - 0x2e5  :  120 - 0x78
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "10000000", --  744 - 0x2e8  :  128 - 0x80 -- plane 1
    "11110000", --  745 - 0x2e9  :  240 - 0xf0
    "11000000", --  746 - 0x2ea  :  192 - 0xc0
    "10111000", --  747 - 0x2eb  :  184 - 0xb8
    "11011100", --  748 - 0x2ec  :  220 - 0xdc
    "10000000", --  749 - 0x2ed  :  128 - 0x80
    "11110000", --  750 - 0x2ee  :  240 - 0xf0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "11110000", --  752 - 0x2f0  :  240 - 0xf0 -- Sprite 0x2f
    "11100000", --  753 - 0x2f1  :  224 - 0xe0
    "11100000", --  754 - 0x2f2  :  224 - 0xe0
    "11110000", --  755 - 0x2f3  :  240 - 0xf0
    "11111010", --  756 - 0x2f4  :  250 - 0xfa
    "11111110", --  757 - 0x2f5  :  254 - 0xfe
    "11111100", --  758 - 0x2f6  :  252 - 0xfc
    "11011000", --  759 - 0x2f7  :  216 - 0xd8
    "10001111", --  760 - 0x2f8  :  143 - 0x8f -- plane 1
    "11100111", --  761 - 0x2f9  :  231 - 0xe7
    "11100000", --  762 - 0x2fa  :  224 - 0xe0
    "11110000", --  763 - 0x2fb  :  240 - 0xf0
    "11001000", --  764 - 0x2fc  :  200 - 0xc8
    "10001000", --  765 - 0x2fd  :  136 - 0x88
    "00010000", --  766 - 0x2fe  :   16 - 0x10
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000111", --  770 - 0x302  :    7 - 0x7
    "00001000", --  771 - 0x303  :    8 - 0x8
    "00010000", --  772 - 0x304  :   16 - 0x10
    "00100000", --  773 - 0x305  :   32 - 0x20
    "01000000", --  774 - 0x306  :   64 - 0x40
    "01000000", --  775 - 0x307  :   64 - 0x40
    "00000000", --  776 - 0x308  :    0 - 0x0 -- plane 1
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000111", --  779 - 0x30b  :    7 - 0x7
    "00001000", --  780 - 0x30c  :    8 - 0x8
    "00010000", --  781 - 0x30d  :   16 - 0x10
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "00100000", --  783 - 0x30f  :   32 - 0x20
    "01000000", --  784 - 0x310  :   64 - 0x40 -- Sprite 0x31
    "01000000", --  785 - 0x311  :   64 - 0x40
    "00100000", --  786 - 0x312  :   32 - 0x20
    "00010000", --  787 - 0x313  :   16 - 0x10
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00000111", --  789 - 0x315  :    7 - 0x7
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00100000", --  792 - 0x318  :   32 - 0x20 -- plane 1
    "00100000", --  793 - 0x319  :   32 - 0x20
    "00010000", --  794 - 0x31a  :   16 - 0x10
    "00001000", --  795 - 0x31b  :    8 - 0x8
    "00000111", --  796 - 0x31c  :    7 - 0x7
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  801 - 0x321  :    0 - 0x0
    "11100000", --  802 - 0x322  :  224 - 0xe0
    "00010000", --  803 - 0x323  :   16 - 0x10
    "00001000", --  804 - 0x324  :    8 - 0x8
    "00000100", --  805 - 0x325  :    4 - 0x4
    "00000010", --  806 - 0x326  :    2 - 0x2
    "00000010", --  807 - 0x327  :    2 - 0x2
    "00000000", --  808 - 0x328  :    0 - 0x0 -- plane 1
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "11100000", --  811 - 0x32b  :  224 - 0xe0
    "00010000", --  812 - 0x32c  :   16 - 0x10
    "00001000", --  813 - 0x32d  :    8 - 0x8
    "00000100", --  814 - 0x32e  :    4 - 0x4
    "00000100", --  815 - 0x32f  :    4 - 0x4
    "00000010", --  816 - 0x330  :    2 - 0x2 -- Sprite 0x33
    "00000010", --  817 - 0x331  :    2 - 0x2
    "00000100", --  818 - 0x332  :    4 - 0x4
    "00001000", --  819 - 0x333  :    8 - 0x8
    "00010000", --  820 - 0x334  :   16 - 0x10
    "11100000", --  821 - 0x335  :  224 - 0xe0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000100", --  824 - 0x338  :    4 - 0x4 -- plane 1
    "00000100", --  825 - 0x339  :    4 - 0x4
    "00001000", --  826 - 0x33a  :    8 - 0x8
    "00010000", --  827 - 0x33b  :   16 - 0x10
    "11100000", --  828 - 0x33c  :  224 - 0xe0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000011", --  836 - 0x344  :    3 - 0x3
    "00000100", --  837 - 0x345  :    4 - 0x4
    "00001000", --  838 - 0x346  :    8 - 0x8
    "00010000", --  839 - 0x347  :   16 - 0x10
    "00000000", --  840 - 0x348  :    0 - 0x0 -- plane 1
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000011", --  845 - 0x34d  :    3 - 0x3
    "00000100", --  846 - 0x34e  :    4 - 0x4
    "00001000", --  847 - 0x34f  :    8 - 0x8
    "00010000", --  848 - 0x350  :   16 - 0x10 -- Sprite 0x35
    "00001000", --  849 - 0x351  :    8 - 0x8
    "00000100", --  850 - 0x352  :    4 - 0x4
    "00000011", --  851 - 0x353  :    3 - 0x3
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00001000", --  856 - 0x358  :    8 - 0x8 -- plane 1
    "00000100", --  857 - 0x359  :    4 - 0x4
    "00000011", --  858 - 0x35a  :    3 - 0x3
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "11000000", --  868 - 0x364  :  192 - 0xc0
    "00100000", --  869 - 0x365  :   32 - 0x20
    "00010000", --  870 - 0x366  :   16 - 0x10
    "00001000", --  871 - 0x367  :    8 - 0x8
    "00000000", --  872 - 0x368  :    0 - 0x0 -- plane 1
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "11000000", --  877 - 0x36d  :  192 - 0xc0
    "00100000", --  878 - 0x36e  :   32 - 0x20
    "00010000", --  879 - 0x36f  :   16 - 0x10
    "00001000", --  880 - 0x370  :    8 - 0x8 -- Sprite 0x37
    "00010000", --  881 - 0x371  :   16 - 0x10
    "00100000", --  882 - 0x372  :   32 - 0x20
    "11000000", --  883 - 0x373  :  192 - 0xc0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00010000", --  888 - 0x378  :   16 - 0x10 -- plane 1
    "00100000", --  889 - 0x379  :   32 - 0x20
    "11000000", --  890 - 0x37a  :  192 - 0xc0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000001", --  903 - 0x387  :    1 - 0x1
    "00000000", --  904 - 0x388  :    0 - 0x0 -- plane 1
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000010", --  912 - 0x390  :    2 - 0x2 -- Sprite 0x39
    "00000001", --  913 - 0x391  :    1 - 0x1
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000001", --  920 - 0x398  :    1 - 0x1 -- plane 1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "10000000", --  944 - 0x3b0  :  128 - 0x80 -- Sprite 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- plane 1
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000001", --  963 - 0x3c3  :    1 - 0x1
    "00100001", --  964 - 0x3c4  :   33 - 0x21
    "00010000", --  965 - 0x3c5  :   16 - 0x10
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000001", --  969 - 0x3c9  :    1 - 0x1
    "00000001", --  970 - 0x3ca  :    1 - 0x1
    "01000000", --  971 - 0x3cb  :   64 - 0x40
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "01100000", --  976 - 0x3d0  :   96 - 0x60 -- Sprite 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00010000", --  979 - 0x3d3  :   16 - 0x10
    "00100001", --  980 - 0x3d4  :   33 - 0x21
    "00000001", --  981 - 0x3d5  :    1 - 0x1
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "10000000", --  984 - 0x3d8  :  128 - 0x80 -- plane 1
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "01000000", --  989 - 0x3dd  :   64 - 0x40
    "00000001", --  990 - 0x3de  :    1 - 0x1
    "00000001", --  991 - 0x3df  :    1 - 0x1
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00001000", --  996 - 0x3e4  :    8 - 0x8
    "00010000", --  997 - 0x3e5  :   16 - 0x10
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000100", -- 1003 - 0x3eb  :    4 - 0x4
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00001100", -- 1008 - 0x3f0  :   12 - 0xc -- Sprite 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00010000", -- 1011 - 0x3f3  :   16 - 0x10
    "00001000", -- 1012 - 0x3f4  :    8 - 0x8
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000010", -- 1016 - 0x3f8  :    2 - 0x2 -- plane 1
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000100", -- 1021 - 0x3fd  :    4 - 0x4
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000100", -- 1024 - 0x400  :    4 - 0x4 -- Sprite 0x40
    "00000010", -- 1025 - 0x401  :    2 - 0x2
    "00000001", -- 1026 - 0x402  :    1 - 0x1
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00001111", -- 1032 - 0x408  :   15 - 0xf -- plane 1
    "00000111", -- 1033 - 0x409  :    7 - 0x7
    "00000011", -- 1034 - 0x40a  :    3 - 0x3
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000001", -- 1037 - 0x40d  :    1 - 0x1
    "00000001", -- 1038 - 0x40e  :    1 - 0x1
    "00000001", -- 1039 - 0x40f  :    1 - 0x1
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x41
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000001", -- 1046 - 0x416  :    1 - 0x1
    "00000011", -- 1047 - 0x417  :    3 - 0x3
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- plane 1
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000001", -- 1054 - 0x41e  :    1 - 0x1
    "00000011", -- 1055 - 0x41f  :    3 - 0x3
    "00000111", -- 1056 - 0x420  :    7 - 0x7 -- Sprite 0x42
    "00000111", -- 1057 - 0x421  :    7 - 0x7
    "00000111", -- 1058 - 0x422  :    7 - 0x7
    "00000011", -- 1059 - 0x423  :    3 - 0x3
    "00000001", -- 1060 - 0x424  :    1 - 0x1
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000111", -- 1064 - 0x428  :    7 - 0x7 -- plane 1
    "00000111", -- 1065 - 0x429  :    7 - 0x7
    "00000111", -- 1066 - 0x42a  :    7 - 0x7
    "00000111", -- 1067 - 0x42b  :    7 - 0x7
    "00000011", -- 1068 - 0x42c  :    3 - 0x3
    "00000001", -- 1069 - 0x42d  :    1 - 0x1
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x43
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- plane 1
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x44
    "01000010", -- 1089 - 0x441  :   66 - 0x42
    "00111001", -- 1090 - 0x442  :   57 - 0x39
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- plane 1
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11111111", -- 1100 - 0x44c  :  255 - 0xff
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "01111111", -- 1104 - 0x450  :  127 - 0x7f -- Sprite 0x45
    "00111111", -- 1105 - 0x451  :   63 - 0x3f
    "00011111", -- 1106 - 0x452  :   31 - 0x1f
    "00001111", -- 1107 - 0x453  :   15 - 0xf
    "00011111", -- 1108 - 0x454  :   31 - 0x1f
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- plane 1
    "01111111", -- 1113 - 0x459  :  127 - 0x7f
    "00111111", -- 1114 - 0x45a  :   63 - 0x3f
    "00011111", -- 1115 - 0x45b  :   31 - 0x1f
    "00011111", -- 1116 - 0x45c  :   31 - 0x1f
    "11111111", -- 1117 - 0x45d  :  255 - 0xff
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11111111", -- 1119 - 0x45f  :  255 - 0xff
    "11111000", -- 1120 - 0x460  :  248 - 0xf8 -- Sprite 0x46
    "11110111", -- 1121 - 0x461  :  247 - 0xf7
    "11101111", -- 1122 - 0x462  :  239 - 0xef
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "11111110", -- 1125 - 0x465  :  254 - 0xfe
    "01111110", -- 1126 - 0x466  :  126 - 0x7e
    "00111110", -- 1127 - 0x467  :   62 - 0x3e
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- plane 1
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "11111111", -- 1130 - 0x46a  :  255 - 0xff
    "11111111", -- 1131 - 0x46b  :  255 - 0xff
    "11111111", -- 1132 - 0x46c  :  255 - 0xff
    "11111111", -- 1133 - 0x46d  :  255 - 0xff
    "11111111", -- 1134 - 0x46e  :  255 - 0xff
    "01111111", -- 1135 - 0x46f  :  127 - 0x7f
    "00000111", -- 1136 - 0x470  :    7 - 0x7 -- Sprite 0x47
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000111", -- 1144 - 0x478  :    7 - 0x7 -- plane 1
    "00000011", -- 1145 - 0x479  :    3 - 0x3
    "00000011", -- 1146 - 0x47a  :    3 - 0x3
    "00000001", -- 1147 - 0x47b  :    1 - 0x1
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x48
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "11000000", -- 1155 - 0x483  :  192 - 0xc0
    "11100000", -- 1156 - 0x484  :  224 - 0xe0
    "11110000", -- 1157 - 0x485  :  240 - 0xf0
    "11011011", -- 1158 - 0x486  :  219 - 0xdb
    "11110110", -- 1159 - 0x487  :  246 - 0xf6
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- plane 1
    "10000000", -- 1161 - 0x489  :  128 - 0x80
    "10000000", -- 1162 - 0x48a  :  128 - 0x80
    "11000000", -- 1163 - 0x48b  :  192 - 0xc0
    "11100000", -- 1164 - 0x48c  :  224 - 0xe0
    "11110000", -- 1165 - 0x48d  :  240 - 0xf0
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11001011", -- 1168 - 0x490  :  203 - 0xcb -- Sprite 0x49
    "11100000", -- 1169 - 0x491  :  224 - 0xe0
    "11000100", -- 1170 - 0x492  :  196 - 0xc4
    "00000010", -- 1171 - 0x493  :    2 - 0x2
    "11010001", -- 1172 - 0x494  :  209 - 0xd1
    "11100001", -- 1173 - 0x495  :  225 - 0xe1
    "11010001", -- 1174 - 0x496  :  209 - 0xd1
    "10000011", -- 1175 - 0x497  :  131 - 0x83
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- plane 1
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11111111", -- 1179 - 0x49b  :  255 - 0xff
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "00001111", -- 1184 - 0x4a0  :   15 - 0xf -- Sprite 0x4a
    "11111111", -- 1185 - 0x4a1  :  255 - 0xff
    "11100000", -- 1186 - 0x4a2  :  224 - 0xe0
    "10001111", -- 1187 - 0x4a3  :  143 - 0x8f
    "01101110", -- 1188 - 0x4a4  :  110 - 0x6e
    "01000100", -- 1189 - 0x4a5  :   68 - 0x44
    "11101110", -- 1190 - 0x4a6  :  238 - 0xee
    "01100000", -- 1191 - 0x4a7  :   96 - 0x60
    "11111111", -- 1192 - 0x4a8  :  255 - 0xff -- plane 1
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "11111111", -- 1194 - 0x4aa  :  255 - 0xff
    "11110000", -- 1195 - 0x4ab  :  240 - 0xf0
    "10000000", -- 1196 - 0x4ac  :  128 - 0x80
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "10011111", -- 1199 - 0x4af  :  159 - 0x9f
    "10000011", -- 1200 - 0x4b0  :  131 - 0x83 -- Sprite 0x4b
    "11100000", -- 1201 - 0x4b1  :  224 - 0xe0
    "11100100", -- 1202 - 0x4b2  :  228 - 0xe4
    "11000110", -- 1203 - 0x4b3  :  198 - 0xc6
    "01100001", -- 1204 - 0x4b4  :   97 - 0x61
    "00110011", -- 1205 - 0x4b5  :   51 - 0x33
    "00011111", -- 1206 - 0x4b6  :   31 - 0x1f
    "00001111", -- 1207 - 0x4b7  :   15 - 0xf
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- plane 1
    "11111111", -- 1209 - 0x4b9  :  255 - 0xff
    "11111001", -- 1210 - 0x4ba  :  249 - 0xf9
    "11111001", -- 1211 - 0x4bb  :  249 - 0xf9
    "01111111", -- 1212 - 0x4bc  :  127 - 0x7f
    "00111111", -- 1213 - 0x4bd  :   63 - 0x3f
    "00011111", -- 1214 - 0x4be  :   31 - 0x1f
    "00001111", -- 1215 - 0x4bf  :   15 - 0xf
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x4c
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000011", -- 1219 - 0x4c3  :    3 - 0x3
    "00000111", -- 1220 - 0x4c4  :    7 - 0x7
    "00001111", -- 1221 - 0x4c5  :   15 - 0xf
    "01011011", -- 1222 - 0x4c6  :   91 - 0x5b
    "10100111", -- 1223 - 0x4c7  :  167 - 0xa7
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- plane 1
    "00000001", -- 1225 - 0x4c9  :    1 - 0x1
    "00000001", -- 1226 - 0x4ca  :    1 - 0x1
    "00000011", -- 1227 - 0x4cb  :    3 - 0x3
    "00000111", -- 1228 - 0x4cc  :    7 - 0x7
    "00001111", -- 1229 - 0x4cd  :   15 - 0xf
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "01110011", -- 1232 - 0x4d0  :  115 - 0x73 -- Sprite 0x4d
    "00000111", -- 1233 - 0x4d1  :    7 - 0x7
    "00100111", -- 1234 - 0x4d2  :   39 - 0x27
    "01000000", -- 1235 - 0x4d3  :   64 - 0x40
    "10001011", -- 1236 - 0x4d4  :  139 - 0x8b
    "10000111", -- 1237 - 0x4d5  :  135 - 0x87
    "10001011", -- 1238 - 0x4d6  :  139 - 0x8b
    "11000001", -- 1239 - 0x4d7  :  193 - 0xc1
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- plane 1
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11111111", -- 1244 - 0x4dc  :  255 - 0xff
    "11111111", -- 1245 - 0x4dd  :  255 - 0xff
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11110000", -- 1248 - 0x4e0  :  240 - 0xf0 -- Sprite 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "00001111", -- 1250 - 0x4e2  :   15 - 0xf
    "11100001", -- 1251 - 0x4e3  :  225 - 0xe1
    "11101100", -- 1252 - 0x4e4  :  236 - 0xec
    "01000100", -- 1253 - 0x4e5  :   68 - 0x44
    "11101110", -- 1254 - 0x4e6  :  238 - 0xee
    "00001100", -- 1255 - 0x4e7  :   12 - 0xc
    "11111111", -- 1256 - 0x4e8  :  255 - 0xff -- plane 1
    "11111111", -- 1257 - 0x4e9  :  255 - 0xff
    "11111111", -- 1258 - 0x4ea  :  255 - 0xff
    "00011111", -- 1259 - 0x4eb  :   31 - 0x1f
    "00000011", -- 1260 - 0x4ec  :    3 - 0x3
    "00000001", -- 1261 - 0x4ed  :    1 - 0x1
    "00000001", -- 1262 - 0x4ee  :    1 - 0x1
    "11110011", -- 1263 - 0x4ef  :  243 - 0xf3
    "10000000", -- 1264 - 0x4f0  :  128 - 0x80 -- Sprite 0x4f
    "00001110", -- 1265 - 0x4f1  :   14 - 0xe
    "01001110", -- 1266 - 0x4f2  :   78 - 0x4e
    "11000110", -- 1267 - 0x4f3  :  198 - 0xc6
    "00001100", -- 1268 - 0x4f4  :   12 - 0xc
    "10011000", -- 1269 - 0x4f5  :  152 - 0x98
    "11110000", -- 1270 - 0x4f6  :  240 - 0xf0
    "11100000", -- 1271 - 0x4f7  :  224 - 0xe0
    "11111111", -- 1272 - 0x4f8  :  255 - 0xff -- plane 1
    "11111111", -- 1273 - 0x4f9  :  255 - 0xff
    "00111111", -- 1274 - 0x4fa  :   63 - 0x3f
    "00111111", -- 1275 - 0x4fb  :   63 - 0x3f
    "11111100", -- 1276 - 0x4fc  :  252 - 0xfc
    "11111000", -- 1277 - 0x4fd  :  248 - 0xf8
    "11110000", -- 1278 - 0x4fe  :  240 - 0xf0
    "11100000", -- 1279 - 0x4ff  :  224 - 0xe0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0x50
    "01000010", -- 1281 - 0x501  :   66 - 0x42
    "10011100", -- 1282 - 0x502  :  156 - 0x9c
    "11111111", -- 1283 - 0x503  :  255 - 0xff
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "11111111", -- 1288 - 0x508  :  255 - 0xff -- plane 1
    "11111111", -- 1289 - 0x509  :  255 - 0xff
    "11111111", -- 1290 - 0x50a  :  255 - 0xff
    "11111111", -- 1291 - 0x50b  :  255 - 0xff
    "11111111", -- 1292 - 0x50c  :  255 - 0xff
    "11111111", -- 1293 - 0x50d  :  255 - 0xff
    "11111111", -- 1294 - 0x50e  :  255 - 0xff
    "11111111", -- 1295 - 0x50f  :  255 - 0xff
    "11111110", -- 1296 - 0x510  :  254 - 0xfe -- Sprite 0x51
    "11111100", -- 1297 - 0x511  :  252 - 0xfc
    "11111000", -- 1298 - 0x512  :  248 - 0xf8
    "11110000", -- 1299 - 0x513  :  240 - 0xf0
    "11111000", -- 1300 - 0x514  :  248 - 0xf8
    "11111111", -- 1301 - 0x515  :  255 - 0xff
    "11111111", -- 1302 - 0x516  :  255 - 0xff
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "11111111", -- 1304 - 0x518  :  255 - 0xff -- plane 1
    "11111110", -- 1305 - 0x519  :  254 - 0xfe
    "11111100", -- 1306 - 0x51a  :  252 - 0xfc
    "11111000", -- 1307 - 0x51b  :  248 - 0xf8
    "11111000", -- 1308 - 0x51c  :  248 - 0xf8
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "00011111", -- 1312 - 0x520  :   31 - 0x1f -- Sprite 0x52
    "11101111", -- 1313 - 0x521  :  239 - 0xef
    "11110111", -- 1314 - 0x522  :  247 - 0xf7
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111110", -- 1317 - 0x525  :  254 - 0xfe
    "01111100", -- 1318 - 0x526  :  124 - 0x7c
    "01110000", -- 1319 - 0x527  :  112 - 0x70
    "11111111", -- 1320 - 0x528  :  255 - 0xff -- plane 1
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11111111", -- 1325 - 0x52d  :  255 - 0xff
    "11111110", -- 1326 - 0x52e  :  254 - 0xfe
    "11111100", -- 1327 - 0x52f  :  252 - 0xfc
    "11100000", -- 1328 - 0x530  :  224 - 0xe0 -- Sprite 0x53
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "11100000", -- 1336 - 0x538  :  224 - 0xe0 -- plane 1
    "10000000", -- 1337 - 0x539  :  128 - 0x80
    "10000000", -- 1338 - 0x53a  :  128 - 0x80
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00100000", -- 1344 - 0x540  :   32 - 0x20 -- Sprite 0x54
    "01000000", -- 1345 - 0x541  :   64 - 0x40
    "10000000", -- 1346 - 0x542  :  128 - 0x80
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "11110000", -- 1352 - 0x548  :  240 - 0xf0 -- plane 1
    "11100000", -- 1353 - 0x549  :  224 - 0xe0
    "11000000", -- 1354 - 0x54a  :  192 - 0xc0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "10000000", -- 1357 - 0x54d  :  128 - 0x80
    "10000000", -- 1358 - 0x54e  :  128 - 0x80
    "10000000", -- 1359 - 0x54f  :  128 - 0x80
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0x55
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "10000000", -- 1366 - 0x556  :  128 - 0x80
    "11000000", -- 1367 - 0x557  :  192 - 0xc0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- plane 1
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "10000000", -- 1374 - 0x55e  :  128 - 0x80
    "11000000", -- 1375 - 0x55f  :  192 - 0xc0
    "11100000", -- 1376 - 0x560  :  224 - 0xe0 -- Sprite 0x56
    "11100000", -- 1377 - 0x561  :  224 - 0xe0
    "11100000", -- 1378 - 0x562  :  224 - 0xe0
    "11000000", -- 1379 - 0x563  :  192 - 0xc0
    "10000000", -- 1380 - 0x564  :  128 - 0x80
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "11100000", -- 1384 - 0x568  :  224 - 0xe0 -- plane 1
    "11100000", -- 1385 - 0x569  :  224 - 0xe0
    "11100000", -- 1386 - 0x56a  :  224 - 0xe0
    "11100000", -- 1387 - 0x56b  :  224 - 0xe0
    "11000000", -- 1388 - 0x56c  :  192 - 0xc0
    "10000000", -- 1389 - 0x56d  :  128 - 0x80
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0x57
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- plane 1
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Sprite 0x58
    "11111111", -- 1409 - 0x581  :  255 - 0xff
    "11111111", -- 1410 - 0x582  :  255 - 0xff
    "11111111", -- 1411 - 0x583  :  255 - 0xff
    "11111111", -- 1412 - 0x584  :  255 - 0xff
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "11111111", -- 1416 - 0x588  :  255 - 0xff -- plane 1
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11111111", -- 1418 - 0x58a  :  255 - 0xff
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11111111", -- 1421 - 0x58d  :  255 - 0xff
    "11111111", -- 1422 - 0x58e  :  255 - 0xff
    "11111111", -- 1423 - 0x58f  :  255 - 0xff
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Sprite 0x59
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "11111111", -- 1426 - 0x592  :  255 - 0xff
    "11111111", -- 1427 - 0x593  :  255 - 0xff
    "11111111", -- 1428 - 0x594  :  255 - 0xff
    "11111111", -- 1429 - 0x595  :  255 - 0xff
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff -- plane 1
    "11111111", -- 1433 - 0x599  :  255 - 0xff
    "11111111", -- 1434 - 0x59a  :  255 - 0xff
    "11111111", -- 1435 - 0x59b  :  255 - 0xff
    "11111111", -- 1436 - 0x59c  :  255 - 0xff
    "11111111", -- 1437 - 0x59d  :  255 - 0xff
    "11111111", -- 1438 - 0x59e  :  255 - 0xff
    "11111111", -- 1439 - 0x59f  :  255 - 0xff
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Sprite 0x5a
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "11111111", -- 1442 - 0x5a2  :  255 - 0xff
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "11111111", -- 1445 - 0x5a5  :  255 - 0xff
    "11111111", -- 1446 - 0x5a6  :  255 - 0xff
    "11111111", -- 1447 - 0x5a7  :  255 - 0xff
    "11111111", -- 1448 - 0x5a8  :  255 - 0xff -- plane 1
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111111", -- 1450 - 0x5aa  :  255 - 0xff
    "11111111", -- 1451 - 0x5ab  :  255 - 0xff
    "11111111", -- 1452 - 0x5ac  :  255 - 0xff
    "11111111", -- 1453 - 0x5ad  :  255 - 0xff
    "11111111", -- 1454 - 0x5ae  :  255 - 0xff
    "11111111", -- 1455 - 0x5af  :  255 - 0xff
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0x5b
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11111111", -- 1461 - 0x5b5  :  255 - 0xff
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- plane 1
    "11111111", -- 1465 - 0x5b9  :  255 - 0xff
    "11111111", -- 1466 - 0x5ba  :  255 - 0xff
    "11111111", -- 1467 - 0x5bb  :  255 - 0xff
    "11111111", -- 1468 - 0x5bc  :  255 - 0xff
    "11111111", -- 1469 - 0x5bd  :  255 - 0xff
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0x5c
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "11111111", -- 1478 - 0x5c6  :  255 - 0xff
    "11111111", -- 1479 - 0x5c7  :  255 - 0xff
    "11111111", -- 1480 - 0x5c8  :  255 - 0xff -- plane 1
    "11111111", -- 1481 - 0x5c9  :  255 - 0xff
    "11111111", -- 1482 - 0x5ca  :  255 - 0xff
    "11111111", -- 1483 - 0x5cb  :  255 - 0xff
    "11111111", -- 1484 - 0x5cc  :  255 - 0xff
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "11111111", -- 1486 - 0x5ce  :  255 - 0xff
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0x5d
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "11111111", -- 1490 - 0x5d2  :  255 - 0xff
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "11111111", -- 1492 - 0x5d4  :  255 - 0xff
    "11111111", -- 1493 - 0x5d5  :  255 - 0xff
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "11111111", -- 1496 - 0x5d8  :  255 - 0xff -- plane 1
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111111", -- 1499 - 0x5db  :  255 - 0xff
    "11111111", -- 1500 - 0x5dc  :  255 - 0xff
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0x5e
    "11111111", -- 1505 - 0x5e1  :  255 - 0xff
    "11111111", -- 1506 - 0x5e2  :  255 - 0xff
    "11111111", -- 1507 - 0x5e3  :  255 - 0xff
    "11111111", -- 1508 - 0x5e4  :  255 - 0xff
    "11111111", -- 1509 - 0x5e5  :  255 - 0xff
    "11111111", -- 1510 - 0x5e6  :  255 - 0xff
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "11111111", -- 1512 - 0x5e8  :  255 - 0xff -- plane 1
    "11111111", -- 1513 - 0x5e9  :  255 - 0xff
    "11111111", -- 1514 - 0x5ea  :  255 - 0xff
    "11111111", -- 1515 - 0x5eb  :  255 - 0xff
    "11111111", -- 1516 - 0x5ec  :  255 - 0xff
    "11111111", -- 1517 - 0x5ed  :  255 - 0xff
    "11111111", -- 1518 - 0x5ee  :  255 - 0xff
    "11111111", -- 1519 - 0x5ef  :  255 - 0xff
    "11111111", -- 1520 - 0x5f0  :  255 - 0xff -- Sprite 0x5f
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "11111111", -- 1522 - 0x5f2  :  255 - 0xff
    "11111111", -- 1523 - 0x5f3  :  255 - 0xff
    "11111111", -- 1524 - 0x5f4  :  255 - 0xff
    "11111111", -- 1525 - 0x5f5  :  255 - 0xff
    "11111111", -- 1526 - 0x5f6  :  255 - 0xff
    "11111111", -- 1527 - 0x5f7  :  255 - 0xff
    "11111111", -- 1528 - 0x5f8  :  255 - 0xff -- plane 1
    "11111111", -- 1529 - 0x5f9  :  255 - 0xff
    "11111111", -- 1530 - 0x5fa  :  255 - 0xff
    "11111111", -- 1531 - 0x5fb  :  255 - 0xff
    "11111111", -- 1532 - 0x5fc  :  255 - 0xff
    "11111111", -- 1533 - 0x5fd  :  255 - 0xff
    "11111111", -- 1534 - 0x5fe  :  255 - 0xff
    "11111111", -- 1535 - 0x5ff  :  255 - 0xff
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00011111", -- 1538 - 0x602  :   31 - 0x1f
    "00111111", -- 1539 - 0x603  :   63 - 0x3f
    "00111111", -- 1540 - 0x604  :   63 - 0x3f
    "01111111", -- 1541 - 0x605  :  127 - 0x7f
    "01111111", -- 1542 - 0x606  :  127 - 0x7f
    "01111111", -- 1543 - 0x607  :  127 - 0x7f
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- plane 1
    "00001111", -- 1545 - 0x609  :   15 - 0xf
    "00101000", -- 1546 - 0x60a  :   40 - 0x28
    "01011100", -- 1547 - 0x60b  :   92 - 0x5c
    "00111111", -- 1548 - 0x60c  :   63 - 0x3f
    "01111111", -- 1549 - 0x60d  :  127 - 0x7f
    "01111111", -- 1550 - 0x60e  :  127 - 0x7f
    "01111111", -- 1551 - 0x60f  :  127 - 0x7f
    "01111111", -- 1552 - 0x610  :  127 - 0x7f -- Sprite 0x61
    "00111110", -- 1553 - 0x611  :   62 - 0x3e
    "00011111", -- 1554 - 0x612  :   31 - 0x1f
    "00011111", -- 1555 - 0x613  :   31 - 0x1f
    "00001111", -- 1556 - 0x614  :   15 - 0xf
    "00001111", -- 1557 - 0x615  :   15 - 0xf
    "00001111", -- 1558 - 0x616  :   15 - 0xf
    "00000111", -- 1559 - 0x617  :    7 - 0x7
    "01111111", -- 1560 - 0x618  :  127 - 0x7f -- plane 1
    "00111110", -- 1561 - 0x619  :   62 - 0x3e
    "00011111", -- 1562 - 0x61a  :   31 - 0x1f
    "00011111", -- 1563 - 0x61b  :   31 - 0x1f
    "00001000", -- 1564 - 0x61c  :    8 - 0x8
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0x62
    "01100000", -- 1569 - 0x621  :   96 - 0x60
    "11110000", -- 1570 - 0x622  :  240 - 0xf0
    "11111000", -- 1571 - 0x623  :  248 - 0xf8
    "11111000", -- 1572 - 0x624  :  248 - 0xf8
    "11111000", -- 1573 - 0x625  :  248 - 0xf8
    "11111100", -- 1574 - 0x626  :  252 - 0xfc
    "11111100", -- 1575 - 0x627  :  252 - 0xfc
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- plane 1
    "10000000", -- 1577 - 0x629  :  128 - 0x80
    "01000000", -- 1578 - 0x62a  :   64 - 0x40
    "11000100", -- 1579 - 0x62b  :  196 - 0xc4
    "11110110", -- 1580 - 0x62c  :  246 - 0xf6
    "11111110", -- 1581 - 0x62d  :  254 - 0xfe
    "11111100", -- 1582 - 0x62e  :  252 - 0xfc
    "11111100", -- 1583 - 0x62f  :  252 - 0xfc
    "11111000", -- 1584 - 0x630  :  248 - 0xf8 -- Sprite 0x63
    "11110000", -- 1585 - 0x631  :  240 - 0xf0
    "11110000", -- 1586 - 0x632  :  240 - 0xf0
    "11100000", -- 1587 - 0x633  :  224 - 0xe0
    "10000000", -- 1588 - 0x634  :  128 - 0x80
    "10000000", -- 1589 - 0x635  :  128 - 0x80
    "11000000", -- 1590 - 0x636  :  192 - 0xc0
    "11000000", -- 1591 - 0x637  :  192 - 0xc0
    "11111000", -- 1592 - 0x638  :  248 - 0xf8 -- plane 1
    "11110000", -- 1593 - 0x639  :  240 - 0xf0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "10000000", -- 1596 - 0x63c  :  128 - 0x80
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00011111", -- 1601 - 0x641  :   31 - 0x1f
    "00111111", -- 1602 - 0x642  :   63 - 0x3f
    "01111111", -- 1603 - 0x643  :  127 - 0x7f
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "11111111", -- 1605 - 0x645  :  255 - 0xff
    "00111110", -- 1606 - 0x646  :   62 - 0x3e
    "00001111", -- 1607 - 0x647  :   15 - 0xf
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- plane 1
    "00011100", -- 1609 - 0x649  :   28 - 0x1c
    "00111111", -- 1610 - 0x64a  :   63 - 0x3f
    "01111111", -- 1611 - 0x64b  :  127 - 0x7f
    "11111111", -- 1612 - 0x64c  :  255 - 0xff
    "11111111", -- 1613 - 0x64d  :  255 - 0xff
    "00111110", -- 1614 - 0x64e  :   62 - 0x3e
    "01110000", -- 1615 - 0x64f  :  112 - 0x70
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000001", -- 1619 - 0x653  :    1 - 0x1
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- plane 1
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0x66
    "11100000", -- 1633 - 0x661  :  224 - 0xe0
    "11110000", -- 1634 - 0x662  :  240 - 0xf0
    "11111100", -- 1635 - 0x663  :  252 - 0xfc
    "11111110", -- 1636 - 0x664  :  254 - 0xfe
    "11111110", -- 1637 - 0x665  :  254 - 0xfe
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "11111100", -- 1639 - 0x667  :  252 - 0xfc
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- plane 1
    "01100000", -- 1641 - 0x669  :   96 - 0x60
    "11110000", -- 1642 - 0x66a  :  240 - 0xf0
    "11111000", -- 1643 - 0x66b  :  248 - 0xf8
    "11111100", -- 1644 - 0x66c  :  252 - 0xfc
    "11111100", -- 1645 - 0x66d  :  252 - 0xfc
    "11111100", -- 1646 - 0x66e  :  252 - 0xfc
    "11111111", -- 1647 - 0x66f  :  255 - 0xff
    "01111100", -- 1648 - 0x670  :  124 - 0x7c -- Sprite 0x67
    "11111100", -- 1649 - 0x671  :  252 - 0xfc
    "11111000", -- 1650 - 0x672  :  248 - 0xf8
    "11110000", -- 1651 - 0x673  :  240 - 0xf0
    "11100000", -- 1652 - 0x674  :  224 - 0xe0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "01111100", -- 1656 - 0x678  :  124 - 0x7c -- plane 1
    "11111100", -- 1657 - 0x679  :  252 - 0xfc
    "10001000", -- 1658 - 0x67a  :  136 - 0x88
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0x68
    "00000111", -- 1665 - 0x681  :    7 - 0x7
    "00000111", -- 1666 - 0x682  :    7 - 0x7
    "00001111", -- 1667 - 0x683  :   15 - 0xf
    "00001111", -- 1668 - 0x684  :   15 - 0xf
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00011111", -- 1670 - 0x686  :   31 - 0x1f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- plane 1
    "00000111", -- 1673 - 0x689  :    7 - 0x7
    "00000011", -- 1674 - 0x68a  :    3 - 0x3
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000111", -- 1677 - 0x68d  :    7 - 0x7
    "00000100", -- 1678 - 0x68e  :    4 - 0x4
    "00000100", -- 1679 - 0x68f  :    4 - 0x4
    "01111111", -- 1680 - 0x690  :  127 - 0x7f -- Sprite 0x69
    "01111111", -- 1681 - 0x691  :  127 - 0x7f
    "00011111", -- 1682 - 0x692  :   31 - 0x1f
    "00011111", -- 1683 - 0x693  :   31 - 0x1f
    "00011111", -- 1684 - 0x694  :   31 - 0x1f
    "00011110", -- 1685 - 0x695  :   30 - 0x1e
    "00001111", -- 1686 - 0x696  :   15 - 0xf
    "00011111", -- 1687 - 0x697  :   31 - 0x1f
    "00001100", -- 1688 - 0x698  :   12 - 0xc -- plane 1
    "10011110", -- 1689 - 0x699  :  158 - 0x9e
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "00011111", -- 1691 - 0x69b  :   31 - 0x1f
    "00011111", -- 1692 - 0x69c  :   31 - 0x1f
    "00011110", -- 1693 - 0x69d  :   30 - 0x1e
    "00001111", -- 1694 - 0x69e  :   15 - 0xf
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "11100000", -- 1697 - 0x6a1  :  224 - 0xe0
    "11100000", -- 1698 - 0x6a2  :  224 - 0xe0
    "11110000", -- 1699 - 0x6a3  :  240 - 0xf0
    "11110000", -- 1700 - 0x6a4  :  240 - 0xf0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "11111000", -- 1702 - 0x6a6  :  248 - 0xf8
    "11111100", -- 1703 - 0x6a7  :  252 - 0xfc
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- plane 1
    "11100000", -- 1705 - 0x6a9  :  224 - 0xe0
    "11000000", -- 1706 - 0x6aa  :  192 - 0xc0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "11100000", -- 1709 - 0x6ad  :  224 - 0xe0
    "00100000", -- 1710 - 0x6ae  :   32 - 0x20
    "00100000", -- 1711 - 0x6af  :   32 - 0x20
    "11111110", -- 1712 - 0x6b0  :  254 - 0xfe -- Sprite 0x6b
    "11111110", -- 1713 - 0x6b1  :  254 - 0xfe
    "11111000", -- 1714 - 0x6b2  :  248 - 0xf8
    "11111000", -- 1715 - 0x6b3  :  248 - 0xf8
    "11111000", -- 1716 - 0x6b4  :  248 - 0xf8
    "01111000", -- 1717 - 0x6b5  :  120 - 0x78
    "11110000", -- 1718 - 0x6b6  :  240 - 0xf0
    "11111000", -- 1719 - 0x6b7  :  248 - 0xf8
    "00110000", -- 1720 - 0x6b8  :   48 - 0x30 -- plane 1
    "01111001", -- 1721 - 0x6b9  :  121 - 0x79
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111000", -- 1723 - 0x6bb  :  248 - 0xf8
    "11111000", -- 1724 - 0x6bc  :  248 - 0xf8
    "01111000", -- 1725 - 0x6bd  :  120 - 0x78
    "11110000", -- 1726 - 0x6be  :  240 - 0xf0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000011", -- 1728 - 0x6c0  :    3 - 0x3 -- Sprite 0x6c
    "00000111", -- 1729 - 0x6c1  :    7 - 0x7
    "00000101", -- 1730 - 0x6c2  :    5 - 0x5
    "00001000", -- 1731 - 0x6c3  :    8 - 0x8
    "00011011", -- 1732 - 0x6c4  :   27 - 0x1b
    "00011001", -- 1733 - 0x6c5  :   25 - 0x19
    "00000101", -- 1734 - 0x6c6  :    5 - 0x5
    "00111111", -- 1735 - 0x6c7  :   63 - 0x3f
    "00000011", -- 1736 - 0x6c8  :    3 - 0x3 -- plane 1
    "00000111", -- 1737 - 0x6c9  :    7 - 0x7
    "00000010", -- 1738 - 0x6ca  :    2 - 0x2
    "00000111", -- 1739 - 0x6cb  :    7 - 0x7
    "00000100", -- 1740 - 0x6cc  :    4 - 0x4
    "01000110", -- 1741 - 0x6cd  :   70 - 0x46
    "11100011", -- 1742 - 0x6ce  :  227 - 0xe3
    "11000010", -- 1743 - 0x6cf  :  194 - 0xc2
    "00111111", -- 1744 - 0x6d0  :   63 - 0x3f -- Sprite 0x6d
    "00001111", -- 1745 - 0x6d1  :   15 - 0xf
    "00000101", -- 1746 - 0x6d2  :    5 - 0x5
    "00110111", -- 1747 - 0x6d3  :   55 - 0x37
    "00111111", -- 1748 - 0x6d4  :   63 - 0x3f
    "00111111", -- 1749 - 0x6d5  :   63 - 0x3f
    "00111110", -- 1750 - 0x6d6  :   62 - 0x3e
    "00011100", -- 1751 - 0x6d7  :   28 - 0x1c
    "01000010", -- 1752 - 0x6d8  :   66 - 0x42 -- plane 1
    "00000111", -- 1753 - 0x6d9  :    7 - 0x7
    "00000111", -- 1754 - 0x6da  :    7 - 0x7
    "00000111", -- 1755 - 0x6db  :    7 - 0x7
    "00000111", -- 1756 - 0x6dc  :    7 - 0x7
    "00000011", -- 1757 - 0x6dd  :    3 - 0x3
    "00000010", -- 1758 - 0x6de  :    2 - 0x2
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "11100000", -- 1760 - 0x6e0  :  224 - 0xe0 -- Sprite 0x6e
    "11110000", -- 1761 - 0x6e1  :  240 - 0xf0
    "01010000", -- 1762 - 0x6e2  :   80 - 0x50
    "00001000", -- 1763 - 0x6e3  :    8 - 0x8
    "01101100", -- 1764 - 0x6e4  :  108 - 0x6c
    "11001100", -- 1765 - 0x6e5  :  204 - 0xcc
    "11010000", -- 1766 - 0x6e6  :  208 - 0xd0
    "11111110", -- 1767 - 0x6e7  :  254 - 0xfe
    "11100000", -- 1768 - 0x6e8  :  224 - 0xe0 -- plane 1
    "11110000", -- 1769 - 0x6e9  :  240 - 0xf0
    "10100000", -- 1770 - 0x6ea  :  160 - 0xa0
    "11110000", -- 1771 - 0x6eb  :  240 - 0xf0
    "10010000", -- 1772 - 0x6ec  :  144 - 0x90
    "00110010", -- 1773 - 0x6ed  :   50 - 0x32
    "11100011", -- 1774 - 0x6ee  :  227 - 0xe3
    "00100001", -- 1775 - 0x6ef  :   33 - 0x21
    "11111110", -- 1776 - 0x6f0  :  254 - 0xfe -- Sprite 0x6f
    "11111000", -- 1777 - 0x6f1  :  248 - 0xf8
    "11010000", -- 1778 - 0x6f2  :  208 - 0xd0
    "11111011", -- 1779 - 0x6f3  :  251 - 0xfb
    "11111111", -- 1780 - 0x6f4  :  255 - 0xff
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "00111110", -- 1782 - 0x6f6  :   62 - 0x3e
    "00001100", -- 1783 - 0x6f7  :   12 - 0xc
    "00100000", -- 1784 - 0x6f8  :   32 - 0x20 -- plane 1
    "01110000", -- 1785 - 0x6f9  :  112 - 0x70
    "11110000", -- 1786 - 0x6fa  :  240 - 0xf0
    "11111000", -- 1787 - 0x6fb  :  248 - 0xf8
    "11111000", -- 1788 - 0x6fc  :  248 - 0xf8
    "11110000", -- 1789 - 0x6fd  :  240 - 0xf0
    "00110000", -- 1790 - 0x6fe  :   48 - 0x30
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0x70
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "01111001", -- 1794 - 0x702  :  121 - 0x79
    "11111001", -- 1795 - 0x703  :  249 - 0xf9
    "11110011", -- 1796 - 0x704  :  243 - 0xf3
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "01111011", -- 1798 - 0x706  :  123 - 0x7b
    "00111111", -- 1799 - 0x707  :   63 - 0x3f
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- plane 1
    "00000001", -- 1801 - 0x709  :    1 - 0x1
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00011110", -- 1805 - 0x70d  :   30 - 0x1e
    "01111111", -- 1806 - 0x70e  :  127 - 0x7f
    "00111110", -- 1807 - 0x70f  :   62 - 0x3e
    "00111111", -- 1808 - 0x710  :   63 - 0x3f -- Sprite 0x71
    "00111111", -- 1809 - 0x711  :   63 - 0x3f
    "01111011", -- 1810 - 0x712  :  123 - 0x7b
    "01111111", -- 1811 - 0x713  :  127 - 0x7f
    "11111011", -- 1812 - 0x714  :  251 - 0xfb
    "11110001", -- 1813 - 0x715  :  241 - 0xf1
    "01111001", -- 1814 - 0x716  :  121 - 0x79
    "00111000", -- 1815 - 0x717  :   56 - 0x38
    "00111100", -- 1816 - 0x718  :   60 - 0x3c -- plane 1
    "00111110", -- 1817 - 0x719  :   62 - 0x3e
    "01111111", -- 1818 - 0x71a  :  127 - 0x7f
    "01111110", -- 1819 - 0x71b  :  126 - 0x7e
    "00011000", -- 1820 - 0x71c  :   24 - 0x18
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0x72
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "10000000", -- 1826 - 0x722  :  128 - 0x80
    "10110000", -- 1827 - 0x723  :  176 - 0xb0
    "10111000", -- 1828 - 0x724  :  184 - 0xb8
    "11000110", -- 1829 - 0x725  :  198 - 0xc6
    "10010011", -- 1830 - 0x726  :  147 - 0x93
    "11110111", -- 1831 - 0x727  :  247 - 0xf7
    "11000000", -- 1832 - 0x728  :  192 - 0xc0 -- plane 1
    "11100000", -- 1833 - 0x729  :  224 - 0xe0
    "01000000", -- 1834 - 0x72a  :   64 - 0x40
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00111010", -- 1837 - 0x72d  :   58 - 0x3a
    "11101111", -- 1838 - 0x72e  :  239 - 0xef
    "01001011", -- 1839 - 0x72f  :   75 - 0x4b
    "11100011", -- 1840 - 0x730  :  227 - 0xe3 -- Sprite 0x73
    "11110111", -- 1841 - 0x731  :  247 - 0xf7
    "10010011", -- 1842 - 0x732  :  147 - 0x93
    "11000110", -- 1843 - 0x733  :  198 - 0xc6
    "10111000", -- 1844 - 0x734  :  184 - 0xb8
    "10110000", -- 1845 - 0x735  :  176 - 0xb0
    "10000000", -- 1846 - 0x736  :  128 - 0x80
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "01011111", -- 1848 - 0x738  :   95 - 0x5f -- plane 1
    "01001011", -- 1849 - 0x739  :   75 - 0x4b
    "11101111", -- 1850 - 0x73a  :  239 - 0xef
    "00111010", -- 1851 - 0x73b  :   58 - 0x3a
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "01100000", -- 1854 - 0x73e  :   96 - 0x60
    "11000000", -- 1855 - 0x73f  :  192 - 0xc0
    "00110000", -- 1856 - 0x740  :   48 - 0x30 -- Sprite 0x74
    "01111100", -- 1857 - 0x741  :  124 - 0x7c
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11011111", -- 1860 - 0x744  :  223 - 0xdf
    "00001011", -- 1861 - 0x745  :   11 - 0xb
    "00011111", -- 1862 - 0x746  :   31 - 0x1f
    "01111111", -- 1863 - 0x747  :  127 - 0x7f
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- plane 1
    "00001100", -- 1865 - 0x749  :   12 - 0xc
    "00001111", -- 1866 - 0x74a  :   15 - 0xf
    "00011111", -- 1867 - 0x74b  :   31 - 0x1f
    "00011111", -- 1868 - 0x74c  :   31 - 0x1f
    "00001111", -- 1869 - 0x74d  :   15 - 0xf
    "00001110", -- 1870 - 0x74e  :   14 - 0xe
    "00000100", -- 1871 - 0x74f  :    4 - 0x4
    "01111111", -- 1872 - 0x750  :  127 - 0x7f -- Sprite 0x75
    "00001011", -- 1873 - 0x751  :   11 - 0xb
    "00110011", -- 1874 - 0x752  :   51 - 0x33
    "00110110", -- 1875 - 0x753  :   54 - 0x36
    "00010000", -- 1876 - 0x754  :   16 - 0x10
    "00001010", -- 1877 - 0x755  :   10 - 0xa
    "00001111", -- 1878 - 0x756  :   15 - 0xf
    "00000111", -- 1879 - 0x757  :    7 - 0x7
    "10000100", -- 1880 - 0x758  :  132 - 0x84 -- plane 1
    "11000111", -- 1881 - 0x759  :  199 - 0xc7
    "01001100", -- 1882 - 0x75a  :   76 - 0x4c
    "00001001", -- 1883 - 0x75b  :    9 - 0x9
    "00001111", -- 1884 - 0x75c  :   15 - 0xf
    "00000101", -- 1885 - 0x75d  :    5 - 0x5
    "00001111", -- 1886 - 0x75e  :   15 - 0xf
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "00111000", -- 1888 - 0x760  :   56 - 0x38 -- Sprite 0x76
    "01111100", -- 1889 - 0x761  :  124 - 0x7c
    "11111100", -- 1890 - 0x762  :  252 - 0xfc
    "11111100", -- 1891 - 0x763  :  252 - 0xfc
    "11101100", -- 1892 - 0x764  :  236 - 0xec
    "10100000", -- 1893 - 0x765  :  160 - 0xa0
    "11110000", -- 1894 - 0x766  :  240 - 0xf0
    "11111100", -- 1895 - 0x767  :  252 - 0xfc
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- plane 1
    "01000000", -- 1897 - 0x769  :   64 - 0x40
    "11000000", -- 1898 - 0x76a  :  192 - 0xc0
    "11100000", -- 1899 - 0x76b  :  224 - 0xe0
    "11100000", -- 1900 - 0x76c  :  224 - 0xe0
    "11100000", -- 1901 - 0x76d  :  224 - 0xe0
    "11100000", -- 1902 - 0x76e  :  224 - 0xe0
    "01000010", -- 1903 - 0x76f  :   66 - 0x42
    "11111100", -- 1904 - 0x770  :  252 - 0xfc -- Sprite 0x77
    "10100000", -- 1905 - 0x771  :  160 - 0xa0
    "10011000", -- 1906 - 0x772  :  152 - 0x98
    "11011000", -- 1907 - 0x773  :  216 - 0xd8
    "00010000", -- 1908 - 0x774  :   16 - 0x10
    "10100000", -- 1909 - 0x775  :  160 - 0xa0
    "11100000", -- 1910 - 0x776  :  224 - 0xe0
    "11000000", -- 1911 - 0x777  :  192 - 0xc0
    "01000011", -- 1912 - 0x778  :   67 - 0x43 -- plane 1
    "11000111", -- 1913 - 0x779  :  199 - 0xc7
    "01100010", -- 1914 - 0x77a  :   98 - 0x62
    "00100000", -- 1915 - 0x77b  :   32 - 0x20
    "11100000", -- 1916 - 0x77c  :  224 - 0xe0
    "01000000", -- 1917 - 0x77d  :   64 - 0x40
    "11100000", -- 1918 - 0x77e  :  224 - 0xe0
    "11000000", -- 1919 - 0x77f  :  192 - 0xc0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0x78
    "00000001", -- 1921 - 0x781  :    1 - 0x1
    "00001101", -- 1922 - 0x782  :   13 - 0xd
    "00011101", -- 1923 - 0x783  :   29 - 0x1d
    "01100011", -- 1924 - 0x784  :   99 - 0x63
    "11001001", -- 1925 - 0x785  :  201 - 0xc9
    "11101111", -- 1926 - 0x786  :  239 - 0xef
    "11000111", -- 1927 - 0x787  :  199 - 0xc7
    "00000011", -- 1928 - 0x788  :    3 - 0x3 -- plane 1
    "00000100", -- 1929 - 0x789  :    4 - 0x4
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "01011100", -- 1932 - 0x78c  :   92 - 0x5c
    "11110111", -- 1933 - 0x78d  :  247 - 0xf7
    "11010010", -- 1934 - 0x78e  :  210 - 0xd2
    "11111010", -- 1935 - 0x78f  :  250 - 0xfa
    "11101111", -- 1936 - 0x790  :  239 - 0xef -- Sprite 0x79
    "11001001", -- 1937 - 0x791  :  201 - 0xc9
    "01100011", -- 1938 - 0x792  :   99 - 0x63
    "00011101", -- 1939 - 0x793  :   29 - 0x1d
    "00001101", -- 1940 - 0x794  :   13 - 0xd
    "00000001", -- 1941 - 0x795  :    1 - 0x1
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "11010010", -- 1944 - 0x798  :  210 - 0xd2 -- plane 1
    "11110111", -- 1945 - 0x799  :  247 - 0xf7
    "01011100", -- 1946 - 0x79a  :   92 - 0x5c
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000010", -- 1949 - 0x79d  :    2 - 0x2
    "00000111", -- 1950 - 0x79e  :    7 - 0x7
    "00000011", -- 1951 - 0x79f  :    3 - 0x3
    "00011100", -- 1952 - 0x7a0  :   28 - 0x1c -- Sprite 0x7a
    "10011110", -- 1953 - 0x7a1  :  158 - 0x9e
    "10001111", -- 1954 - 0x7a2  :  143 - 0x8f
    "11011111", -- 1955 - 0x7a3  :  223 - 0xdf
    "11111110", -- 1956 - 0x7a4  :  254 - 0xfe
    "11011110", -- 1957 - 0x7a5  :  222 - 0xde
    "11111100", -- 1958 - 0x7a6  :  252 - 0xfc
    "11111100", -- 1959 - 0x7a7  :  252 - 0xfc
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00011000", -- 1963 - 0x7ab  :   24 - 0x18
    "01111110", -- 1964 - 0x7ac  :  126 - 0x7e
    "11111110", -- 1965 - 0x7ad  :  254 - 0xfe
    "01111100", -- 1966 - 0x7ae  :  124 - 0x7c
    "00111100", -- 1967 - 0x7af  :   60 - 0x3c
    "11111100", -- 1968 - 0x7b0  :  252 - 0xfc -- Sprite 0x7b
    "11011110", -- 1969 - 0x7b1  :  222 - 0xde
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11001111", -- 1971 - 0x7b3  :  207 - 0xcf
    "10011111", -- 1972 - 0x7b4  :  159 - 0x9f
    "10011110", -- 1973 - 0x7b5  :  158 - 0x9e
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "01111100", -- 1976 - 0x7b8  :  124 - 0x7c -- plane 1
    "11111110", -- 1977 - 0x7b9  :  254 - 0xfe
    "01111000", -- 1978 - 0x7ba  :  120 - 0x78
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "10000000", -- 1982 - 0x7be  :  128 - 0x80
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00011110", -- 1988 - 0x7c4  :   30 - 0x1e
    "00111111", -- 1989 - 0x7c5  :   63 - 0x3f
    "01111101", -- 1990 - 0x7c6  :  125 - 0x7d
    "01111000", -- 1991 - 0x7c7  :  120 - 0x78
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000001", -- 1994 - 0x7ca  :    1 - 0x1
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00100000", -- 1997 - 0x7cd  :   32 - 0x20
    "01111100", -- 1998 - 0x7ce  :  124 - 0x7c
    "01111000", -- 1999 - 0x7cf  :  120 - 0x78
    "01111100", -- 2000 - 0x7d0  :  124 - 0x7c -- Sprite 0x7d
    "11111011", -- 2001 - 0x7d1  :  251 - 0xfb
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "01011111", -- 2004 - 0x7d4  :   95 - 0x5f
    "00011111", -- 2005 - 0x7d5  :   31 - 0x1f
    "00011111", -- 2006 - 0x7d6  :   31 - 0x1f
    "00011111", -- 2007 - 0x7d7  :   31 - 0x1f
    "01111100", -- 2008 - 0x7d8  :  124 - 0x7c -- plane 1
    "11111110", -- 2009 - 0x7d9  :  254 - 0xfe
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111110", -- 2011 - 0x7db  :  254 - 0xfe
    "01111100", -- 2012 - 0x7dc  :  124 - 0x7c
    "01100000", -- 2013 - 0x7dd  :   96 - 0x60
    "11100000", -- 2014 - 0x7de  :  224 - 0xe0
    "11100001", -- 2015 - 0x7df  :  225 - 0xe1
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "10000000", -- 2021 - 0x7e5  :  128 - 0x80
    "10000000", -- 2022 - 0x7e6  :  128 - 0x80
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "01111100", -- 2024 - 0x7e8  :  124 - 0x7c -- plane 1
    "10000010", -- 2025 - 0x7e9  :  130 - 0x82
    "00000001", -- 2026 - 0x7ea  :    1 - 0x1
    "10000010", -- 2027 - 0x7eb  :  130 - 0x82
    "01111100", -- 2028 - 0x7ec  :  124 - 0x7c
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0x7f
    "00100001", -- 2033 - 0x7f1  :   33 - 0x21
    "10100010", -- 2034 - 0x7f2  :  162 - 0xa2
    "10100011", -- 2035 - 0x7f3  :  163 - 0xa3
    "10110011", -- 2036 - 0x7f4  :  179 - 0xb3
    "10001111", -- 2037 - 0x7f5  :  143 - 0x8f
    "00100111", -- 2038 - 0x7f6  :   39 - 0x27
    "11111110", -- 2039 - 0x7f7  :  254 - 0xfe
    "00010000", -- 2040 - 0x7f8  :   16 - 0x10 -- plane 1
    "00011001", -- 2041 - 0x7f9  :   25 - 0x19
    "01011010", -- 2042 - 0x7fa  :   90 - 0x5a
    "11011111", -- 2043 - 0x7fb  :  223 - 0xdf
    "01001111", -- 2044 - 0x7fc  :   79 - 0x4f
    "01110011", -- 2045 - 0x7fd  :  115 - 0x73
    "11011011", -- 2046 - 0x7fe  :  219 - 0xdb
    "00000010", -- 2047 - 0x7ff  :    2 - 0x2
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Sprite 0x80
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000000", -- 2050 - 0x802  :    0 - 0x0
    "00000000", -- 2051 - 0x803  :    0 - 0x0
    "00000011", -- 2052 - 0x804  :    3 - 0x3
    "00001111", -- 2053 - 0x805  :   15 - 0xf
    "00011111", -- 2054 - 0x806  :   31 - 0x1f
    "00011111", -- 2055 - 0x807  :   31 - 0x1f
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- plane 1
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000011", -- 2059 - 0x80b  :    3 - 0x3
    "00001100", -- 2060 - 0x80c  :   12 - 0xc
    "00010000", -- 2061 - 0x80d  :   16 - 0x10
    "00100010", -- 2062 - 0x80e  :   34 - 0x22
    "00100000", -- 2063 - 0x80f  :   32 - 0x20
    "00011111", -- 2064 - 0x810  :   31 - 0x1f -- Sprite 0x81
    "00011111", -- 2065 - 0x811  :   31 - 0x1f
    "00001111", -- 2066 - 0x812  :   15 - 0xf
    "00000011", -- 2067 - 0x813  :    3 - 0x3
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00100001", -- 2072 - 0x818  :   33 - 0x21 -- plane 1
    "00100011", -- 2073 - 0x819  :   35 - 0x23
    "00010000", -- 2074 - 0x81a  :   16 - 0x10
    "00001100", -- 2075 - 0x81b  :   12 - 0xc
    "00000011", -- 2076 - 0x81c  :    3 - 0x3
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00000000", -- 2080 - 0x820  :    0 - 0x0 -- Sprite 0x82
    "00000000", -- 2081 - 0x821  :    0 - 0x0
    "00000000", -- 2082 - 0x822  :    0 - 0x0
    "00000000", -- 2083 - 0x823  :    0 - 0x0
    "11000000", -- 2084 - 0x824  :  192 - 0xc0
    "11110000", -- 2085 - 0x825  :  240 - 0xf0
    "11111000", -- 2086 - 0x826  :  248 - 0xf8
    "11111000", -- 2087 - 0x827  :  248 - 0xf8
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- plane 1
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "11000000", -- 2091 - 0x82b  :  192 - 0xc0
    "00110000", -- 2092 - 0x82c  :   48 - 0x30
    "00001000", -- 2093 - 0x82d  :    8 - 0x8
    "01100100", -- 2094 - 0x82e  :  100 - 0x64
    "11000100", -- 2095 - 0x82f  :  196 - 0xc4
    "11111000", -- 2096 - 0x830  :  248 - 0xf8 -- Sprite 0x83
    "11111000", -- 2097 - 0x831  :  248 - 0xf8
    "11110000", -- 2098 - 0x832  :  240 - 0xf0
    "11000000", -- 2099 - 0x833  :  192 - 0xc0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "10000100", -- 2104 - 0x838  :  132 - 0x84 -- plane 1
    "00000100", -- 2105 - 0x839  :    4 - 0x4
    "00001000", -- 2106 - 0x83a  :    8 - 0x8
    "00110000", -- 2107 - 0x83b  :   48 - 0x30
    "11000000", -- 2108 - 0x83c  :  192 - 0xc0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0 -- Sprite 0x84
    "00000000", -- 2113 - 0x841  :    0 - 0x0
    "00000000", -- 2114 - 0x842  :    0 - 0x0
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000011", -- 2116 - 0x844  :    3 - 0x3
    "00001111", -- 2117 - 0x845  :   15 - 0xf
    "00011111", -- 2118 - 0x846  :   31 - 0x1f
    "00011111", -- 2119 - 0x847  :   31 - 0x1f
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- plane 1
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000011", -- 2123 - 0x84b  :    3 - 0x3
    "00001100", -- 2124 - 0x84c  :   12 - 0xc
    "00010000", -- 2125 - 0x84d  :   16 - 0x10
    "00100110", -- 2126 - 0x84e  :   38 - 0x26
    "00100011", -- 2127 - 0x84f  :   35 - 0x23
    "00011111", -- 2128 - 0x850  :   31 - 0x1f -- Sprite 0x85
    "00011111", -- 2129 - 0x851  :   31 - 0x1f
    "00001111", -- 2130 - 0x852  :   15 - 0xf
    "00000011", -- 2131 - 0x853  :    3 - 0x3
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00100001", -- 2136 - 0x858  :   33 - 0x21 -- plane 1
    "00100000", -- 2137 - 0x859  :   32 - 0x20
    "00010000", -- 2138 - 0x85a  :   16 - 0x10
    "00001100", -- 2139 - 0x85b  :   12 - 0xc
    "00000011", -- 2140 - 0x85c  :    3 - 0x3
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "11000000", -- 2148 - 0x864  :  192 - 0xc0
    "11110000", -- 2149 - 0x865  :  240 - 0xf0
    "11111000", -- 2150 - 0x866  :  248 - 0xf8
    "11111000", -- 2151 - 0x867  :  248 - 0xf8
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- plane 1
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "11000000", -- 2155 - 0x86b  :  192 - 0xc0
    "00110000", -- 2156 - 0x86c  :   48 - 0x30
    "00001000", -- 2157 - 0x86d  :    8 - 0x8
    "01000100", -- 2158 - 0x86e  :   68 - 0x44
    "00000100", -- 2159 - 0x86f  :    4 - 0x4
    "11111000", -- 2160 - 0x870  :  248 - 0xf8 -- Sprite 0x87
    "11111000", -- 2161 - 0x871  :  248 - 0xf8
    "11110000", -- 2162 - 0x872  :  240 - 0xf0
    "11000000", -- 2163 - 0x873  :  192 - 0xc0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "10000100", -- 2168 - 0x878  :  132 - 0x84 -- plane 1
    "11000100", -- 2169 - 0x879  :  196 - 0xc4
    "00001000", -- 2170 - 0x87a  :    8 - 0x8
    "00110000", -- 2171 - 0x87b  :   48 - 0x30
    "11000000", -- 2172 - 0x87c  :  192 - 0xc0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Sprite 0x88
    "00000000", -- 2177 - 0x881  :    0 - 0x0
    "00000000", -- 2178 - 0x882  :    0 - 0x0
    "00000000", -- 2179 - 0x883  :    0 - 0x0
    "00000011", -- 2180 - 0x884  :    3 - 0x3
    "00001111", -- 2181 - 0x885  :   15 - 0xf
    "00011111", -- 2182 - 0x886  :   31 - 0x1f
    "00011111", -- 2183 - 0x887  :   31 - 0x1f
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000011", -- 2187 - 0x88b  :    3 - 0x3
    "00001100", -- 2188 - 0x88c  :   12 - 0xc
    "00010000", -- 2189 - 0x88d  :   16 - 0x10
    "00100000", -- 2190 - 0x88e  :   32 - 0x20
    "00100001", -- 2191 - 0x88f  :   33 - 0x21
    "00011111", -- 2192 - 0x890  :   31 - 0x1f -- Sprite 0x89
    "00011111", -- 2193 - 0x891  :   31 - 0x1f
    "00001111", -- 2194 - 0x892  :   15 - 0xf
    "00000011", -- 2195 - 0x893  :    3 - 0x3
    "00000000", -- 2196 - 0x894  :    0 - 0x0
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00100011", -- 2200 - 0x898  :   35 - 0x23 -- plane 1
    "00100110", -- 2201 - 0x899  :   38 - 0x26
    "00010000", -- 2202 - 0x89a  :   16 - 0x10
    "00001100", -- 2203 - 0x89b  :   12 - 0xc
    "00000011", -- 2204 - 0x89c  :    3 - 0x3
    "00000000", -- 2205 - 0x89d  :    0 - 0x0
    "00000000", -- 2206 - 0x89e  :    0 - 0x0
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Sprite 0x8a
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "11000000", -- 2212 - 0x8a4  :  192 - 0xc0
    "11110000", -- 2213 - 0x8a5  :  240 - 0xf0
    "11111000", -- 2214 - 0x8a6  :  248 - 0xf8
    "11111000", -- 2215 - 0x8a7  :  248 - 0xf8
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "11000000", -- 2219 - 0x8ab  :  192 - 0xc0
    "00110000", -- 2220 - 0x8ac  :   48 - 0x30
    "00001000", -- 2221 - 0x8ad  :    8 - 0x8
    "11000100", -- 2222 - 0x8ae  :  196 - 0xc4
    "10000100", -- 2223 - 0x8af  :  132 - 0x84
    "11111000", -- 2224 - 0x8b0  :  248 - 0xf8 -- Sprite 0x8b
    "11111000", -- 2225 - 0x8b1  :  248 - 0xf8
    "11110000", -- 2226 - 0x8b2  :  240 - 0xf0
    "11000000", -- 2227 - 0x8b3  :  192 - 0xc0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "00000000", -- 2230 - 0x8b6  :    0 - 0x0
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00000100", -- 2232 - 0x8b8  :    4 - 0x4 -- plane 1
    "01000100", -- 2233 - 0x8b9  :   68 - 0x44
    "00001000", -- 2234 - 0x8ba  :    8 - 0x8
    "00110000", -- 2235 - 0x8bb  :   48 - 0x30
    "11000000", -- 2236 - 0x8bc  :  192 - 0xc0
    "00000000", -- 2237 - 0x8bd  :    0 - 0x0
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Sprite 0x8c
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000011", -- 2244 - 0x8c4  :    3 - 0x3
    "00001111", -- 2245 - 0x8c5  :   15 - 0xf
    "00011111", -- 2246 - 0x8c6  :   31 - 0x1f
    "00011111", -- 2247 - 0x8c7  :   31 - 0x1f
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000011", -- 2251 - 0x8cb  :    3 - 0x3
    "00001100", -- 2252 - 0x8cc  :   12 - 0xc
    "00010000", -- 2253 - 0x8cd  :   16 - 0x10
    "00100011", -- 2254 - 0x8ce  :   35 - 0x23
    "00100001", -- 2255 - 0x8cf  :   33 - 0x21
    "00011111", -- 2256 - 0x8d0  :   31 - 0x1f -- Sprite 0x8d
    "00011111", -- 2257 - 0x8d1  :   31 - 0x1f
    "00001111", -- 2258 - 0x8d2  :   15 - 0xf
    "00000011", -- 2259 - 0x8d3  :    3 - 0x3
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00100000", -- 2264 - 0x8d8  :   32 - 0x20 -- plane 1
    "00100010", -- 2265 - 0x8d9  :   34 - 0x22
    "00010000", -- 2266 - 0x8da  :   16 - 0x10
    "00001100", -- 2267 - 0x8db  :   12 - 0xc
    "00000011", -- 2268 - 0x8dc  :    3 - 0x3
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000000", -- 2270 - 0x8de  :    0 - 0x0
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Sprite 0x8e
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "11000000", -- 2276 - 0x8e4  :  192 - 0xc0
    "11110000", -- 2277 - 0x8e5  :  240 - 0xf0
    "11111000", -- 2278 - 0x8e6  :  248 - 0xf8
    "11111000", -- 2279 - 0x8e7  :  248 - 0xf8
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "11000000", -- 2283 - 0x8eb  :  192 - 0xc0
    "00110000", -- 2284 - 0x8ec  :   48 - 0x30
    "00001000", -- 2285 - 0x8ed  :    8 - 0x8
    "00000100", -- 2286 - 0x8ee  :    4 - 0x4
    "10000100", -- 2287 - 0x8ef  :  132 - 0x84
    "11111000", -- 2288 - 0x8f0  :  248 - 0xf8 -- Sprite 0x8f
    "11111000", -- 2289 - 0x8f1  :  248 - 0xf8
    "11110000", -- 2290 - 0x8f2  :  240 - 0xf0
    "11000000", -- 2291 - 0x8f3  :  192 - 0xc0
    "00000000", -- 2292 - 0x8f4  :    0 - 0x0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "11000100", -- 2296 - 0x8f8  :  196 - 0xc4 -- plane 1
    "01100100", -- 2297 - 0x8f9  :  100 - 0x64
    "00001000", -- 2298 - 0x8fa  :    8 - 0x8
    "00110000", -- 2299 - 0x8fb  :   48 - 0x30
    "11000000", -- 2300 - 0x8fc  :  192 - 0xc0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00001111", -- 2307 - 0x903  :   15 - 0xf
    "00110000", -- 2308 - 0x904  :   48 - 0x30
    "01100000", -- 2309 - 0x905  :   96 - 0x60
    "00111111", -- 2310 - 0x906  :   63 - 0x3f
    "01111111", -- 2311 - 0x907  :  127 - 0x7f
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- plane 1
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00101111", -- 2316 - 0x90c  :   47 - 0x2f
    "00111111", -- 2317 - 0x90d  :   63 - 0x3f
    "01100000", -- 2318 - 0x90e  :   96 - 0x60
    "00100000", -- 2319 - 0x90f  :   32 - 0x20
    "01111111", -- 2320 - 0x910  :  127 - 0x7f -- Sprite 0x91
    "00111111", -- 2321 - 0x911  :   63 - 0x3f
    "01100000", -- 2322 - 0x912  :   96 - 0x60
    "00110000", -- 2323 - 0x913  :   48 - 0x30
    "00001111", -- 2324 - 0x914  :   15 - 0xf
    "00000000", -- 2325 - 0x915  :    0 - 0x0
    "00000000", -- 2326 - 0x916  :    0 - 0x0
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "00100000", -- 2328 - 0x918  :   32 - 0x20 -- plane 1
    "01100000", -- 2329 - 0x919  :   96 - 0x60
    "00111111", -- 2330 - 0x91a  :   63 - 0x3f
    "00101111", -- 2331 - 0x91b  :   47 - 0x2f
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Sprite 0x92
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "11111000", -- 2339 - 0x923  :  248 - 0xf8
    "00000110", -- 2340 - 0x924  :    6 - 0x6
    "00000011", -- 2341 - 0x925  :    3 - 0x3
    "11111110", -- 2342 - 0x926  :  254 - 0xfe
    "11111111", -- 2343 - 0x927  :  255 - 0xff
    "00000000", -- 2344 - 0x928  :    0 - 0x0 -- plane 1
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "11111010", -- 2348 - 0x92c  :  250 - 0xfa
    "11111110", -- 2349 - 0x92d  :  254 - 0xfe
    "00000011", -- 2350 - 0x92e  :    3 - 0x3
    "00000010", -- 2351 - 0x92f  :    2 - 0x2
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Sprite 0x93
    "11111110", -- 2353 - 0x931  :  254 - 0xfe
    "00000011", -- 2354 - 0x932  :    3 - 0x3
    "00000110", -- 2355 - 0x933  :    6 - 0x6
    "11111000", -- 2356 - 0x934  :  248 - 0xf8
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000010", -- 2360 - 0x938  :    2 - 0x2 -- plane 1
    "00000011", -- 2361 - 0x939  :    3 - 0x3
    "11111110", -- 2362 - 0x93a  :  254 - 0xfe
    "11111010", -- 2363 - 0x93b  :  250 - 0xfa
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00101111", -- 2372 - 0x944  :   47 - 0x2f
    "00111111", -- 2373 - 0x945  :   63 - 0x3f
    "01100000", -- 2374 - 0x946  :   96 - 0x60
    "00100000", -- 2375 - 0x947  :   32 - 0x20
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- plane 1
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00001111", -- 2379 - 0x94b  :   15 - 0xf
    "00110000", -- 2380 - 0x94c  :   48 - 0x30
    "01100000", -- 2381 - 0x94d  :   96 - 0x60
    "00111111", -- 2382 - 0x94e  :   63 - 0x3f
    "01111111", -- 2383 - 0x94f  :  127 - 0x7f
    "00100000", -- 2384 - 0x950  :   32 - 0x20 -- Sprite 0x95
    "01100000", -- 2385 - 0x951  :   96 - 0x60
    "00111111", -- 2386 - 0x952  :   63 - 0x3f
    "00101111", -- 2387 - 0x953  :   47 - 0x2f
    "00000000", -- 2388 - 0x954  :    0 - 0x0
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "00000000", -- 2391 - 0x957  :    0 - 0x0
    "01111111", -- 2392 - 0x958  :  127 - 0x7f -- plane 1
    "00111111", -- 2393 - 0x959  :   63 - 0x3f
    "01100000", -- 2394 - 0x95a  :   96 - 0x60
    "00110000", -- 2395 - 0x95b  :   48 - 0x30
    "00001111", -- 2396 - 0x95c  :   15 - 0xf
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "11111010", -- 2404 - 0x964  :  250 - 0xfa
    "11111110", -- 2405 - 0x965  :  254 - 0xfe
    "00000011", -- 2406 - 0x966  :    3 - 0x3
    "00000010", -- 2407 - 0x967  :    2 - 0x2
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- plane 1
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "00000000", -- 2410 - 0x96a  :    0 - 0x0
    "11111000", -- 2411 - 0x96b  :  248 - 0xf8
    "00000110", -- 2412 - 0x96c  :    6 - 0x6
    "00000011", -- 2413 - 0x96d  :    3 - 0x3
    "11111110", -- 2414 - 0x96e  :  254 - 0xfe
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00000010", -- 2416 - 0x970  :    2 - 0x2 -- Sprite 0x97
    "00000011", -- 2417 - 0x971  :    3 - 0x3
    "11111110", -- 2418 - 0x972  :  254 - 0xfe
    "11111010", -- 2419 - 0x973  :  250 - 0xfa
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "11111111", -- 2424 - 0x978  :  255 - 0xff -- plane 1
    "11111110", -- 2425 - 0x979  :  254 - 0xfe
    "00000011", -- 2426 - 0x97a  :    3 - 0x3
    "00000110", -- 2427 - 0x97b  :    6 - 0x6
    "11111000", -- 2428 - 0x97c  :  248 - 0xf8
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Sprite 0x98
    "01000100", -- 2433 - 0x981  :   68 - 0x44
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "01000001", -- 2435 - 0x983  :   65 - 0x41
    "00100000", -- 2436 - 0x984  :   32 - 0x20
    "01001011", -- 2437 - 0x985  :   75 - 0x4b
    "00100111", -- 2438 - 0x986  :   39 - 0x27
    "00011111", -- 2439 - 0x987  :   31 - 0x1f
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- plane 1
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "01000000", -- 2443 - 0x98b  :   64 - 0x40
    "00100000", -- 2444 - 0x98c  :   32 - 0x20
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000001", -- 2447 - 0x98f  :    1 - 0x1
    "00001111", -- 2448 - 0x990  :   15 - 0xf -- Sprite 0x99
    "00011110", -- 2449 - 0x991  :   30 - 0x1e
    "00011111", -- 2450 - 0x992  :   31 - 0x1f
    "00011111", -- 2451 - 0x993  :   31 - 0x1f
    "00011111", -- 2452 - 0x994  :   31 - 0x1f
    "00001111", -- 2453 - 0x995  :   15 - 0xf
    "00001111", -- 2454 - 0x996  :   15 - 0xf
    "00000011", -- 2455 - 0x997  :    3 - 0x3
    "00000011", -- 2456 - 0x998  :    3 - 0x3 -- plane 1
    "00000111", -- 2457 - 0x999  :    7 - 0x7
    "00000110", -- 2458 - 0x99a  :    6 - 0x6
    "00000110", -- 2459 - 0x99b  :    6 - 0x6
    "00000111", -- 2460 - 0x99c  :    7 - 0x7
    "00000011", -- 2461 - 0x99d  :    3 - 0x3
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Sprite 0x9a
    "00100000", -- 2465 - 0x9a1  :   32 - 0x20
    "01010000", -- 2466 - 0x9a2  :   80 - 0x50
    "00100000", -- 2467 - 0x9a3  :   32 - 0x20
    "01100000", -- 2468 - 0x9a4  :   96 - 0x60
    "01001000", -- 2469 - 0x9a5  :   72 - 0x48
    "11100000", -- 2470 - 0x9a6  :  224 - 0xe0
    "11110000", -- 2471 - 0x9a7  :  240 - 0xf0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "01000000", -- 2474 - 0x9aa  :   64 - 0x40
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00001000", -- 2477 - 0x9ad  :    8 - 0x8
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "01000000", -- 2479 - 0x9af  :   64 - 0x40
    "11111000", -- 2480 - 0x9b0  :  248 - 0xf8 -- Sprite 0x9b
    "01111000", -- 2481 - 0x9b1  :  120 - 0x78
    "00111100", -- 2482 - 0x9b2  :   60 - 0x3c
    "00111100", -- 2483 - 0x9b3  :   60 - 0x3c
    "00111100", -- 2484 - 0x9b4  :   60 - 0x3c
    "11111100", -- 2485 - 0x9b5  :  252 - 0xfc
    "11111000", -- 2486 - 0x9b6  :  248 - 0xf8
    "11100000", -- 2487 - 0x9b7  :  224 - 0xe0
    "11100000", -- 2488 - 0x9b8  :  224 - 0xe0 -- plane 1
    "11110000", -- 2489 - 0x9b9  :  240 - 0xf0
    "11010000", -- 2490 - 0x9ba  :  208 - 0xd0
    "11010000", -- 2491 - 0x9bb  :  208 - 0xd0
    "11110000", -- 2492 - 0x9bc  :  240 - 0xf0
    "11100000", -- 2493 - 0x9bd  :  224 - 0xe0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00010000", -- 2496 - 0x9c0  :   16 - 0x10 -- Sprite 0x9c
    "00000001", -- 2497 - 0x9c1  :    1 - 0x1
    "00101010", -- 2498 - 0x9c2  :   42 - 0x2a
    "00001100", -- 2499 - 0x9c3  :   12 - 0xc
    "10100110", -- 2500 - 0x9c4  :  166 - 0xa6
    "00010111", -- 2501 - 0x9c5  :   23 - 0x17
    "00011111", -- 2502 - 0x9c6  :   31 - 0x1f
    "00011111", -- 2503 - 0x9c7  :   31 - 0x1f
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- plane 1
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000010", -- 2506 - 0x9ca  :    2 - 0x2
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "10000000", -- 2508 - 0x9cc  :  128 - 0x80
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000011", -- 2510 - 0x9ce  :    3 - 0x3
    "00000111", -- 2511 - 0x9cf  :    7 - 0x7
    "01011110", -- 2512 - 0x9d0  :   94 - 0x5e -- Sprite 0x9d
    "00111100", -- 2513 - 0x9d1  :   60 - 0x3c
    "00111101", -- 2514 - 0x9d2  :   61 - 0x3d
    "00111101", -- 2515 - 0x9d3  :   61 - 0x3d
    "00111110", -- 2516 - 0x9d4  :   62 - 0x3e
    "00011111", -- 2517 - 0x9d5  :   31 - 0x1f
    "00001111", -- 2518 - 0x9d6  :   15 - 0xf
    "00000111", -- 2519 - 0x9d7  :    7 - 0x7
    "00000111", -- 2520 - 0x9d8  :    7 - 0x7 -- plane 1
    "00001111", -- 2521 - 0x9d9  :   15 - 0xf
    "00001110", -- 2522 - 0x9da  :   14 - 0xe
    "00001110", -- 2523 - 0x9db  :   14 - 0xe
    "00001111", -- 2524 - 0x9dc  :   15 - 0xf
    "00000111", -- 2525 - 0x9dd  :    7 - 0x7
    "00000011", -- 2526 - 0x9de  :    3 - 0x3
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Sprite 0x9e
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "10000000", -- 2530 - 0x9e2  :  128 - 0x80
    "11001000", -- 2531 - 0x9e3  :  200 - 0xc8
    "01100000", -- 2532 - 0x9e4  :   96 - 0x60
    "11100000", -- 2533 - 0x9e5  :  224 - 0xe0
    "11110100", -- 2534 - 0x9e6  :  244 - 0xf4
    "11111000", -- 2535 - 0x9e7  :  248 - 0xf8
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00001000", -- 2539 - 0x9eb  :    8 - 0x8
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "10000000", -- 2541 - 0x9ed  :  128 - 0x80
    "00100100", -- 2542 - 0x9ee  :   36 - 0x24
    "11000000", -- 2543 - 0x9ef  :  192 - 0xc0
    "01111100", -- 2544 - 0x9f0  :  124 - 0x7c -- Sprite 0x9f
    "00011100", -- 2545 - 0x9f1  :   28 - 0x1c
    "00101110", -- 2546 - 0x9f2  :   46 - 0x2e
    "00101110", -- 2547 - 0x9f3  :   46 - 0x2e
    "00011110", -- 2548 - 0x9f4  :   30 - 0x1e
    "11111100", -- 2549 - 0x9f5  :  252 - 0xfc
    "11111000", -- 2550 - 0x9f6  :  248 - 0xf8
    "11100000", -- 2551 - 0x9f7  :  224 - 0xe0
    "11110000", -- 2552 - 0x9f8  :  240 - 0xf0 -- plane 1
    "11111000", -- 2553 - 0x9f9  :  248 - 0xf8
    "11011000", -- 2554 - 0x9fa  :  216 - 0xd8
    "11011000", -- 2555 - 0x9fb  :  216 - 0xd8
    "11111000", -- 2556 - 0x9fc  :  248 - 0xf8
    "11110000", -- 2557 - 0x9fd  :  240 - 0xf0
    "11000000", -- 2558 - 0x9fe  :  192 - 0xc0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "11111111", -- 2560 - 0xa00  :  255 - 0xff -- Sprite 0xa0
    "11111111", -- 2561 - 0xa01  :  255 - 0xff
    "00111000", -- 2562 - 0xa02  :   56 - 0x38
    "01101100", -- 2563 - 0xa03  :  108 - 0x6c
    "11000110", -- 2564 - 0xa04  :  198 - 0xc6
    "10000011", -- 2565 - 0xa05  :  131 - 0x83
    "11111111", -- 2566 - 0xa06  :  255 - 0xff
    "11111111", -- 2567 - 0xa07  :  255 - 0xff
    "11111111", -- 2568 - 0xa08  :  255 - 0xff -- plane 1
    "11111111", -- 2569 - 0xa09  :  255 - 0xff
    "00111000", -- 2570 - 0xa0a  :   56 - 0x38
    "01101100", -- 2571 - 0xa0b  :  108 - 0x6c
    "11000110", -- 2572 - 0xa0c  :  198 - 0xc6
    "10000011", -- 2573 - 0xa0d  :  131 - 0x83
    "11111111", -- 2574 - 0xa0e  :  255 - 0xff
    "11111111", -- 2575 - 0xa0f  :  255 - 0xff
    "11111111", -- 2576 - 0xa10  :  255 - 0xff -- Sprite 0xa1
    "11111111", -- 2577 - 0xa11  :  255 - 0xff
    "00111000", -- 2578 - 0xa12  :   56 - 0x38
    "01101100", -- 2579 - 0xa13  :  108 - 0x6c
    "11000110", -- 2580 - 0xa14  :  198 - 0xc6
    "10000011", -- 2581 - 0xa15  :  131 - 0x83
    "11111111", -- 2582 - 0xa16  :  255 - 0xff
    "11111111", -- 2583 - 0xa17  :  255 - 0xff
    "11111111", -- 2584 - 0xa18  :  255 - 0xff -- plane 1
    "11111111", -- 2585 - 0xa19  :  255 - 0xff
    "00111000", -- 2586 - 0xa1a  :   56 - 0x38
    "01101100", -- 2587 - 0xa1b  :  108 - 0x6c
    "11000110", -- 2588 - 0xa1c  :  198 - 0xc6
    "10000011", -- 2589 - 0xa1d  :  131 - 0x83
    "11111111", -- 2590 - 0xa1e  :  255 - 0xff
    "11111111", -- 2591 - 0xa1f  :  255 - 0xff
    "10010010", -- 2592 - 0xa20  :  146 - 0x92 -- Sprite 0xa2
    "01010100", -- 2593 - 0xa21  :   84 - 0x54
    "00111000", -- 2594 - 0xa22  :   56 - 0x38
    "11111110", -- 2595 - 0xa23  :  254 - 0xfe
    "00111000", -- 2596 - 0xa24  :   56 - 0x38
    "01010100", -- 2597 - 0xa25  :   84 - 0x54
    "10010010", -- 2598 - 0xa26  :  146 - 0x92
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- plane 1
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "11111111", -- 2608 - 0xa30  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 2609 - 0xa31  :  255 - 0xff
    "11111111", -- 2610 - 0xa32  :  255 - 0xff
    "11111111", -- 2611 - 0xa33  :  255 - 0xff
    "11111111", -- 2612 - 0xa34  :  255 - 0xff
    "11111111", -- 2613 - 0xa35  :  255 - 0xff
    "11111111", -- 2614 - 0xa36  :  255 - 0xff
    "11111111", -- 2615 - 0xa37  :  255 - 0xff
    "11111111", -- 2616 - 0xa38  :  255 - 0xff -- plane 1
    "11111111", -- 2617 - 0xa39  :  255 - 0xff
    "11111111", -- 2618 - 0xa3a  :  255 - 0xff
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "11111111", -- 2624 - 0xa40  :  255 - 0xff -- Sprite 0xa4
    "11111111", -- 2625 - 0xa41  :  255 - 0xff
    "11111111", -- 2626 - 0xa42  :  255 - 0xff
    "11111111", -- 2627 - 0xa43  :  255 - 0xff
    "11111111", -- 2628 - 0xa44  :  255 - 0xff
    "11111111", -- 2629 - 0xa45  :  255 - 0xff
    "11111111", -- 2630 - 0xa46  :  255 - 0xff
    "11111111", -- 2631 - 0xa47  :  255 - 0xff
    "11111111", -- 2632 - 0xa48  :  255 - 0xff -- plane 1
    "11111111", -- 2633 - 0xa49  :  255 - 0xff
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11111111", -- 2635 - 0xa4b  :  255 - 0xff
    "11111111", -- 2636 - 0xa4c  :  255 - 0xff
    "11111111", -- 2637 - 0xa4d  :  255 - 0xff
    "11111111", -- 2638 - 0xa4e  :  255 - 0xff
    "11111111", -- 2639 - 0xa4f  :  255 - 0xff
    "11111111", -- 2640 - 0xa50  :  255 - 0xff -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "11111111", -- 2643 - 0xa53  :  255 - 0xff
    "11111111", -- 2644 - 0xa54  :  255 - 0xff
    "11111111", -- 2645 - 0xa55  :  255 - 0xff
    "11111111", -- 2646 - 0xa56  :  255 - 0xff
    "11111111", -- 2647 - 0xa57  :  255 - 0xff
    "11111111", -- 2648 - 0xa58  :  255 - 0xff -- plane 1
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "11111111", -- 2652 - 0xa5c  :  255 - 0xff
    "11111111", -- 2653 - 0xa5d  :  255 - 0xff
    "11111111", -- 2654 - 0xa5e  :  255 - 0xff
    "11111111", -- 2655 - 0xa5f  :  255 - 0xff
    "11111111", -- 2656 - 0xa60  :  255 - 0xff -- Sprite 0xa6
    "11111111", -- 2657 - 0xa61  :  255 - 0xff
    "11111111", -- 2658 - 0xa62  :  255 - 0xff
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "11111111", -- 2660 - 0xa64  :  255 - 0xff
    "11111111", -- 2661 - 0xa65  :  255 - 0xff
    "11111111", -- 2662 - 0xa66  :  255 - 0xff
    "11111111", -- 2663 - 0xa67  :  255 - 0xff
    "11111111", -- 2664 - 0xa68  :  255 - 0xff -- plane 1
    "11111111", -- 2665 - 0xa69  :  255 - 0xff
    "11111111", -- 2666 - 0xa6a  :  255 - 0xff
    "11111111", -- 2667 - 0xa6b  :  255 - 0xff
    "11111111", -- 2668 - 0xa6c  :  255 - 0xff
    "11111111", -- 2669 - 0xa6d  :  255 - 0xff
    "11111111", -- 2670 - 0xa6e  :  255 - 0xff
    "11111111", -- 2671 - 0xa6f  :  255 - 0xff
    "11111111", -- 2672 - 0xa70  :  255 - 0xff -- Sprite 0xa7
    "11111111", -- 2673 - 0xa71  :  255 - 0xff
    "11111111", -- 2674 - 0xa72  :  255 - 0xff
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111111", -- 2676 - 0xa74  :  255 - 0xff
    "11111111", -- 2677 - 0xa75  :  255 - 0xff
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "11111111", -- 2680 - 0xa78  :  255 - 0xff -- plane 1
    "11111111", -- 2681 - 0xa79  :  255 - 0xff
    "11111111", -- 2682 - 0xa7a  :  255 - 0xff
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111111", -- 2684 - 0xa7c  :  255 - 0xff
    "11111111", -- 2685 - 0xa7d  :  255 - 0xff
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00100011", -- 2693 - 0xa85  :   35 - 0x23
    "10010111", -- 2694 - 0xa86  :  151 - 0x97
    "00101111", -- 2695 - 0xa87  :   47 - 0x2f
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- plane 1
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000001", -- 2702 - 0xa8e  :    1 - 0x1
    "00000011", -- 2703 - 0xa8f  :    3 - 0x3
    "01101110", -- 2704 - 0xa90  :  110 - 0x6e -- Sprite 0xa9
    "11101111", -- 2705 - 0xa91  :  239 - 0xef
    "11110111", -- 2706 - 0xa92  :  247 - 0xf7
    "11111111", -- 2707 - 0xa93  :  255 - 0xff
    "01111111", -- 2708 - 0xa94  :  127 - 0x7f
    "00111111", -- 2709 - 0xa95  :   63 - 0x3f
    "01011111", -- 2710 - 0xa96  :   95 - 0x5f
    "00001111", -- 2711 - 0xa97  :   15 - 0xf
    "00000111", -- 2712 - 0xa98  :    7 - 0x7 -- plane 1
    "00000111", -- 2713 - 0xa99  :    7 - 0x7
    "00000011", -- 2714 - 0xa9a  :    3 - 0x3
    "00100111", -- 2715 - 0xa9b  :   39 - 0x27
    "00011111", -- 2716 - 0xa9c  :   31 - 0x1f
    "00000111", -- 2717 - 0xa9d  :    7 - 0x7
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "11111000", -- 2724 - 0xaa4  :  248 - 0xf8
    "11111100", -- 2725 - 0xaa5  :  252 - 0xfc
    "11111110", -- 2726 - 0xaa6  :  254 - 0xfe
    "01011110", -- 2727 - 0xaa7  :   94 - 0x5e
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- plane 1
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "11110000", -- 2733 - 0xaad  :  240 - 0xf0
    "11111000", -- 2734 - 0xaae  :  248 - 0xf8
    "10101100", -- 2735 - 0xaaf  :  172 - 0xac
    "01011110", -- 2736 - 0xab0  :   94 - 0x5e -- Sprite 0xab
    "00001100", -- 2737 - 0xab1  :   12 - 0xc
    "10011110", -- 2738 - 0xab2  :  158 - 0x9e
    "11111110", -- 2739 - 0xab3  :  254 - 0xfe
    "11111110", -- 2740 - 0xab4  :  254 - 0xfe
    "11111110", -- 2741 - 0xab5  :  254 - 0xfe
    "11111000", -- 2742 - 0xab6  :  248 - 0xf8
    "11000000", -- 2743 - 0xab7  :  192 - 0xc0
    "10101100", -- 2744 - 0xab8  :  172 - 0xac -- plane 1
    "11111000", -- 2745 - 0xab9  :  248 - 0xf8
    "11111000", -- 2746 - 0xaba  :  248 - 0xf8
    "11111000", -- 2747 - 0xabb  :  248 - 0xf8
    "11110000", -- 2748 - 0xabc  :  240 - 0xf0
    "11000000", -- 2749 - 0xabd  :  192 - 0xc0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000011", -- 2757 - 0xac5  :    3 - 0x3
    "00000111", -- 2758 - 0xac6  :    7 - 0x7
    "00101111", -- 2759 - 0xac7  :   47 - 0x2f
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- plane 1
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000001", -- 2766 - 0xace  :    1 - 0x1
    "00000011", -- 2767 - 0xacf  :    3 - 0x3
    "01001110", -- 2768 - 0xad0  :   78 - 0x4e -- Sprite 0xad
    "01101110", -- 2769 - 0xad1  :  110 - 0x6e
    "11111110", -- 2770 - 0xad2  :  254 - 0xfe
    "01111111", -- 2771 - 0xad3  :  127 - 0x7f
    "00111111", -- 2772 - 0xad4  :   63 - 0x3f
    "00011111", -- 2773 - 0xad5  :   31 - 0x1f
    "00001111", -- 2774 - 0xad6  :   15 - 0xf
    "00000011", -- 2775 - 0xad7  :    3 - 0x3
    "00000111", -- 2776 - 0xad8  :    7 - 0x7 -- plane 1
    "00000111", -- 2777 - 0xad9  :    7 - 0x7
    "00000111", -- 2778 - 0xada  :    7 - 0x7
    "00100111", -- 2779 - 0xadb  :   39 - 0x27
    "00011111", -- 2780 - 0xadc  :   31 - 0x1f
    "00000111", -- 2781 - 0xadd  :    7 - 0x7
    "00000001", -- 2782 - 0xade  :    1 - 0x1
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000000", -- 2786 - 0xae2  :    0 - 0x0
    "00000000", -- 2787 - 0xae3  :    0 - 0x0
    "11111000", -- 2788 - 0xae4  :  248 - 0xf8
    "11111100", -- 2789 - 0xae5  :  252 - 0xfc
    "11111110", -- 2790 - 0xae6  :  254 - 0xfe
    "01010110", -- 2791 - 0xae7  :   86 - 0x56
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- plane 1
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "11110000", -- 2797 - 0xaed  :  240 - 0xf0
    "11111000", -- 2798 - 0xaee  :  248 - 0xf8
    "10101100", -- 2799 - 0xaef  :  172 - 0xac
    "01010110", -- 2800 - 0xaf0  :   86 - 0x56 -- Sprite 0xaf
    "00001100", -- 2801 - 0xaf1  :   12 - 0xc
    "00001110", -- 2802 - 0xaf2  :   14 - 0xe
    "00011111", -- 2803 - 0xaf3  :   31 - 0x1f
    "11111111", -- 2804 - 0xaf4  :  255 - 0xff
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111110", -- 2806 - 0xaf6  :  254 - 0xfe
    "11111000", -- 2807 - 0xaf7  :  248 - 0xf8
    "10101100", -- 2808 - 0xaf8  :  172 - 0xac -- plane 1
    "11111000", -- 2809 - 0xaf9  :  248 - 0xf8
    "11111000", -- 2810 - 0xafa  :  248 - 0xf8
    "11111100", -- 2811 - 0xafb  :  252 - 0xfc
    "11111100", -- 2812 - 0xafc  :  252 - 0xfc
    "11111000", -- 2813 - 0xafd  :  248 - 0xf8
    "11110000", -- 2814 - 0xafe  :  240 - 0xf0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "11111111", -- 2816 - 0xb00  :  255 - 0xff -- Sprite 0xb0
    "11111111", -- 2817 - 0xb01  :  255 - 0xff
    "11111111", -- 2818 - 0xb02  :  255 - 0xff
    "11111111", -- 2819 - 0xb03  :  255 - 0xff
    "11111111", -- 2820 - 0xb04  :  255 - 0xff
    "11111111", -- 2821 - 0xb05  :  255 - 0xff
    "11111111", -- 2822 - 0xb06  :  255 - 0xff
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "11111111", -- 2824 - 0xb08  :  255 - 0xff -- plane 1
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11111111", -- 2826 - 0xb0a  :  255 - 0xff
    "11111111", -- 2827 - 0xb0b  :  255 - 0xff
    "11111111", -- 2828 - 0xb0c  :  255 - 0xff
    "11111111", -- 2829 - 0xb0d  :  255 - 0xff
    "11111111", -- 2830 - 0xb0e  :  255 - 0xff
    "11111111", -- 2831 - 0xb0f  :  255 - 0xff
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Sprite 0xb1
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "11111111", -- 2834 - 0xb12  :  255 - 0xff
    "11111111", -- 2835 - 0xb13  :  255 - 0xff
    "11111111", -- 2836 - 0xb14  :  255 - 0xff
    "11111111", -- 2837 - 0xb15  :  255 - 0xff
    "11111111", -- 2838 - 0xb16  :  255 - 0xff
    "11111111", -- 2839 - 0xb17  :  255 - 0xff
    "11111111", -- 2840 - 0xb18  :  255 - 0xff -- plane 1
    "11111111", -- 2841 - 0xb19  :  255 - 0xff
    "11111111", -- 2842 - 0xb1a  :  255 - 0xff
    "11111111", -- 2843 - 0xb1b  :  255 - 0xff
    "11111111", -- 2844 - 0xb1c  :  255 - 0xff
    "11111111", -- 2845 - 0xb1d  :  255 - 0xff
    "11111111", -- 2846 - 0xb1e  :  255 - 0xff
    "11111111", -- 2847 - 0xb1f  :  255 - 0xff
    "11111111", -- 2848 - 0xb20  :  255 - 0xff -- Sprite 0xb2
    "11111111", -- 2849 - 0xb21  :  255 - 0xff
    "11111111", -- 2850 - 0xb22  :  255 - 0xff
    "11111111", -- 2851 - 0xb23  :  255 - 0xff
    "11111111", -- 2852 - 0xb24  :  255 - 0xff
    "11111111", -- 2853 - 0xb25  :  255 - 0xff
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "11111111", -- 2855 - 0xb27  :  255 - 0xff
    "11111111", -- 2856 - 0xb28  :  255 - 0xff -- plane 1
    "11111111", -- 2857 - 0xb29  :  255 - 0xff
    "11111111", -- 2858 - 0xb2a  :  255 - 0xff
    "11111111", -- 2859 - 0xb2b  :  255 - 0xff
    "11111111", -- 2860 - 0xb2c  :  255 - 0xff
    "11111111", -- 2861 - 0xb2d  :  255 - 0xff
    "11111111", -- 2862 - 0xb2e  :  255 - 0xff
    "11111111", -- 2863 - 0xb2f  :  255 - 0xff
    "11111111", -- 2864 - 0xb30  :  255 - 0xff -- Sprite 0xb3
    "11111111", -- 2865 - 0xb31  :  255 - 0xff
    "11111111", -- 2866 - 0xb32  :  255 - 0xff
    "11111111", -- 2867 - 0xb33  :  255 - 0xff
    "11111111", -- 2868 - 0xb34  :  255 - 0xff
    "11111111", -- 2869 - 0xb35  :  255 - 0xff
    "11111111", -- 2870 - 0xb36  :  255 - 0xff
    "11111111", -- 2871 - 0xb37  :  255 - 0xff
    "11111111", -- 2872 - 0xb38  :  255 - 0xff -- plane 1
    "11111111", -- 2873 - 0xb39  :  255 - 0xff
    "11111111", -- 2874 - 0xb3a  :  255 - 0xff
    "11111111", -- 2875 - 0xb3b  :  255 - 0xff
    "11111111", -- 2876 - 0xb3c  :  255 - 0xff
    "11111111", -- 2877 - 0xb3d  :  255 - 0xff
    "11111111", -- 2878 - 0xb3e  :  255 - 0xff
    "11111111", -- 2879 - 0xb3f  :  255 - 0xff
    "11111111", -- 2880 - 0xb40  :  255 - 0xff -- Sprite 0xb4
    "11111111", -- 2881 - 0xb41  :  255 - 0xff
    "11111111", -- 2882 - 0xb42  :  255 - 0xff
    "11111111", -- 2883 - 0xb43  :  255 - 0xff
    "11111111", -- 2884 - 0xb44  :  255 - 0xff
    "11111111", -- 2885 - 0xb45  :  255 - 0xff
    "11111111", -- 2886 - 0xb46  :  255 - 0xff
    "11111111", -- 2887 - 0xb47  :  255 - 0xff
    "11111111", -- 2888 - 0xb48  :  255 - 0xff -- plane 1
    "11111111", -- 2889 - 0xb49  :  255 - 0xff
    "11111111", -- 2890 - 0xb4a  :  255 - 0xff
    "11111111", -- 2891 - 0xb4b  :  255 - 0xff
    "11111111", -- 2892 - 0xb4c  :  255 - 0xff
    "11111111", -- 2893 - 0xb4d  :  255 - 0xff
    "11111111", -- 2894 - 0xb4e  :  255 - 0xff
    "11111111", -- 2895 - 0xb4f  :  255 - 0xff
    "11111111", -- 2896 - 0xb50  :  255 - 0xff -- Sprite 0xb5
    "11111111", -- 2897 - 0xb51  :  255 - 0xff
    "11111111", -- 2898 - 0xb52  :  255 - 0xff
    "11111111", -- 2899 - 0xb53  :  255 - 0xff
    "11111111", -- 2900 - 0xb54  :  255 - 0xff
    "11111111", -- 2901 - 0xb55  :  255 - 0xff
    "11111111", -- 2902 - 0xb56  :  255 - 0xff
    "11111111", -- 2903 - 0xb57  :  255 - 0xff
    "11111111", -- 2904 - 0xb58  :  255 - 0xff -- plane 1
    "11111111", -- 2905 - 0xb59  :  255 - 0xff
    "11111111", -- 2906 - 0xb5a  :  255 - 0xff
    "11111111", -- 2907 - 0xb5b  :  255 - 0xff
    "11111111", -- 2908 - 0xb5c  :  255 - 0xff
    "11111111", -- 2909 - 0xb5d  :  255 - 0xff
    "11111111", -- 2910 - 0xb5e  :  255 - 0xff
    "11111111", -- 2911 - 0xb5f  :  255 - 0xff
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Sprite 0xb6
    "11111111", -- 2913 - 0xb61  :  255 - 0xff
    "11111111", -- 2914 - 0xb62  :  255 - 0xff
    "11111111", -- 2915 - 0xb63  :  255 - 0xff
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11111111", -- 2917 - 0xb65  :  255 - 0xff
    "11111111", -- 2918 - 0xb66  :  255 - 0xff
    "11111111", -- 2919 - 0xb67  :  255 - 0xff
    "11111111", -- 2920 - 0xb68  :  255 - 0xff -- plane 1
    "11111111", -- 2921 - 0xb69  :  255 - 0xff
    "11111111", -- 2922 - 0xb6a  :  255 - 0xff
    "11111111", -- 2923 - 0xb6b  :  255 - 0xff
    "11111111", -- 2924 - 0xb6c  :  255 - 0xff
    "11111111", -- 2925 - 0xb6d  :  255 - 0xff
    "11111111", -- 2926 - 0xb6e  :  255 - 0xff
    "11111111", -- 2927 - 0xb6f  :  255 - 0xff
    "11111111", -- 2928 - 0xb70  :  255 - 0xff -- Sprite 0xb7
    "11111111", -- 2929 - 0xb71  :  255 - 0xff
    "11111111", -- 2930 - 0xb72  :  255 - 0xff
    "11111111", -- 2931 - 0xb73  :  255 - 0xff
    "11111111", -- 2932 - 0xb74  :  255 - 0xff
    "11111111", -- 2933 - 0xb75  :  255 - 0xff
    "11111111", -- 2934 - 0xb76  :  255 - 0xff
    "11111111", -- 2935 - 0xb77  :  255 - 0xff
    "11111111", -- 2936 - 0xb78  :  255 - 0xff -- plane 1
    "11111111", -- 2937 - 0xb79  :  255 - 0xff
    "11111111", -- 2938 - 0xb7a  :  255 - 0xff
    "11111111", -- 2939 - 0xb7b  :  255 - 0xff
    "11111111", -- 2940 - 0xb7c  :  255 - 0xff
    "11111111", -- 2941 - 0xb7d  :  255 - 0xff
    "11111111", -- 2942 - 0xb7e  :  255 - 0xff
    "11111111", -- 2943 - 0xb7f  :  255 - 0xff
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Sprite 0xb8
    "00000111", -- 2945 - 0xb81  :    7 - 0x7
    "00001000", -- 2946 - 0xb82  :    8 - 0x8
    "00010000", -- 2947 - 0xb83  :   16 - 0x10
    "00010000", -- 2948 - 0xb84  :   16 - 0x10
    "00100000", -- 2949 - 0xb85  :   32 - 0x20
    "00100000", -- 2950 - 0xb86  :   32 - 0x20
    "00100000", -- 2951 - 0xb87  :   32 - 0x20
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- plane 1
    "00000111", -- 2953 - 0xb89  :    7 - 0x7
    "00001000", -- 2954 - 0xb8a  :    8 - 0x8
    "00010000", -- 2955 - 0xb8b  :   16 - 0x10
    "00010000", -- 2956 - 0xb8c  :   16 - 0x10
    "00100000", -- 2957 - 0xb8d  :   32 - 0x20
    "00100000", -- 2958 - 0xb8e  :   32 - 0x20
    "00100000", -- 2959 - 0xb8f  :   32 - 0x20
    "00011111", -- 2960 - 0xb90  :   31 - 0x1f -- Sprite 0xb9
    "00101111", -- 2961 - 0xb91  :   47 - 0x2f
    "00110111", -- 2962 - 0xb92  :   55 - 0x37
    "00111010", -- 2963 - 0xb93  :   58 - 0x3a
    "00111101", -- 2964 - 0xb94  :   61 - 0x3d
    "00111110", -- 2965 - 0xb95  :   62 - 0x3e
    "00111111", -- 2966 - 0xb96  :   63 - 0x3f
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00011111", -- 2968 - 0xb98  :   31 - 0x1f -- plane 1
    "00111111", -- 2969 - 0xb99  :   63 - 0x3f
    "00111111", -- 2970 - 0xb9a  :   63 - 0x3f
    "00111111", -- 2971 - 0xb9b  :   63 - 0x3f
    "00111110", -- 2972 - 0xb9c  :   62 - 0x3e
    "00111111", -- 2973 - 0xb9d  :   63 - 0x3f
    "00111111", -- 2974 - 0xb9e  :   63 - 0x3f
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Sprite 0xba
    "00000101", -- 2977 - 0xba1  :    5 - 0x5
    "00011001", -- 2978 - 0xba2  :   25 - 0x19
    "00110011", -- 2979 - 0xba3  :   51 - 0x33
    "01100011", -- 2980 - 0xba4  :   99 - 0x63
    "11000111", -- 2981 - 0xba5  :  199 - 0xc7
    "11000111", -- 2982 - 0xba6  :  199 - 0xc7
    "11000100", -- 2983 - 0xba7  :  196 - 0xc4
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- plane 1
    "00000111", -- 2985 - 0xba9  :    7 - 0x7
    "00011111", -- 2986 - 0xbaa  :   31 - 0x1f
    "00111111", -- 2987 - 0xbab  :   63 - 0x3f
    "01111111", -- 2988 - 0xbac  :  127 - 0x7f
    "11111111", -- 2989 - 0xbad  :  255 - 0xff
    "11111111", -- 2990 - 0xbae  :  255 - 0xff
    "11011101", -- 2991 - 0xbaf  :  221 - 0xdd
    "10000000", -- 2992 - 0xbb0  :  128 - 0x80 -- Sprite 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000011", -- 2997 - 0xbb5  :    3 - 0x3
    "00000011", -- 2998 - 0xbb6  :    3 - 0x3
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "10001001", -- 3000 - 0xbb8  :  137 - 0x89 -- plane 1
    "00000001", -- 3001 - 0xbb9  :    1 - 0x1
    "00000001", -- 3002 - 0xbba  :    1 - 0x1
    "00000001", -- 3003 - 0xbbb  :    1 - 0x1
    "00000001", -- 3004 - 0xbbc  :    1 - 0x1
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Sprite 0xbc
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000011", -- 3022 - 0xbce  :    3 - 0x3
    "00000111", -- 3023 - 0xbcf  :    7 - 0x7
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00001111", -- 3026 - 0xbd2  :   15 - 0xf
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "10000000", -- 3028 - 0xbd4  :  128 - 0x80
    "01100011", -- 3029 - 0xbd5  :   99 - 0x63
    "00011110", -- 3030 - 0xbd6  :   30 - 0x1e
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00001111", -- 3032 - 0xbd8  :   15 - 0xf -- plane 1
    "00001111", -- 3033 - 0xbd9  :   15 - 0xf
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00011111", -- 3035 - 0xbdb  :   31 - 0x1f
    "01111111", -- 3036 - 0xbdc  :  127 - 0x7f
    "00011100", -- 3037 - 0xbdd  :   28 - 0x1c
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000001", -- 3040 - 0xbe0  :    1 - 0x1 -- Sprite 0xbe
    "00000011", -- 3041 - 0xbe1  :    3 - 0x3
    "00011001", -- 3042 - 0xbe2  :   25 - 0x19
    "00111100", -- 3043 - 0xbe3  :   60 - 0x3c
    "00011001", -- 3044 - 0xbe4  :   25 - 0x19
    "00100011", -- 3045 - 0xbe5  :   35 - 0x23
    "01010001", -- 3046 - 0xbe6  :   81 - 0x51
    "00100000", -- 3047 - 0xbe7  :   32 - 0x20
    "00000001", -- 3048 - 0xbe8  :    1 - 0x1 -- plane 1
    "00000010", -- 3049 - 0xbe9  :    2 - 0x2
    "00011001", -- 3050 - 0xbea  :   25 - 0x19
    "00100100", -- 3051 - 0xbeb  :   36 - 0x24
    "00011001", -- 3052 - 0xbec  :   25 - 0x19
    "00100010", -- 3053 - 0xbed  :   34 - 0x22
    "00010001", -- 3054 - 0xbee  :   17 - 0x11
    "00101100", -- 3055 - 0xbef  :   44 - 0x2c
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00011111", -- 3064 - 0xbf8  :   31 - 0x1f -- plane 1
    "00000111", -- 3065 - 0xbf9  :    7 - 0x7
    "00000011", -- 3066 - 0xbfa  :    3 - 0x3
    "00000011", -- 3067 - 0xbfb  :    3 - 0x3
    "00000001", -- 3068 - 0xbfc  :    1 - 0x1
    "00000001", -- 3069 - 0xbfd  :    1 - 0x1
    "00000001", -- 3070 - 0xbfe  :    1 - 0x1
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Sprite 0xc0
    "00111111", -- 3073 - 0xc01  :   63 - 0x3f
    "00011111", -- 3074 - 0xc02  :   31 - 0x1f
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000001", -- 3076 - 0xc04  :    1 - 0x1
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "00000001", -- 3078 - 0xc06  :    1 - 0x1
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- plane 1
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000001", -- 3083 - 0xc0b  :    1 - 0x1
    "00000011", -- 3084 - 0xc0c  :    3 - 0x3
    "00000111", -- 3085 - 0xc0d  :    7 - 0x7
    "00001101", -- 3086 - 0xc0e  :   13 - 0xd
    "00011001", -- 3087 - 0xc0f  :   25 - 0x19
    "00010001", -- 3088 - 0xc10  :   17 - 0x11 -- Sprite 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000001", -- 3090 - 0xc12  :    1 - 0x1
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000001", -- 3092 - 0xc14  :    1 - 0x1
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00011111", -- 3094 - 0xc16  :   31 - 0x1f
    "00111111", -- 3095 - 0xc17  :   63 - 0x3f
    "00101001", -- 3096 - 0xc18  :   41 - 0x29 -- plane 1
    "00011001", -- 3097 - 0xc19  :   25 - 0x19
    "00001101", -- 3098 - 0xc1a  :   13 - 0xd
    "00000111", -- 3099 - 0xc1b  :    7 - 0x7
    "00000011", -- 3100 - 0xc1c  :    3 - 0x3
    "00000001", -- 3101 - 0xc1d  :    1 - 0x1
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Sprite 0xc2
    "11111100", -- 3105 - 0xc21  :  252 - 0xfc
    "11111000", -- 3106 - 0xc22  :  248 - 0xf8
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "10000000", -- 3108 - 0xc24  :  128 - 0x80
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "10000000", -- 3110 - 0xc26  :  128 - 0x80
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- plane 1
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "10000000", -- 3115 - 0xc2b  :  128 - 0x80
    "11000000", -- 3116 - 0xc2c  :  192 - 0xc0
    "11100000", -- 3117 - 0xc2d  :  224 - 0xe0
    "10110000", -- 3118 - 0xc2e  :  176 - 0xb0
    "10011000", -- 3119 - 0xc2f  :  152 - 0x98
    "10001000", -- 3120 - 0xc30  :  136 - 0x88 -- Sprite 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "10000000", -- 3122 - 0xc32  :  128 - 0x80
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "10000000", -- 3124 - 0xc34  :  128 - 0x80
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "11111000", -- 3126 - 0xc36  :  248 - 0xf8
    "11111100", -- 3127 - 0xc37  :  252 - 0xfc
    "10010100", -- 3128 - 0xc38  :  148 - 0x94 -- plane 1
    "10011000", -- 3129 - 0xc39  :  152 - 0x98
    "10110000", -- 3130 - 0xc3a  :  176 - 0xb0
    "11100000", -- 3131 - 0xc3b  :  224 - 0xe0
    "11000000", -- 3132 - 0xc3c  :  192 - 0xc0
    "10000000", -- 3133 - 0xc3d  :  128 - 0x80
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00111111", -- 3141 - 0xc45  :   63 - 0x3f
    "00011111", -- 3142 - 0xc46  :   31 - 0x1f
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0 -- plane 1
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000001", -- 3151 - 0xc4f  :    1 - 0x1
    "00000001", -- 3152 - 0xc50  :    1 - 0x1 -- Sprite 0xc5
    "00000001", -- 3153 - 0xc51  :    1 - 0x1
    "01000001", -- 3154 - 0xc52  :   65 - 0x41
    "00000001", -- 3155 - 0xc53  :    1 - 0x1
    "00000001", -- 3156 - 0xc54  :    1 - 0x1
    "00000000", -- 3157 - 0xc55  :    0 - 0x0
    "00011111", -- 3158 - 0xc56  :   31 - 0x1f
    "00111111", -- 3159 - 0xc57  :   63 - 0x3f
    "00001111", -- 3160 - 0xc58  :   15 - 0xf -- plane 1
    "01111001", -- 3161 - 0xc59  :  121 - 0x79
    "10100001", -- 3162 - 0xc5a  :  161 - 0xa1
    "01111001", -- 3163 - 0xc5b  :  121 - 0x79
    "00001111", -- 3164 - 0xc5c  :   15 - 0xf
    "00000001", -- 3165 - 0xc5d  :    1 - 0x1
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "11111100", -- 3173 - 0xc65  :  252 - 0xfc
    "11111000", -- 3174 - 0xc66  :  248 - 0xf8
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0 -- plane 1
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "00000000", -- 3181 - 0xc6d  :    0 - 0x0
    "00000000", -- 3182 - 0xc6e  :    0 - 0x0
    "10000000", -- 3183 - 0xc6f  :  128 - 0x80
    "10000000", -- 3184 - 0xc70  :  128 - 0x80 -- Sprite 0xc7
    "10000000", -- 3185 - 0xc71  :  128 - 0x80
    "10000010", -- 3186 - 0xc72  :  130 - 0x82
    "10000000", -- 3187 - 0xc73  :  128 - 0x80
    "10000000", -- 3188 - 0xc74  :  128 - 0x80
    "00000000", -- 3189 - 0xc75  :    0 - 0x0
    "11111000", -- 3190 - 0xc76  :  248 - 0xf8
    "11111100", -- 3191 - 0xc77  :  252 - 0xfc
    "11110000", -- 3192 - 0xc78  :  240 - 0xf0 -- plane 1
    "10011110", -- 3193 - 0xc79  :  158 - 0x9e
    "10000101", -- 3194 - 0xc7a  :  133 - 0x85
    "10011110", -- 3195 - 0xc7b  :  158 - 0x9e
    "11110000", -- 3196 - 0xc7c  :  240 - 0xf0
    "10000000", -- 3197 - 0xc7d  :  128 - 0x80
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00011110", -- 3203 - 0xc83  :   30 - 0x1e
    "00111111", -- 3204 - 0xc84  :   63 - 0x3f
    "00111111", -- 3205 - 0xc85  :   63 - 0x3f
    "00111111", -- 3206 - 0xc86  :   63 - 0x3f
    "00111111", -- 3207 - 0xc87  :   63 - 0x3f
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- plane 1
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00011110", -- 3211 - 0xc8b  :   30 - 0x1e
    "00111111", -- 3212 - 0xc8c  :   63 - 0x3f
    "00111111", -- 3213 - 0xc8d  :   63 - 0x3f
    "00111111", -- 3214 - 0xc8e  :   63 - 0x3f
    "00111111", -- 3215 - 0xc8f  :   63 - 0x3f
    "00011111", -- 3216 - 0xc90  :   31 - 0x1f -- Sprite 0xc9
    "00001111", -- 3217 - 0xc91  :   15 - 0xf
    "00000111", -- 3218 - 0xc92  :    7 - 0x7
    "00000011", -- 3219 - 0xc93  :    3 - 0x3
    "00000001", -- 3220 - 0xc94  :    1 - 0x1
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00011111", -- 3224 - 0xc98  :   31 - 0x1f -- plane 1
    "00001111", -- 3225 - 0xc99  :   15 - 0xf
    "00000111", -- 3226 - 0xc9a  :    7 - 0x7
    "00000011", -- 3227 - 0xc9b  :    3 - 0x3
    "00000001", -- 3228 - 0xc9c  :    1 - 0x1
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00111100", -- 3235 - 0xca3  :   60 - 0x3c
    "01111110", -- 3236 - 0xca4  :  126 - 0x7e
    "11111110", -- 3237 - 0xca5  :  254 - 0xfe
    "11111110", -- 3238 - 0xca6  :  254 - 0xfe
    "11111110", -- 3239 - 0xca7  :  254 - 0xfe
    "00000000", -- 3240 - 0xca8  :    0 - 0x0 -- plane 1
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00111100", -- 3243 - 0xcab  :   60 - 0x3c
    "01111110", -- 3244 - 0xcac  :  126 - 0x7e
    "11111110", -- 3245 - 0xcad  :  254 - 0xfe
    "11111110", -- 3246 - 0xcae  :  254 - 0xfe
    "11111110", -- 3247 - 0xcaf  :  254 - 0xfe
    "11111100", -- 3248 - 0xcb0  :  252 - 0xfc -- Sprite 0xcb
    "11111000", -- 3249 - 0xcb1  :  248 - 0xf8
    "11110000", -- 3250 - 0xcb2  :  240 - 0xf0
    "11100000", -- 3251 - 0xcb3  :  224 - 0xe0
    "11000000", -- 3252 - 0xcb4  :  192 - 0xc0
    "10000000", -- 3253 - 0xcb5  :  128 - 0x80
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "11111100", -- 3256 - 0xcb8  :  252 - 0xfc -- plane 1
    "11111000", -- 3257 - 0xcb9  :  248 - 0xf8
    "11110000", -- 3258 - 0xcba  :  240 - 0xf0
    "11100000", -- 3259 - 0xcbb  :  224 - 0xe0
    "11000000", -- 3260 - 0xcbc  :  192 - 0xc0
    "10000000", -- 3261 - 0xcbd  :  128 - 0x80
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff -- Sprite 0xcc
    "11111111", -- 3265 - 0xcc1  :  255 - 0xff
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111111", -- 3267 - 0xcc3  :  255 - 0xff
    "11111111", -- 3268 - 0xcc4  :  255 - 0xff
    "11111111", -- 3269 - 0xcc5  :  255 - 0xff
    "11111111", -- 3270 - 0xcc6  :  255 - 0xff
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "11111111", -- 3272 - 0xcc8  :  255 - 0xff -- plane 1
    "11111111", -- 3273 - 0xcc9  :  255 - 0xff
    "11111111", -- 3274 - 0xcca  :  255 - 0xff
    "11111111", -- 3275 - 0xccb  :  255 - 0xff
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "11111111", -- 3277 - 0xccd  :  255 - 0xff
    "11111111", -- 3278 - 0xcce  :  255 - 0xff
    "11111111", -- 3279 - 0xccf  :  255 - 0xff
    "11111111", -- 3280 - 0xcd0  :  255 - 0xff -- Sprite 0xcd
    "11111111", -- 3281 - 0xcd1  :  255 - 0xff
    "11111111", -- 3282 - 0xcd2  :  255 - 0xff
    "11111111", -- 3283 - 0xcd3  :  255 - 0xff
    "11111111", -- 3284 - 0xcd4  :  255 - 0xff
    "11111111", -- 3285 - 0xcd5  :  255 - 0xff
    "11111111", -- 3286 - 0xcd6  :  255 - 0xff
    "11111111", -- 3287 - 0xcd7  :  255 - 0xff
    "11111111", -- 3288 - 0xcd8  :  255 - 0xff -- plane 1
    "11111111", -- 3289 - 0xcd9  :  255 - 0xff
    "11111111", -- 3290 - 0xcda  :  255 - 0xff
    "11111111", -- 3291 - 0xcdb  :  255 - 0xff
    "11111111", -- 3292 - 0xcdc  :  255 - 0xff
    "11111111", -- 3293 - 0xcdd  :  255 - 0xff
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "11111111", -- 3296 - 0xce0  :  255 - 0xff -- Sprite 0xce
    "11111111", -- 3297 - 0xce1  :  255 - 0xff
    "11111111", -- 3298 - 0xce2  :  255 - 0xff
    "11111111", -- 3299 - 0xce3  :  255 - 0xff
    "11111111", -- 3300 - 0xce4  :  255 - 0xff
    "11111111", -- 3301 - 0xce5  :  255 - 0xff
    "11111111", -- 3302 - 0xce6  :  255 - 0xff
    "11111111", -- 3303 - 0xce7  :  255 - 0xff
    "11111111", -- 3304 - 0xce8  :  255 - 0xff -- plane 1
    "11111111", -- 3305 - 0xce9  :  255 - 0xff
    "11111111", -- 3306 - 0xcea  :  255 - 0xff
    "11111111", -- 3307 - 0xceb  :  255 - 0xff
    "11111111", -- 3308 - 0xcec  :  255 - 0xff
    "11111111", -- 3309 - 0xced  :  255 - 0xff
    "11111111", -- 3310 - 0xcee  :  255 - 0xff
    "11111111", -- 3311 - 0xcef  :  255 - 0xff
    "11111111", -- 3312 - 0xcf0  :  255 - 0xff -- Sprite 0xcf
    "11111111", -- 3313 - 0xcf1  :  255 - 0xff
    "11111111", -- 3314 - 0xcf2  :  255 - 0xff
    "11111111", -- 3315 - 0xcf3  :  255 - 0xff
    "11111111", -- 3316 - 0xcf4  :  255 - 0xff
    "11111111", -- 3317 - 0xcf5  :  255 - 0xff
    "11111111", -- 3318 - 0xcf6  :  255 - 0xff
    "11111111", -- 3319 - 0xcf7  :  255 - 0xff
    "11111111", -- 3320 - 0xcf8  :  255 - 0xff -- plane 1
    "11111111", -- 3321 - 0xcf9  :  255 - 0xff
    "11111111", -- 3322 - 0xcfa  :  255 - 0xff
    "11111111", -- 3323 - 0xcfb  :  255 - 0xff
    "11111111", -- 3324 - 0xcfc  :  255 - 0xff
    "11111111", -- 3325 - 0xcfd  :  255 - 0xff
    "11111111", -- 3326 - 0xcfe  :  255 - 0xff
    "11111111", -- 3327 - 0xcff  :  255 - 0xff
    "00001000", -- 3328 - 0xd00  :    8 - 0x8 -- Sprite 0xd0
    "00011001", -- 3329 - 0xd01  :   25 - 0x19
    "00001001", -- 3330 - 0xd02  :    9 - 0x9
    "00001001", -- 3331 - 0xd03  :    9 - 0x9
    "00001001", -- 3332 - 0xd04  :    9 - 0x9
    "00001001", -- 3333 - 0xd05  :    9 - 0x9
    "00011100", -- 3334 - 0xd06  :   28 - 0x1c
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- plane 1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00111000", -- 3344 - 0xd10  :   56 - 0x38 -- Sprite 0xd1
    "00000101", -- 3345 - 0xd11  :    5 - 0x5
    "00000101", -- 3346 - 0xd12  :    5 - 0x5
    "00011001", -- 3347 - 0xd13  :   25 - 0x19
    "00000101", -- 3348 - 0xd14  :    5 - 0x5
    "00000101", -- 3349 - 0xd15  :    5 - 0x5
    "00111000", -- 3350 - 0xd16  :   56 - 0x38
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0 -- plane 1
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00111100", -- 3360 - 0xd20  :   60 - 0x3c -- Sprite 0xd2
    "00100001", -- 3361 - 0xd21  :   33 - 0x21
    "00100001", -- 3362 - 0xd22  :   33 - 0x21
    "00111101", -- 3363 - 0xd23  :   61 - 0x3d
    "00000101", -- 3364 - 0xd24  :    5 - 0x5
    "00000101", -- 3365 - 0xd25  :    5 - 0x5
    "00111000", -- 3366 - 0xd26  :   56 - 0x38
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- plane 1
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000000", -- 3372 - 0xd2c  :    0 - 0x0
    "00000000", -- 3373 - 0xd2d  :    0 - 0x0
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00011000", -- 3376 - 0xd30  :   24 - 0x18 -- Sprite 0xd3
    "00100101", -- 3377 - 0xd31  :   37 - 0x25
    "00100101", -- 3378 - 0xd32  :   37 - 0x25
    "00011001", -- 3379 - 0xd33  :   25 - 0x19
    "00100101", -- 3380 - 0xd34  :   37 - 0x25
    "00100101", -- 3381 - 0xd35  :   37 - 0x25
    "00011000", -- 3382 - 0xd36  :   24 - 0x18
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "00000000", -- 3384 - 0xd38  :    0 - 0x0 -- plane 1
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "00000000", -- 3386 - 0xd3a  :    0 - 0x0
    "00000000", -- 3387 - 0xd3b  :    0 - 0x0
    "00000000", -- 3388 - 0xd3c  :    0 - 0x0
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "11000110", -- 3392 - 0xd40  :  198 - 0xc6 -- Sprite 0xd4
    "00101001", -- 3393 - 0xd41  :   41 - 0x29
    "00101001", -- 3394 - 0xd42  :   41 - 0x29
    "00101001", -- 3395 - 0xd43  :   41 - 0x29
    "00101001", -- 3396 - 0xd44  :   41 - 0x29
    "00101001", -- 3397 - 0xd45  :   41 - 0x29
    "11000110", -- 3398 - 0xd46  :  198 - 0xc6
    "00000000", -- 3399 - 0xd47  :    0 - 0x0
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- plane 1
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- plane 1
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000001", -- 3419 - 0xd5b  :    1 - 0x1
    "00000011", -- 3420 - 0xd5c  :    3 - 0x3
    "01100011", -- 3421 - 0xd5d  :   99 - 0x63
    "00110001", -- 3422 - 0xd5e  :   49 - 0x31
    "00011111", -- 3423 - 0xd5f  :   31 - 0x1f
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "00000000", -- 3427 - 0xd63  :    0 - 0x0
    "00111100", -- 3428 - 0xd64  :   60 - 0x3c
    "10110110", -- 3429 - 0xd65  :  182 - 0xb6
    "01111100", -- 3430 - 0xd66  :  124 - 0x7c
    "11111000", -- 3431 - 0xd67  :  248 - 0xf8
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- plane 1
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "11111100", -- 3434 - 0xd6a  :  252 - 0xfc
    "11111110", -- 3435 - 0xd6b  :  254 - 0xfe
    "11000000", -- 3436 - 0xd6c  :  192 - 0xc0
    "01000000", -- 3437 - 0xd6d  :   64 - 0x40
    "10000000", -- 3438 - 0xd6e  :  128 - 0x80
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "00000011", -- 3440 - 0xd70  :    3 - 0x3 -- Sprite 0xd7
    "00000011", -- 3441 - 0xd71  :    3 - 0x3
    "00000011", -- 3442 - 0xd72  :    3 - 0x3
    "00000111", -- 3443 - 0xd73  :    7 - 0x7
    "00001100", -- 3444 - 0xd74  :   12 - 0xc
    "00011011", -- 3445 - 0xd75  :   27 - 0x1b
    "01110111", -- 3446 - 0xd76  :  119 - 0x77
    "00000111", -- 3447 - 0xd77  :    7 - 0x7
    "01111111", -- 3448 - 0xd78  :  127 - 0x7f -- plane 1
    "00111111", -- 3449 - 0xd79  :   63 - 0x3f
    "01010011", -- 3450 - 0xd7a  :   83 - 0x53
    "00000111", -- 3451 - 0xd7b  :    7 - 0x7
    "00001100", -- 3452 - 0xd7c  :   12 - 0xc
    "00011011", -- 3453 - 0xd7d  :   27 - 0x1b
    "00000111", -- 3454 - 0xd7e  :    7 - 0x7
    "00000111", -- 3455 - 0xd7f  :    7 - 0x7
    "00001111", -- 3456 - 0xd80  :   15 - 0xf -- Sprite 0xd8
    "00001111", -- 3457 - 0xd81  :   15 - 0xf
    "00011111", -- 3458 - 0xd82  :   31 - 0x1f
    "00111111", -- 3459 - 0xd83  :   63 - 0x3f
    "01111111", -- 3460 - 0xd84  :  127 - 0x7f
    "00111111", -- 3461 - 0xd85  :   63 - 0x3f
    "00000000", -- 3462 - 0xd86  :    0 - 0x0
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00001111", -- 3464 - 0xd88  :   15 - 0xf -- plane 1
    "00001111", -- 3465 - 0xd89  :   15 - 0xf
    "00000011", -- 3466 - 0xd8a  :    3 - 0x3
    "00111000", -- 3467 - 0xd8b  :   56 - 0x38
    "00111111", -- 3468 - 0xd8c  :   63 - 0x3f
    "00001110", -- 3469 - 0xd8d  :   14 - 0xe
    "00011100", -- 3470 - 0xd8e  :   28 - 0x1c
    "00001110", -- 3471 - 0xd8f  :   14 - 0xe
    "11100000", -- 3472 - 0xd90  :  224 - 0xe0 -- Sprite 0xd9
    "11110000", -- 3473 - 0xd91  :  240 - 0xf0
    "11110000", -- 3474 - 0xd92  :  240 - 0xf0
    "11110000", -- 3475 - 0xd93  :  240 - 0xf0
    "00011000", -- 3476 - 0xd94  :   24 - 0x18
    "11111100", -- 3477 - 0xd95  :  252 - 0xfc
    "11111100", -- 3478 - 0xd96  :  252 - 0xfc
    "11111100", -- 3479 - 0xd97  :  252 - 0xfc
    "00000000", -- 3480 - 0xd98  :    0 - 0x0 -- plane 1
    "10010000", -- 3481 - 0xd99  :  144 - 0x90
    "11110000", -- 3482 - 0xd9a  :  240 - 0xf0
    "11110000", -- 3483 - 0xd9b  :  240 - 0xf0
    "00011000", -- 3484 - 0xd9c  :   24 - 0x18
    "11111100", -- 3485 - 0xd9d  :  252 - 0xfc
    "11110000", -- 3486 - 0xd9e  :  240 - 0xf0
    "11111000", -- 3487 - 0xd9f  :  248 - 0xf8
    "11111000", -- 3488 - 0xda0  :  248 - 0xf8 -- Sprite 0xda
    "11111100", -- 3489 - 0xda1  :  252 - 0xfc
    "11111111", -- 3490 - 0xda2  :  255 - 0xff
    "11111111", -- 3491 - 0xda3  :  255 - 0xff
    "11111110", -- 3492 - 0xda4  :  254 - 0xfe
    "11110000", -- 3493 - 0xda5  :  240 - 0xf0
    "00000000", -- 3494 - 0xda6  :    0 - 0x0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "11111000", -- 3496 - 0xda8  :  248 - 0xf8 -- plane 1
    "11110000", -- 3497 - 0xda9  :  240 - 0xf0
    "10000111", -- 3498 - 0xdaa  :  135 - 0x87
    "00111101", -- 3499 - 0xdab  :   61 - 0x3d
    "11111110", -- 3500 - 0xdac  :  254 - 0xfe
    "00011100", -- 3501 - 0xdad  :   28 - 0x1c
    "00001000", -- 3502 - 0xdae  :    8 - 0x8
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000011", -- 3504 - 0xdb0  :    3 - 0x3 -- Sprite 0xdb
    "00000011", -- 3505 - 0xdb1  :    3 - 0x3
    "00000011", -- 3506 - 0xdb2  :    3 - 0x3
    "00000011", -- 3507 - 0xdb3  :    3 - 0x3
    "00000001", -- 3508 - 0xdb4  :    1 - 0x1
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000111", -- 3510 - 0xdb6  :    7 - 0x7
    "00011111", -- 3511 - 0xdb7  :   31 - 0x1f
    "01111111", -- 3512 - 0xdb8  :  127 - 0x7f -- plane 1
    "00111111", -- 3513 - 0xdb9  :   63 - 0x3f
    "01010011", -- 3514 - 0xdba  :   83 - 0x53
    "00000011", -- 3515 - 0xdbb  :    3 - 0x3
    "00000001", -- 3516 - 0xdbc  :    1 - 0x1
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000111", -- 3518 - 0xdbe  :    7 - 0x7
    "00011111", -- 3519 - 0xdbf  :   31 - 0x1f
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Sprite 0xdc
    "11111111", -- 3521 - 0xdc1  :  255 - 0xff
    "01111111", -- 3522 - 0xdc2  :  127 - 0x7f
    "00111111", -- 3523 - 0xdc3  :   63 - 0x3f
    "00001111", -- 3524 - 0xdc4  :   15 - 0xf
    "00000011", -- 3525 - 0xdc5  :    3 - 0x3
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "11001111", -- 3528 - 0xdc8  :  207 - 0xcf -- plane 1
    "01100011", -- 3529 - 0xdc9  :   99 - 0x63
    "00111000", -- 3530 - 0xdca  :   56 - 0x38
    "00111110", -- 3531 - 0xdcb  :   62 - 0x3e
    "01111011", -- 3532 - 0xdcc  :  123 - 0x7b
    "00110000", -- 3533 - 0xdcd  :   48 - 0x30
    "00011000", -- 3534 - 0xdce  :   24 - 0x18
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "11100000", -- 3536 - 0xdd0  :  224 - 0xe0 -- Sprite 0xdd
    "11110000", -- 3537 - 0xdd1  :  240 - 0xf0
    "11110000", -- 3538 - 0xdd2  :  240 - 0xf0
    "11100000", -- 3539 - 0xdd3  :  224 - 0xe0
    "11111110", -- 3540 - 0xdd4  :  254 - 0xfe
    "00111100", -- 3541 - 0xdd5  :   60 - 0x3c
    "11110000", -- 3542 - 0xdd6  :  240 - 0xf0
    "11111100", -- 3543 - 0xdd7  :  252 - 0xfc
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0 -- plane 1
    "10010000", -- 3545 - 0xdd9  :  144 - 0x90
    "11110000", -- 3546 - 0xdda  :  240 - 0xf0
    "11100000", -- 3547 - 0xddb  :  224 - 0xe0
    "11111000", -- 3548 - 0xddc  :  248 - 0xf8
    "00111000", -- 3549 - 0xddd  :   56 - 0x38
    "11110000", -- 3550 - 0xdde  :  240 - 0xf0
    "11110000", -- 3551 - 0xddf  :  240 - 0xf0
    "11111100", -- 3552 - 0xde0  :  252 - 0xfc -- Sprite 0xde
    "11111000", -- 3553 - 0xde1  :  248 - 0xf8
    "11111000", -- 3554 - 0xde2  :  248 - 0xf8
    "11111000", -- 3555 - 0xde3  :  248 - 0xf8
    "11111000", -- 3556 - 0xde4  :  248 - 0xf8
    "11111000", -- 3557 - 0xde5  :  248 - 0xf8
    "11111000", -- 3558 - 0xde6  :  248 - 0xf8
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "11111000", -- 3560 - 0xde8  :  248 - 0xf8 -- plane 1
    "11111000", -- 3561 - 0xde9  :  248 - 0xf8
    "11111000", -- 3562 - 0xdea  :  248 - 0xf8
    "00111000", -- 3563 - 0xdeb  :   56 - 0x38
    "10000000", -- 3564 - 0xdec  :  128 - 0x80
    "11111000", -- 3565 - 0xded  :  248 - 0xf8
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "01011100", -- 3567 - 0xdef  :   92 - 0x5c
    "11111111", -- 3568 - 0xdf0  :  255 - 0xff -- Sprite 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "11111111", -- 3570 - 0xdf2  :  255 - 0xff
    "11111111", -- 3571 - 0xdf3  :  255 - 0xff
    "11111111", -- 3572 - 0xdf4  :  255 - 0xff
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111111", -- 3575 - 0xdf7  :  255 - 0xff
    "11111111", -- 3576 - 0xdf8  :  255 - 0xff -- plane 1
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11111111", -- 3580 - 0xdfc  :  255 - 0xff
    "11111111", -- 3581 - 0xdfd  :  255 - 0xff
    "11111111", -- 3582 - 0xdfe  :  255 - 0xff
    "11111111", -- 3583 - 0xdff  :  255 - 0xff
    "11111111", -- 3584 - 0xe00  :  255 - 0xff -- Sprite 0xe0
    "11111111", -- 3585 - 0xe01  :  255 - 0xff
    "11111111", -- 3586 - 0xe02  :  255 - 0xff
    "11111111", -- 3587 - 0xe03  :  255 - 0xff
    "11111111", -- 3588 - 0xe04  :  255 - 0xff
    "11111111", -- 3589 - 0xe05  :  255 - 0xff
    "11111111", -- 3590 - 0xe06  :  255 - 0xff
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "11111111", -- 3592 - 0xe08  :  255 - 0xff -- plane 1
    "11111111", -- 3593 - 0xe09  :  255 - 0xff
    "11111111", -- 3594 - 0xe0a  :  255 - 0xff
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "11111111", -- 3596 - 0xe0c  :  255 - 0xff
    "11111111", -- 3597 - 0xe0d  :  255 - 0xff
    "11111111", -- 3598 - 0xe0e  :  255 - 0xff
    "11111111", -- 3599 - 0xe0f  :  255 - 0xff
    "11111111", -- 3600 - 0xe10  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "11111111", -- 3602 - 0xe12  :  255 - 0xff
    "11111111", -- 3603 - 0xe13  :  255 - 0xff
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111111", -- 3605 - 0xe15  :  255 - 0xff
    "11111111", -- 3606 - 0xe16  :  255 - 0xff
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "11111111", -- 3608 - 0xe18  :  255 - 0xff -- plane 1
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "11111111", -- 3610 - 0xe1a  :  255 - 0xff
    "11111111", -- 3611 - 0xe1b  :  255 - 0xff
    "11111111", -- 3612 - 0xe1c  :  255 - 0xff
    "11111111", -- 3613 - 0xe1d  :  255 - 0xff
    "11111111", -- 3614 - 0xe1e  :  255 - 0xff
    "11111111", -- 3615 - 0xe1f  :  255 - 0xff
    "11111111", -- 3616 - 0xe20  :  255 - 0xff -- Sprite 0xe2
    "11111111", -- 3617 - 0xe21  :  255 - 0xff
    "11111111", -- 3618 - 0xe22  :  255 - 0xff
    "11111111", -- 3619 - 0xe23  :  255 - 0xff
    "11111111", -- 3620 - 0xe24  :  255 - 0xff
    "11111111", -- 3621 - 0xe25  :  255 - 0xff
    "11111111", -- 3622 - 0xe26  :  255 - 0xff
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111111", -- 3624 - 0xe28  :  255 - 0xff -- plane 1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "11111111", -- 3631 - 0xe2f  :  255 - 0xff
    "11111111", -- 3632 - 0xe30  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 3633 - 0xe31  :  255 - 0xff
    "11111111", -- 3634 - 0xe32  :  255 - 0xff
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "11111111", -- 3636 - 0xe34  :  255 - 0xff
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "11111111", -- 3640 - 0xe38  :  255 - 0xff -- plane 1
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "11111111", -- 3642 - 0xe3a  :  255 - 0xff
    "11111111", -- 3643 - 0xe3b  :  255 - 0xff
    "11111111", -- 3644 - 0xe3c  :  255 - 0xff
    "11111111", -- 3645 - 0xe3d  :  255 - 0xff
    "11111111", -- 3646 - 0xe3e  :  255 - 0xff
    "11111111", -- 3647 - 0xe3f  :  255 - 0xff
    "11111111", -- 3648 - 0xe40  :  255 - 0xff -- Sprite 0xe4
    "11111111", -- 3649 - 0xe41  :  255 - 0xff
    "11111111", -- 3650 - 0xe42  :  255 - 0xff
    "11111111", -- 3651 - 0xe43  :  255 - 0xff
    "11111111", -- 3652 - 0xe44  :  255 - 0xff
    "11111111", -- 3653 - 0xe45  :  255 - 0xff
    "11111111", -- 3654 - 0xe46  :  255 - 0xff
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11111111", -- 3656 - 0xe48  :  255 - 0xff -- plane 1
    "11111111", -- 3657 - 0xe49  :  255 - 0xff
    "11111111", -- 3658 - 0xe4a  :  255 - 0xff
    "11111111", -- 3659 - 0xe4b  :  255 - 0xff
    "11111111", -- 3660 - 0xe4c  :  255 - 0xff
    "11111111", -- 3661 - 0xe4d  :  255 - 0xff
    "11111111", -- 3662 - 0xe4e  :  255 - 0xff
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "11111111", -- 3664 - 0xe50  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 3665 - 0xe51  :  255 - 0xff
    "11111111", -- 3666 - 0xe52  :  255 - 0xff
    "11111111", -- 3667 - 0xe53  :  255 - 0xff
    "11111111", -- 3668 - 0xe54  :  255 - 0xff
    "11111111", -- 3669 - 0xe55  :  255 - 0xff
    "11111111", -- 3670 - 0xe56  :  255 - 0xff
    "11111111", -- 3671 - 0xe57  :  255 - 0xff
    "11111111", -- 3672 - 0xe58  :  255 - 0xff -- plane 1
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "11111111", -- 3674 - 0xe5a  :  255 - 0xff
    "11111111", -- 3675 - 0xe5b  :  255 - 0xff
    "11111111", -- 3676 - 0xe5c  :  255 - 0xff
    "11111111", -- 3677 - 0xe5d  :  255 - 0xff
    "11111111", -- 3678 - 0xe5e  :  255 - 0xff
    "11111111", -- 3679 - 0xe5f  :  255 - 0xff
    "11111111", -- 3680 - 0xe60  :  255 - 0xff -- Sprite 0xe6
    "11111111", -- 3681 - 0xe61  :  255 - 0xff
    "11111111", -- 3682 - 0xe62  :  255 - 0xff
    "11111111", -- 3683 - 0xe63  :  255 - 0xff
    "11111111", -- 3684 - 0xe64  :  255 - 0xff
    "11111111", -- 3685 - 0xe65  :  255 - 0xff
    "11111111", -- 3686 - 0xe66  :  255 - 0xff
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "11111111", -- 3688 - 0xe68  :  255 - 0xff -- plane 1
    "11111111", -- 3689 - 0xe69  :  255 - 0xff
    "11111111", -- 3690 - 0xe6a  :  255 - 0xff
    "11111111", -- 3691 - 0xe6b  :  255 - 0xff
    "11111111", -- 3692 - 0xe6c  :  255 - 0xff
    "11111111", -- 3693 - 0xe6d  :  255 - 0xff
    "11111111", -- 3694 - 0xe6e  :  255 - 0xff
    "11111111", -- 3695 - 0xe6f  :  255 - 0xff
    "11111111", -- 3696 - 0xe70  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 3697 - 0xe71  :  255 - 0xff
    "11111111", -- 3698 - 0xe72  :  255 - 0xff
    "11111111", -- 3699 - 0xe73  :  255 - 0xff
    "11111111", -- 3700 - 0xe74  :  255 - 0xff
    "11111111", -- 3701 - 0xe75  :  255 - 0xff
    "11111111", -- 3702 - 0xe76  :  255 - 0xff
    "11111111", -- 3703 - 0xe77  :  255 - 0xff
    "11111111", -- 3704 - 0xe78  :  255 - 0xff -- plane 1
    "11111111", -- 3705 - 0xe79  :  255 - 0xff
    "11111111", -- 3706 - 0xe7a  :  255 - 0xff
    "11111111", -- 3707 - 0xe7b  :  255 - 0xff
    "11111111", -- 3708 - 0xe7c  :  255 - 0xff
    "11111111", -- 3709 - 0xe7d  :  255 - 0xff
    "11111111", -- 3710 - 0xe7e  :  255 - 0xff
    "11111111", -- 3711 - 0xe7f  :  255 - 0xff
    "11111111", -- 3712 - 0xe80  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "11111111", -- 3715 - 0xe83  :  255 - 0xff
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11111111", -- 3720 - 0xe88  :  255 - 0xff -- plane 1
    "11111111", -- 3721 - 0xe89  :  255 - 0xff
    "11111111", -- 3722 - 0xe8a  :  255 - 0xff
    "11111111", -- 3723 - 0xe8b  :  255 - 0xff
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11111111", -- 3728 - 0xe90  :  255 - 0xff -- Sprite 0xe9
    "11111111", -- 3729 - 0xe91  :  255 - 0xff
    "11111111", -- 3730 - 0xe92  :  255 - 0xff
    "11111111", -- 3731 - 0xe93  :  255 - 0xff
    "11111111", -- 3732 - 0xe94  :  255 - 0xff
    "11111111", -- 3733 - 0xe95  :  255 - 0xff
    "11111111", -- 3734 - 0xe96  :  255 - 0xff
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111111", -- 3736 - 0xe98  :  255 - 0xff -- plane 1
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111111", -- 3740 - 0xe9c  :  255 - 0xff
    "11111111", -- 3741 - 0xe9d  :  255 - 0xff
    "11111111", -- 3742 - 0xe9e  :  255 - 0xff
    "11111111", -- 3743 - 0xe9f  :  255 - 0xff
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "11111111", -- 3748 - 0xea4  :  255 - 0xff
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "11111111", -- 3751 - 0xea7  :  255 - 0xff
    "11111111", -- 3752 - 0xea8  :  255 - 0xff -- plane 1
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "11111111", -- 3760 - 0xeb0  :  255 - 0xff -- Sprite 0xeb
    "11111111", -- 3761 - 0xeb1  :  255 - 0xff
    "11111111", -- 3762 - 0xeb2  :  255 - 0xff
    "11111111", -- 3763 - 0xeb3  :  255 - 0xff
    "11111111", -- 3764 - 0xeb4  :  255 - 0xff
    "11111111", -- 3765 - 0xeb5  :  255 - 0xff
    "11111111", -- 3766 - 0xeb6  :  255 - 0xff
    "11111111", -- 3767 - 0xeb7  :  255 - 0xff
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff -- plane 1
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "11111111", -- 3772 - 0xebc  :  255 - 0xff
    "11111111", -- 3773 - 0xebd  :  255 - 0xff
    "11111111", -- 3774 - 0xebe  :  255 - 0xff
    "11111111", -- 3775 - 0xebf  :  255 - 0xff
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "00000001", -- 3777 - 0xec1  :    1 - 0x1
    "00000011", -- 3778 - 0xec2  :    3 - 0x3
    "00110011", -- 3779 - 0xec3  :   51 - 0x33
    "00011001", -- 3780 - 0xec4  :   25 - 0x19
    "00001111", -- 3781 - 0xec5  :   15 - 0xf
    "00111111", -- 3782 - 0xec6  :   63 - 0x3f
    "00011111", -- 3783 - 0xec7  :   31 - 0x1f
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "00000001", -- 3785 - 0xec9  :    1 - 0x1
    "00000011", -- 3786 - 0xeca  :    3 - 0x3
    "00110011", -- 3787 - 0xecb  :   51 - 0x33
    "00011001", -- 3788 - 0xecc  :   25 - 0x19
    "00001111", -- 3789 - 0xecd  :   15 - 0xf
    "00111111", -- 3790 - 0xece  :   63 - 0x3f
    "00011111", -- 3791 - 0xecf  :   31 - 0x1f
    "00101011", -- 3792 - 0xed0  :   43 - 0x2b -- Sprite 0xed
    "00000111", -- 3793 - 0xed1  :    7 - 0x7
    "00000101", -- 3794 - 0xed2  :    5 - 0x5
    "00001101", -- 3795 - 0xed3  :   13 - 0xd
    "00001011", -- 3796 - 0xed4  :   11 - 0xb
    "00011011", -- 3797 - 0xed5  :   27 - 0x1b
    "00011011", -- 3798 - 0xed6  :   27 - 0x1b
    "00111011", -- 3799 - 0xed7  :   59 - 0x3b
    "00101011", -- 3800 - 0xed8  :   43 - 0x2b -- plane 1
    "00000111", -- 3801 - 0xed9  :    7 - 0x7
    "00000101", -- 3802 - 0xeda  :    5 - 0x5
    "00001101", -- 3803 - 0xedb  :   13 - 0xd
    "00001011", -- 3804 - 0xedc  :   11 - 0xb
    "00011011", -- 3805 - 0xedd  :   27 - 0x1b
    "00011011", -- 3806 - 0xede  :   27 - 0x1b
    "00000011", -- 3807 - 0xedf  :    3 - 0x3
    "00001001", -- 3808 - 0xee0  :    9 - 0x9 -- Sprite 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000111", -- 3810 - 0xee2  :    7 - 0x7
    "00000111", -- 3811 - 0xee3  :    7 - 0x7
    "00001111", -- 3812 - 0xee4  :   15 - 0xf
    "00001101", -- 3813 - 0xee5  :   13 - 0xd
    "00000001", -- 3814 - 0xee6  :    1 - 0x1
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000001", -- 3816 - 0xee8  :    1 - 0x1 -- plane 1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000011", -- 3818 - 0xeea  :    3 - 0x3
    "00000101", -- 3819 - 0xeeb  :    5 - 0x5
    "00001110", -- 3820 - 0xeec  :   14 - 0xe
    "00001101", -- 3821 - 0xeed  :   13 - 0xd
    "00000001", -- 3822 - 0xeee  :    1 - 0x1
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "11111000", -- 3824 - 0xef0  :  248 - 0xf8 -- Sprite 0xef
    "11111100", -- 3825 - 0xef1  :  252 - 0xfc
    "11111000", -- 3826 - 0xef2  :  248 - 0xf8
    "11101100", -- 3827 - 0xef3  :  236 - 0xec
    "11111000", -- 3828 - 0xef4  :  248 - 0xf8
    "11110000", -- 3829 - 0xef5  :  240 - 0xf0
    "11000000", -- 3830 - 0xef6  :  192 - 0xc0
    "11000000", -- 3831 - 0xef7  :  192 - 0xc0
    "11111000", -- 3832 - 0xef8  :  248 - 0xf8 -- plane 1
    "11111100", -- 3833 - 0xef9  :  252 - 0xfc
    "11000000", -- 3834 - 0xefa  :  192 - 0xc0
    "01000000", -- 3835 - 0xefb  :   64 - 0x40
    "10000000", -- 3836 - 0xefc  :  128 - 0x80
    "10000000", -- 3837 - 0xefd  :  128 - 0x80
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "10000000", -- 3839 - 0xeff  :  128 - 0x80
    "11110000", -- 3840 - 0xf00  :  240 - 0xf0 -- Sprite 0xf0
    "11111000", -- 3841 - 0xf01  :  248 - 0xf8
    "11111000", -- 3842 - 0xf02  :  248 - 0xf8
    "11101000", -- 3843 - 0xf03  :  232 - 0xe8
    "11001100", -- 3844 - 0xf04  :  204 - 0xcc
    "11100110", -- 3845 - 0xf05  :  230 - 0xe6
    "11111011", -- 3846 - 0xf06  :  251 - 0xfb
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11010000", -- 3848 - 0xf08  :  208 - 0xd0 -- plane 1
    "11111000", -- 3849 - 0xf09  :  248 - 0xf8
    "11111000", -- 3850 - 0xf0a  :  248 - 0xf8
    "11101000", -- 3851 - 0xf0b  :  232 - 0xe8
    "11001100", -- 3852 - 0xf0c  :  204 - 0xcc
    "11100110", -- 3853 - 0xf0d  :  230 - 0xe6
    "11111000", -- 3854 - 0xf0e  :  248 - 0xf8
    "11111110", -- 3855 - 0xf0f  :  254 - 0xfe
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Sprite 0xf1
    "11111110", -- 3857 - 0xf11  :  254 - 0xfe
    "11111110", -- 3858 - 0xf12  :  254 - 0xfe
    "11111110", -- 3859 - 0xf13  :  254 - 0xfe
    "11111110", -- 3860 - 0xf14  :  254 - 0xfe
    "10001111", -- 3861 - 0xf15  :  143 - 0x8f
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "11111110", -- 3864 - 0xf18  :  254 - 0xfe -- plane 1
    "11111110", -- 3865 - 0xf19  :  254 - 0xfe
    "00000110", -- 3866 - 0xf1a  :    6 - 0x6
    "11111000", -- 3867 - 0xf1b  :  248 - 0xf8
    "00001110", -- 3868 - 0xf1c  :   14 - 0xe
    "10000000", -- 3869 - 0xf1d  :  128 - 0x80
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000001", -- 3872 - 0xf20  :    1 - 0x1 -- Sprite 0xf2
    "00001111", -- 3873 - 0xf21  :   15 - 0xf
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000100", -- 3876 - 0xf24  :    4 - 0x4
    "00011110", -- 3877 - 0xf25  :   30 - 0x1e
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000011", -- 3879 - 0xf27  :    3 - 0x3
    "00000001", -- 3880 - 0xf28  :    1 - 0x1 -- plane 1
    "00001111", -- 3881 - 0xf29  :   15 - 0xf
    "00000111", -- 3882 - 0xf2a  :    7 - 0x7
    "00011101", -- 3883 - 0xf2b  :   29 - 0x1d
    "00111011", -- 3884 - 0xf2c  :   59 - 0x3b
    "00000001", -- 3885 - 0xf2d  :    1 - 0x1
    "00001111", -- 3886 - 0xf2e  :   15 - 0xf
    "00000010", -- 3887 - 0xf2f  :    2 - 0x2
    "00000111", -- 3888 - 0xf30  :    7 - 0x7 -- Sprite 0xf3
    "00001111", -- 3889 - 0xf31  :   15 - 0xf
    "00011111", -- 3890 - 0xf32  :   31 - 0x1f
    "00001111", -- 3891 - 0xf33  :   15 - 0xf
    "00000111", -- 3892 - 0xf34  :    7 - 0x7
    "00001111", -- 3893 - 0xf35  :   15 - 0xf
    "00001111", -- 3894 - 0xf36  :   15 - 0xf
    "00000011", -- 3895 - 0xf37  :    3 - 0x3
    "00000010", -- 3896 - 0xf38  :    2 - 0x2 -- plane 1
    "00000011", -- 3897 - 0xf39  :    3 - 0x3
    "00000010", -- 3898 - 0xf3a  :    2 - 0x2
    "01110111", -- 3899 - 0xf3b  :  119 - 0x77
    "00010111", -- 3900 - 0xf3c  :   23 - 0x17
    "00000001", -- 3901 - 0xf3d  :    1 - 0x1
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "11100000", -- 3904 - 0xf40  :  224 - 0xe0 -- Sprite 0xf4
    "11110000", -- 3905 - 0xf41  :  240 - 0xf0
    "11110000", -- 3906 - 0xf42  :  240 - 0xf0
    "01001000", -- 3907 - 0xf43  :   72 - 0x48
    "11001000", -- 3908 - 0xf44  :  200 - 0xc8
    "10011100", -- 3909 - 0xf45  :  156 - 0x9c
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "11110000", -- 3911 - 0xf47  :  240 - 0xf0
    "11100000", -- 3912 - 0xf48  :  224 - 0xe0 -- plane 1
    "11110000", -- 3913 - 0xf49  :  240 - 0xf0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "10110000", -- 3915 - 0xf4b  :  176 - 0xb0
    "00110000", -- 3916 - 0xf4c  :   48 - 0x30
    "01100000", -- 3917 - 0xf4d  :   96 - 0x60
    "11110000", -- 3918 - 0xf4e  :  240 - 0xf0
    "00010000", -- 3919 - 0xf4f  :   16 - 0x10
    "11111000", -- 3920 - 0xf50  :  248 - 0xf8 -- Sprite 0xf5
    "11111100", -- 3921 - 0xf51  :  252 - 0xfc
    "11111100", -- 3922 - 0xf52  :  252 - 0xfc
    "11111000", -- 3923 - 0xf53  :  248 - 0xf8
    "11111000", -- 3924 - 0xf54  :  248 - 0xf8
    "01111000", -- 3925 - 0xf55  :  120 - 0x78
    "01110000", -- 3926 - 0xf56  :  112 - 0x70
    "01100000", -- 3927 - 0xf57  :   96 - 0x60
    "00110000", -- 3928 - 0xf58  :   48 - 0x30 -- plane 1
    "11110000", -- 3929 - 0xf59  :  240 - 0xf0
    "11010000", -- 3930 - 0xf5a  :  208 - 0xd0
    "11111100", -- 3931 - 0xf5b  :  252 - 0xfc
    "11111110", -- 3932 - 0xf5c  :  254 - 0xfe
    "00001000", -- 3933 - 0xf5d  :    8 - 0x8
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "01111100", -- 3938 - 0xf62  :  124 - 0x7c
    "10001010", -- 3939 - 0xf63  :  138 - 0x8a
    "11111110", -- 3940 - 0xf64  :  254 - 0xfe
    "11111110", -- 3941 - 0xf65  :  254 - 0xfe
    "11111110", -- 3942 - 0xf66  :  254 - 0xfe
    "11111110", -- 3943 - 0xf67  :  254 - 0xfe
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- plane 1
    "00010000", -- 3945 - 0xf69  :   16 - 0x10
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "01110100", -- 3947 - 0xf6b  :  116 - 0x74
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "11111110", -- 3952 - 0xf70  :  254 - 0xfe -- Sprite 0xf7
    "01111100", -- 3953 - 0xf71  :  124 - 0x7c
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0 -- plane 1
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00010000", -- 3962 - 0xf7a  :   16 - 0x10
    "00010000", -- 3963 - 0xf7b  :   16 - 0x10
    "00010000", -- 3964 - 0xf7c  :   16 - 0x10
    "00010000", -- 3965 - 0xf7d  :   16 - 0x10
    "00010000", -- 3966 - 0xf7e  :   16 - 0x10
    "00010000", -- 3967 - 0xf7f  :   16 - 0x10
    "00000111", -- 3968 - 0xf80  :    7 - 0x7 -- Sprite 0xf8
    "00001011", -- 3969 - 0xf81  :   11 - 0xb
    "00001111", -- 3970 - 0xf82  :   15 - 0xf
    "00001011", -- 3971 - 0xf83  :   11 - 0xb
    "00001011", -- 3972 - 0xf84  :   11 - 0xb
    "00001011", -- 3973 - 0xf85  :   11 - 0xb
    "00001011", -- 3974 - 0xf86  :   11 - 0xb
    "00000111", -- 3975 - 0xf87  :    7 - 0x7
    "00000000", -- 3976 - 0xf88  :    0 - 0x0 -- plane 1
    "00000100", -- 3977 - 0xf89  :    4 - 0x4
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00010100", -- 3979 - 0xf8b  :   20 - 0x14
    "00000100", -- 3980 - 0xf8c  :    4 - 0x4
    "00000100", -- 3981 - 0xf8d  :    4 - 0x4
    "00000100", -- 3982 - 0xf8e  :    4 - 0x4
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "11000000", -- 3984 - 0xf90  :  192 - 0xc0 -- Sprite 0xf9
    "11100000", -- 3985 - 0xf91  :  224 - 0xe0
    "11100000", -- 3986 - 0xf92  :  224 - 0xe0
    "11100000", -- 3987 - 0xf93  :  224 - 0xe0
    "11100000", -- 3988 - 0xf94  :  224 - 0xe0
    "11100000", -- 3989 - 0xf95  :  224 - 0xe0
    "11100000", -- 3990 - 0xf96  :  224 - 0xe0
    "11000000", -- 3991 - 0xf97  :  192 - 0xc0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- plane 1
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00011111", -- 3995 - 0xf9b  :   31 - 0x1f
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000011", -- 4000 - 0xfa0  :    3 - 0x3 -- Sprite 0xfa
    "00000111", -- 4001 - 0xfa1  :    7 - 0x7
    "00000111", -- 4002 - 0xfa2  :    7 - 0x7
    "00000111", -- 4003 - 0xfa3  :    7 - 0x7
    "00000111", -- 4004 - 0xfa4  :    7 - 0x7
    "00000111", -- 4005 - 0xfa5  :    7 - 0x7
    "00000111", -- 4006 - 0xfa6  :    7 - 0x7
    "00000011", -- 4007 - 0xfa7  :    3 - 0x3
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- plane 1
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "11111000", -- 4011 - 0xfab  :  248 - 0xf8
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "11100000", -- 4016 - 0xfb0  :  224 - 0xe0 -- Sprite 0xfb
    "11010000", -- 4017 - 0xfb1  :  208 - 0xd0
    "11010000", -- 4018 - 0xfb2  :  208 - 0xd0
    "11010000", -- 4019 - 0xfb3  :  208 - 0xd0
    "11010000", -- 4020 - 0xfb4  :  208 - 0xd0
    "11110000", -- 4021 - 0xfb5  :  240 - 0xf0
    "11010000", -- 4022 - 0xfb6  :  208 - 0xd0
    "11100000", -- 4023 - 0xfb7  :  224 - 0xe0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- plane 1
    "00100000", -- 4025 - 0xfb9  :   32 - 0x20
    "00100000", -- 4026 - 0xfba  :   32 - 0x20
    "00101000", -- 4027 - 0xfbb  :   40 - 0x28
    "00100000", -- 4028 - 0xfbc  :   32 - 0x20
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00100000", -- 4030 - 0xfbe  :   32 - 0x20
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Sprite 0xfc
    "00000001", -- 4033 - 0xfc1  :    1 - 0x1
    "00010011", -- 4034 - 0xfc2  :   19 - 0x13
    "00110111", -- 4035 - 0xfc3  :   55 - 0x37
    "00111011", -- 4036 - 0xfc4  :   59 - 0x3b
    "01110100", -- 4037 - 0xfc5  :  116 - 0x74
    "01111010", -- 4038 - 0xfc6  :  122 - 0x7a
    "00111110", -- 4039 - 0xfc7  :   62 - 0x3e
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0 -- plane 1
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00001000", -- 4042 - 0xfca  :    8 - 0x8
    "00100101", -- 4043 - 0xfcb  :   37 - 0x25
    "00010010", -- 4044 - 0xfcc  :   18 - 0x12
    "01010011", -- 4045 - 0xfcd  :   83 - 0x53
    "00110011", -- 4046 - 0xfce  :   51 - 0x33
    "00111001", -- 4047 - 0xfcf  :   57 - 0x39
    "11011000", -- 4048 - 0xfd0  :  216 - 0xd8 -- Sprite 0xfd
    "10011000", -- 4049 - 0xfd1  :  152 - 0x98
    "10101000", -- 4050 - 0xfd2  :  168 - 0xa8
    "11011000", -- 4051 - 0xfd3  :  216 - 0xd8
    "11011010", -- 4052 - 0xfd4  :  218 - 0xda
    "01110100", -- 4053 - 0xfd5  :  116 - 0x74
    "00101000", -- 4054 - 0xfd6  :   40 - 0x28
    "11001000", -- 4055 - 0xfd7  :  200 - 0xc8
    "00001000", -- 4056 - 0xfd8  :    8 - 0x8 -- plane 1
    "10000000", -- 4057 - 0xfd9  :  128 - 0x80
    "00110000", -- 4058 - 0xfda  :   48 - 0x30
    "10011100", -- 4059 - 0xfdb  :  156 - 0x9c
    "11001010", -- 4060 - 0xfdc  :  202 - 0xca
    "10111000", -- 4061 - 0xfdd  :  184 - 0xb8
    "10011000", -- 4062 - 0xfde  :  152 - 0x98
    "01111000", -- 4063 - 0xfdf  :  120 - 0x78
    "00001000", -- 4064 - 0xfe0  :    8 - 0x8 -- Sprite 0xfe
    "01011001", -- 4065 - 0xfe1  :   89 - 0x59
    "00110000", -- 4066 - 0xfe2  :   48 - 0x30
    "01110001", -- 4067 - 0xfe3  :  113 - 0x71
    "01111001", -- 4068 - 0xfe4  :  121 - 0x79
    "00101011", -- 4069 - 0xfe5  :   43 - 0x2b
    "00110110", -- 4070 - 0xfe6  :   54 - 0x36
    "00010110", -- 4071 - 0xfe7  :   22 - 0x16
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- plane 1
    "00001000", -- 4073 - 0xfe9  :    8 - 0x8
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "01000000", -- 4075 - 0xfeb  :   64 - 0x40
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00110001", -- 4077 - 0xfed  :   49 - 0x31
    "00111101", -- 4078 - 0xfee  :   61 - 0x3d
    "00011001", -- 4079 - 0xfef  :   25 - 0x19
    "11000110", -- 4080 - 0xff0  :  198 - 0xc6 -- Sprite 0xff
    "11000100", -- 4081 - 0xff1  :  196 - 0xc4
    "11001100", -- 4082 - 0xff2  :  204 - 0xcc
    "11001100", -- 4083 - 0xff3  :  204 - 0xcc
    "10111000", -- 4084 - 0xff4  :  184 - 0xb8
    "01111100", -- 4085 - 0xff5  :  124 - 0x7c
    "11101100", -- 4086 - 0xff6  :  236 - 0xec
    "11001000", -- 4087 - 0xff7  :  200 - 0xc8
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- plane 1
    "10000000", -- 4089 - 0xff9  :  128 - 0x80
    "11000000", -- 4090 - 0xffa  :  192 - 0xc0
    "11000000", -- 4091 - 0xffb  :  192 - 0xc0
    "11000000", -- 4092 - 0xffc  :  192 - 0xc0
    "10001000", -- 4093 - 0xffd  :  136 - 0x88
    "10111000", -- 4094 - 0xffe  :  184 - 0xb8
    "10111000"  -- 4095 - 0xfff  :  184 - 0xb8
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
