--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_menuscr.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE0_SPRILO_MENU is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE0_SPRILO_MENU;

architecture BEHAVIORAL of ROM_NTABLE0_SPRILO_MENU is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11111010", --    3 -  0x3  :  250 - 0xfa
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11111010", --   14 -  0xe  :  250 - 0xfa
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11111010", --   33 - 0x21  :  250 - 0xfa
    "11111010", --   34 - 0x22  :  250 - 0xfa
    "11111010", --   35 - 0x23  :  250 - 0xfa
    "11111010", --   36 - 0x24  :  250 - 0xfa
    "11111010", --   37 - 0x25  :  250 - 0xfa
    "11111010", --   38 - 0x26  :  250 - 0xfa
    "11111001", --   39 - 0x27  :  249 - 0xf9
    "11111010", --   40 - 0x28  :  250 - 0xfa
    "11111010", --   41 - 0x29  :  250 - 0xfa
    "11111010", --   42 - 0x2a  :  250 - 0xfa
    "11111010", --   43 - 0x2b  :  250 - 0xfa
    "11111010", --   44 - 0x2c  :  250 - 0xfa
    "11111010", --   45 - 0x2d  :  250 - 0xfa
    "11111010", --   46 - 0x2e  :  250 - 0xfa
    "11111010", --   47 - 0x2f  :  250 - 0xfa
    "11111010", --   48 - 0x30  :  250 - 0xfa
    "11111001", --   49 - 0x31  :  249 - 0xf9
    "11111010", --   50 - 0x32  :  250 - 0xfa
    "11111010", --   51 - 0x33  :  250 - 0xfa
    "11111010", --   52 - 0x34  :  250 - 0xfa
    "11111010", --   53 - 0x35  :  250 - 0xfa
    "11111010", --   54 - 0x36  :  250 - 0xfa
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11111010", --   57 - 0x39  :  250 - 0xfa
    "11111010", --   58 - 0x3a  :  250 - 0xfa
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111001", --   60 - 0x3c  :  249 - 0xf9
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11111010", --   64 - 0x40  :  250 - 0xfa -- line 0x2
    "11111010", --   65 - 0x41  :  250 - 0xfa
    "11111010", --   66 - 0x42  :  250 - 0xfa
    "11111010", --   67 - 0x43  :  250 - 0xfa
    "11111010", --   68 - 0x44  :  250 - 0xfa
    "11111010", --   69 - 0x45  :  250 - 0xfa
    "11111010", --   70 - 0x46  :  250 - 0xfa
    "11111010", --   71 - 0x47  :  250 - 0xfa
    "11111010", --   72 - 0x48  :  250 - 0xfa
    "11111010", --   73 - 0x49  :  250 - 0xfa
    "11111001", --   74 - 0x4a  :  249 - 0xf9
    "11111010", --   75 - 0x4b  :  250 - 0xfa
    "11111010", --   76 - 0x4c  :  250 - 0xfa
    "11111010", --   77 - 0x4d  :  250 - 0xfa
    "11101010", --   78 - 0x4e  :  234 - 0xea
    "11111010", --   79 - 0x4f  :  250 - 0xfa
    "11111010", --   80 - 0x50  :  250 - 0xfa
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111010", --   83 - 0x53  :  250 - 0xfa
    "11111010", --   84 - 0x54  :  250 - 0xfa
    "11111010", --   85 - 0x55  :  250 - 0xfa
    "11111010", --   86 - 0x56  :  250 - 0xfa
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11111010", --   97 - 0x61  :  250 - 0xfa
    "11111010", --   98 - 0x62  :  250 - 0xfa
    "11111010", --   99 - 0x63  :  250 - 0xfa
    "11111010", --  100 - 0x64  :  250 - 0xfa
    "11111010", --  101 - 0x65  :  250 - 0xfa
    "11111010", --  102 - 0x66  :  250 - 0xfa
    "11111010", --  103 - 0x67  :  250 - 0xfa
    "11111010", --  104 - 0x68  :  250 - 0xfa
    "11111010", --  105 - 0x69  :  250 - 0xfa
    "11111010", --  106 - 0x6a  :  250 - 0xfa
    "11111010", --  107 - 0x6b  :  250 - 0xfa
    "11111010", --  108 - 0x6c  :  250 - 0xfa
    "11111010", --  109 - 0x6d  :  250 - 0xfa
    "11111010", --  110 - 0x6e  :  250 - 0xfa
    "11111010", --  111 - 0x6f  :  250 - 0xfa
    "11111010", --  112 - 0x70  :  250 - 0xfa
    "11111010", --  113 - 0x71  :  250 - 0xfa
    "11111010", --  114 - 0x72  :  250 - 0xfa
    "11111010", --  115 - 0x73  :  250 - 0xfa
    "11111010", --  116 - 0x74  :  250 - 0xfa
    "11111010", --  117 - 0x75  :  250 - 0xfa
    "11111010", --  118 - 0x76  :  250 - 0xfa
    "11111010", --  119 - 0x77  :  250 - 0xfa
    "11111010", --  120 - 0x78  :  250 - 0xfa
    "11101010", --  121 - 0x79  :  234 - 0xea
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11101010", --  125 - 0x7d  :  234 - 0xea
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11111010", --  128 - 0x80  :  250 - 0xfa -- line 0x4
    "11111010", --  129 - 0x81  :  250 - 0xfa
    "11111010", --  130 - 0x82  :  250 - 0xfa
    "11111010", --  131 - 0x83  :  250 - 0xfa
    "11101010", --  132 - 0x84  :  234 - 0xea
    "11111010", --  133 - 0x85  :  250 - 0xfa
    "11111010", --  134 - 0x86  :  250 - 0xfa
    "11111001", --  135 - 0x87  :  249 - 0xf9
    "11111010", --  136 - 0x88  :  250 - 0xfa
    "11111010", --  137 - 0x89  :  250 - 0xfa
    "11111010", --  138 - 0x8a  :  250 - 0xfa
    "11111010", --  139 - 0x8b  :  250 - 0xfa
    "11111010", --  140 - 0x8c  :  250 - 0xfa
    "11111010", --  141 - 0x8d  :  250 - 0xfa
    "11111010", --  142 - 0x8e  :  250 - 0xfa
    "11111010", --  143 - 0x8f  :  250 - 0xfa
    "11111010", --  144 - 0x90  :  250 - 0xfa
    "11111010", --  145 - 0x91  :  250 - 0xfa
    "11111010", --  146 - 0x92  :  250 - 0xfa
    "11111010", --  147 - 0x93  :  250 - 0xfa
    "11111010", --  148 - 0x94  :  250 - 0xfa
    "11111001", --  149 - 0x95  :  249 - 0xf9
    "11111010", --  150 - 0x96  :  250 - 0xfa
    "11111010", --  151 - 0x97  :  250 - 0xfa
    "11111010", --  152 - 0x98  :  250 - 0xfa
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11111010", --  154 - 0x9a  :  250 - 0xfa
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111010", --  156 - 0x9c  :  250 - 0xfa
    "11111010", --  157 - 0x9d  :  250 - 0xfa
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111010", --  161 - 0xa1  :  250 - 0xfa
    "11111010", --  162 - 0xa2  :  250 - 0xfa
    "11111010", --  163 - 0xa3  :  250 - 0xfa
    "11111010", --  164 - 0xa4  :  250 - 0xfa
    "11111010", --  165 - 0xa5  :  250 - 0xfa
    "11111010", --  166 - 0xa6  :  250 - 0xfa
    "11111010", --  167 - 0xa7  :  250 - 0xfa
    "11111010", --  168 - 0xa8  :  250 - 0xfa
    "11111010", --  169 - 0xa9  :  250 - 0xfa
    "11111010", --  170 - 0xaa  :  250 - 0xfa
    "11001101", --  171 - 0xab  :  205 - 0xcd
    "11101101", --  172 - 0xac  :  237 - 0xed
    "11101101", --  173 - 0xad  :  237 - 0xed
    "11101101", --  174 - 0xae  :  237 - 0xed
    "11101101", --  175 - 0xaf  :  237 - 0xed
    "11101101", --  176 - 0xb0  :  237 - 0xed
    "11101101", --  177 - 0xb1  :  237 - 0xed
    "11101101", --  178 - 0xb2  :  237 - 0xed
    "11101101", --  179 - 0xb3  :  237 - 0xed
    "11001110", --  180 - 0xb4  :  206 - 0xce
    "11111010", --  181 - 0xb5  :  250 - 0xfa
    "11111010", --  182 - 0xb6  :  250 - 0xfa
    "11111010", --  183 - 0xb7  :  250 - 0xfa
    "11111010", --  184 - 0xb8  :  250 - 0xfa
    "11111010", --  185 - 0xb9  :  250 - 0xfa
    "11111010", --  186 - 0xba  :  250 - 0xfa
    "11111010", --  187 - 0xbb  :  250 - 0xfa
    "11111010", --  188 - 0xbc  :  250 - 0xfa
    "11111010", --  189 - 0xbd  :  250 - 0xfa
    "11111010", --  190 - 0xbe  :  250 - 0xfa
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111001", --  192 - 0xc0  :  249 - 0xf9 -- line 0x6
    "11111010", --  193 - 0xc1  :  250 - 0xfa
    "11111010", --  194 - 0xc2  :  250 - 0xfa
    "11111010", --  195 - 0xc3  :  250 - 0xfa
    "11111010", --  196 - 0xc4  :  250 - 0xfa
    "11111010", --  197 - 0xc5  :  250 - 0xfa
    "11111010", --  198 - 0xc6  :  250 - 0xfa
    "11111010", --  199 - 0xc7  :  250 - 0xfa
    "11111010", --  200 - 0xc8  :  250 - 0xfa
    "11111010", --  201 - 0xc9  :  250 - 0xfa
    "11111010", --  202 - 0xca  :  250 - 0xfa
    "11101110", --  203 - 0xcb  :  238 - 0xee
    "11111010", --  204 - 0xcc  :  250 - 0xfa
    "11111010", --  205 - 0xcd  :  250 - 0xfa
    "11111010", --  206 - 0xce  :  250 - 0xfa
    "11111010", --  207 - 0xcf  :  250 - 0xfa
    "11111010", --  208 - 0xd0  :  250 - 0xfa
    "11111010", --  209 - 0xd1  :  250 - 0xfa
    "11111010", --  210 - 0xd2  :  250 - 0xfa
    "11111010", --  211 - 0xd3  :  250 - 0xfa
    "11101110", --  212 - 0xd4  :  238 - 0xee
    "11111010", --  213 - 0xd5  :  250 - 0xfa
    "11111010", --  214 - 0xd6  :  250 - 0xfa
    "11111010", --  215 - 0xd7  :  250 - 0xfa
    "11111010", --  216 - 0xd8  :  250 - 0xfa
    "11111010", --  217 - 0xd9  :  250 - 0xfa
    "11111010", --  218 - 0xda  :  250 - 0xfa
    "11111001", --  219 - 0xdb  :  249 - 0xf9
    "11111010", --  220 - 0xdc  :  250 - 0xfa
    "11111010", --  221 - 0xdd  :  250 - 0xfa
    "11111010", --  222 - 0xde  :  250 - 0xfa
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111010", --  225 - 0xe1  :  250 - 0xfa
    "11111010", --  226 - 0xe2  :  250 - 0xfa
    "11111010", --  227 - 0xe3  :  250 - 0xfa
    "11111001", --  228 - 0xe4  :  249 - 0xf9
    "11111010", --  229 - 0xe5  :  250 - 0xfa
    "11111010", --  230 - 0xe6  :  250 - 0xfa
    "11111010", --  231 - 0xe7  :  250 - 0xfa
    "11111010", --  232 - 0xe8  :  250 - 0xfa
    "11111010", --  233 - 0xe9  :  250 - 0xfa
    "11111010", --  234 - 0xea  :  250 - 0xfa
    "11101110", --  235 - 0xeb  :  238 - 0xee
    "11111010", --  236 - 0xec  :  250 - 0xfa
    "00100011", --  237 - 0xed  :   35 - 0x23
    "00100000", --  238 - 0xee  :   32 - 0x20
    "00100010", --  239 - 0xef  :   34 - 0x22
    "00011001", --  240 - 0xf0  :   25 - 0x19
    "00011100", --  241 - 0xf1  :   28 - 0x1c
    "00011111", --  242 - 0xf2  :   31 - 0x1f
    "11111010", --  243 - 0xf3  :  250 - 0xfa
    "11101110", --  244 - 0xf4  :  238 - 0xee
    "11111010", --  245 - 0xf5  :  250 - 0xfa
    "11111010", --  246 - 0xf6  :  250 - 0xfa
    "11111010", --  247 - 0xf7  :  250 - 0xfa
    "11111010", --  248 - 0xf8  :  250 - 0xfa
    "11111010", --  249 - 0xf9  :  250 - 0xfa
    "11111010", --  250 - 0xfa  :  250 - 0xfa
    "11111010", --  251 - 0xfb  :  250 - 0xfa
    "11111010", --  252 - 0xfc  :  250 - 0xfa
    "11111010", --  253 - 0xfd  :  250 - 0xfa
    "11111010", --  254 - 0xfe  :  250 - 0xfa
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111010", --  257 - 0x101  :  250 - 0xfa
    "11111010", --  258 - 0x102  :  250 - 0xfa
    "11111010", --  259 - 0x103  :  250 - 0xfa
    "11111010", --  260 - 0x104  :  250 - 0xfa
    "11111010", --  261 - 0x105  :  250 - 0xfa
    "11111010", --  262 - 0x106  :  250 - 0xfa
    "11111010", --  263 - 0x107  :  250 - 0xfa
    "11111010", --  264 - 0x108  :  250 - 0xfa
    "11111010", --  265 - 0x109  :  250 - 0xfa
    "11111010", --  266 - 0x10a  :  250 - 0xfa
    "11101110", --  267 - 0x10b  :  238 - 0xee
    "11111010", --  268 - 0x10c  :  250 - 0xfa
    "11111010", --  269 - 0x10d  :  250 - 0xfa
    "11111010", --  270 - 0x10e  :  250 - 0xfa
    "11111010", --  271 - 0x10f  :  250 - 0xfa
    "11111010", --  272 - 0x110  :  250 - 0xfa
    "11111010", --  273 - 0x111  :  250 - 0xfa
    "11111010", --  274 - 0x112  :  250 - 0xfa
    "11111010", --  275 - 0x113  :  250 - 0xfa
    "11101110", --  276 - 0x114  :  238 - 0xee
    "11111010", --  277 - 0x115  :  250 - 0xfa
    "11111010", --  278 - 0x116  :  250 - 0xfa
    "11111010", --  279 - 0x117  :  250 - 0xfa
    "11111010", --  280 - 0x118  :  250 - 0xfa
    "11111010", --  281 - 0x119  :  250 - 0xfa
    "11111010", --  282 - 0x11a  :  250 - 0xfa
    "11111010", --  283 - 0x11b  :  250 - 0xfa
    "11111010", --  284 - 0x11c  :  250 - 0xfa
    "11111001", --  285 - 0x11d  :  249 - 0xf9
    "11111010", --  286 - 0x11e  :  250 - 0xfa
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111010", --  289 - 0x121  :  250 - 0xfa
    "11111010", --  290 - 0x122  :  250 - 0xfa
    "11111010", --  291 - 0x123  :  250 - 0xfa
    "11111010", --  292 - 0x124  :  250 - 0xfa
    "11111010", --  293 - 0x125  :  250 - 0xfa
    "11111010", --  294 - 0x126  :  250 - 0xfa
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11111010", --  296 - 0x128  :  250 - 0xfa
    "11111010", --  297 - 0x129  :  250 - 0xfa
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11011101", --  299 - 0x12b  :  221 - 0xdd
    "11101101", --  300 - 0x12c  :  237 - 0xed
    "11101101", --  301 - 0x12d  :  237 - 0xed
    "11101101", --  302 - 0x12e  :  237 - 0xed
    "11101101", --  303 - 0x12f  :  237 - 0xed
    "11101101", --  304 - 0x130  :  237 - 0xed
    "11101101", --  305 - 0x131  :  237 - 0xed
    "11101101", --  306 - 0x132  :  237 - 0xed
    "11101101", --  307 - 0x133  :  237 - 0xed
    "11011110", --  308 - 0x134  :  222 - 0xde
    "11111010", --  309 - 0x135  :  250 - 0xfa
    "11101010", --  310 - 0x136  :  234 - 0xea
    "11111010", --  311 - 0x137  :  250 - 0xfa
    "11111010", --  312 - 0x138  :  250 - 0xfa
    "11111010", --  313 - 0x139  :  250 - 0xfa
    "11111010", --  314 - 0x13a  :  250 - 0xfa
    "11111010", --  315 - 0x13b  :  250 - 0xfa
    "11111010", --  316 - 0x13c  :  250 - 0xfa
    "11111010", --  317 - 0x13d  :  250 - 0xfa
    "11111010", --  318 - 0x13e  :  250 - 0xfa
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111010", --  321 - 0x141  :  250 - 0xfa
    "11111010", --  322 - 0x142  :  250 - 0xfa
    "11111010", --  323 - 0x143  :  250 - 0xfa
    "11111010", --  324 - 0x144  :  250 - 0xfa
    "11111010", --  325 - 0x145  :  250 - 0xfa
    "11111010", --  326 - 0x146  :  250 - 0xfa
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "11111010", --  330 - 0x14a  :  250 - 0xfa
    "11111010", --  331 - 0x14b  :  250 - 0xfa
    "11111010", --  332 - 0x14c  :  250 - 0xfa
    "11111010", --  333 - 0x14d  :  250 - 0xfa
    "11111010", --  334 - 0x14e  :  250 - 0xfa
    "11111010", --  335 - 0x14f  :  250 - 0xfa
    "11111010", --  336 - 0x150  :  250 - 0xfa
    "11111010", --  337 - 0x151  :  250 - 0xfa
    "11111010", --  338 - 0x152  :  250 - 0xfa
    "11111010", --  339 - 0x153  :  250 - 0xfa
    "11111010", --  340 - 0x154  :  250 - 0xfa
    "11111010", --  341 - 0x155  :  250 - 0xfa
    "11111010", --  342 - 0x156  :  250 - 0xfa
    "11111010", --  343 - 0x157  :  250 - 0xfa
    "11111010", --  344 - 0x158  :  250 - 0xfa
    "11111010", --  345 - 0x159  :  250 - 0xfa
    "11111010", --  346 - 0x15a  :  250 - 0xfa
    "11111010", --  347 - 0x15b  :  250 - 0xfa
    "11111010", --  348 - 0x15c  :  250 - 0xfa
    "11111010", --  349 - 0x15d  :  250 - 0xfa
    "11111010", --  350 - 0x15e  :  250 - 0xfa
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111010", --  353 - 0x161  :  250 - 0xfa
    "11111010", --  354 - 0x162  :  250 - 0xfa
    "11111010", --  355 - 0x163  :  250 - 0xfa
    "11111010", --  356 - 0x164  :  250 - 0xfa
    "11111010", --  357 - 0x165  :  250 - 0xfa
    "11111001", --  358 - 0x166  :  249 - 0xf9
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11111010", --  360 - 0x168  :  250 - 0xfa
    "11101010", --  361 - 0x169  :  234 - 0xea
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111010", --  363 - 0x16b  :  250 - 0xfa
    "11111010", --  364 - 0x16c  :  250 - 0xfa
    "11111010", --  365 - 0x16d  :  250 - 0xfa
    "11111010", --  366 - 0x16e  :  250 - 0xfa
    "11111010", --  367 - 0x16f  :  250 - 0xfa
    "11111010", --  368 - 0x170  :  250 - 0xfa
    "11111010", --  369 - 0x171  :  250 - 0xfa
    "11111010", --  370 - 0x172  :  250 - 0xfa
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111010", --  372 - 0x174  :  250 - 0xfa
    "11111010", --  373 - 0x175  :  250 - 0xfa
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11111010", --  375 - 0x177  :  250 - 0xfa
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111010", --  377 - 0x179  :  250 - 0xfa
    "11111010", --  378 - 0x17a  :  250 - 0xfa
    "11111010", --  379 - 0x17b  :  250 - 0xfa
    "11111010", --  380 - 0x17c  :  250 - 0xfa
    "11111010", --  381 - 0x17d  :  250 - 0xfa
    "11111010", --  382 - 0x17e  :  250 - 0xfa
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11111010", --  384 - 0x180  :  250 - 0xfa -- line 0xc
    "11111010", --  385 - 0x181  :  250 - 0xfa
    "11101010", --  386 - 0x182  :  234 - 0xea
    "11111010", --  387 - 0x183  :  250 - 0xfa
    "11111010", --  388 - 0x184  :  250 - 0xfa
    "11111010", --  389 - 0x185  :  250 - 0xfa
    "11111010", --  390 - 0x186  :  250 - 0xfa
    "11111010", --  391 - 0x187  :  250 - 0xfa
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11111010", --  393 - 0x189  :  250 - 0xfa
    "00100000", --  394 - 0x18a  :   32 - 0x20
    "00100010", --  395 - 0x18b  :   34 - 0x22
    "00010101", --  396 - 0x18c  :   21 - 0x15
    "00100011", --  397 - 0x18d  :   35 - 0x23
    "00100011", --  398 - 0x18e  :   35 - 0x23
    "11111010", --  399 - 0x18f  :  250 - 0xfa
    "11111010", --  400 - 0x190  :  250 - 0xfa
    "00100011", --  401 - 0x191  :   35 - 0x23
    "00100100", --  402 - 0x192  :   36 - 0x24
    "00010001", --  403 - 0x193  :   17 - 0x11
    "00100010", --  404 - 0x194  :   34 - 0x22
    "00100100", --  405 - 0x195  :   36 - 0x24
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111010", --  409 - 0x199  :  250 - 0xfa
    "11111010", --  410 - 0x19a  :  250 - 0xfa
    "11101010", --  411 - 0x19b  :  234 - 0xea
    "11111010", --  412 - 0x19c  :  250 - 0xfa
    "11111010", --  413 - 0x19d  :  250 - 0xfa
    "11111010", --  414 - 0x19e  :  250 - 0xfa
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111010", --  417 - 0x1a1  :  250 - 0xfa
    "11111010", --  418 - 0x1a2  :  250 - 0xfa
    "11111010", --  419 - 0x1a3  :  250 - 0xfa
    "11111010", --  420 - 0x1a4  :  250 - 0xfa
    "11111010", --  421 - 0x1a5  :  250 - 0xfa
    "11111010", --  422 - 0x1a6  :  250 - 0xfa
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111010", --  424 - 0x1a8  :  250 - 0xfa
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11111010", --  427 - 0x1ab  :  250 - 0xfa
    "11111010", --  428 - 0x1ac  :  250 - 0xfa
    "11111010", --  429 - 0x1ad  :  250 - 0xfa
    "11101010", --  430 - 0x1ae  :  234 - 0xea
    "11111010", --  431 - 0x1af  :  250 - 0xfa
    "11111010", --  432 - 0x1b0  :  250 - 0xfa
    "11111010", --  433 - 0x1b1  :  250 - 0xfa
    "11111010", --  434 - 0x1b2  :  250 - 0xfa
    "11111010", --  435 - 0x1b3  :  250 - 0xfa
    "11111010", --  436 - 0x1b4  :  250 - 0xfa
    "11111010", --  437 - 0x1b5  :  250 - 0xfa
    "11111010", --  438 - 0x1b6  :  250 - 0xfa
    "11111010", --  439 - 0x1b7  :  250 - 0xfa
    "11111010", --  440 - 0x1b8  :  250 - 0xfa
    "11111010", --  441 - 0x1b9  :  250 - 0xfa
    "11111010", --  442 - 0x1ba  :  250 - 0xfa
    "11111010", --  443 - 0x1bb  :  250 - 0xfa
    "11111010", --  444 - 0x1bc  :  250 - 0xfa
    "11111010", --  445 - 0x1bd  :  250 - 0xfa
    "11111010", --  446 - 0x1be  :  250 - 0xfa
    "11111010", --  447 - 0x1bf  :  250 - 0xfa
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111010", --  449 - 0x1c1  :  250 - 0xfa
    "11111010", --  450 - 0x1c2  :  250 - 0xfa
    "11111010", --  451 - 0x1c3  :  250 - 0xfa
    "11111010", --  452 - 0x1c4  :  250 - 0xfa
    "11111010", --  453 - 0x1c5  :  250 - 0xfa
    "11111010", --  454 - 0x1c6  :  250 - 0xfa
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111001", --  456 - 0x1c8  :  249 - 0xf9
    "11111010", --  457 - 0x1c9  :  250 - 0xfa
    "11111010", --  458 - 0x1ca  :  250 - 0xfa
    "11111010", --  459 - 0x1cb  :  250 - 0xfa
    "00100100", --  460 - 0x1cc  :   36 - 0x24
    "00011111", --  461 - 0x1cd  :   31 - 0x1f
    "11111010", --  462 - 0x1ce  :  250 - 0xfa
    "11111010", --  463 - 0x1cf  :  250 - 0xfa
    "00100010", --  464 - 0x1d0  :   34 - 0x22
    "00010001", --  465 - 0x1d1  :   17 - 0x11
    "00010011", --  466 - 0x1d2  :   19 - 0x13
    "00010101", --  467 - 0x1d3  :   21 - 0x15
    "11111010", --  468 - 0x1d4  :  250 - 0xfa
    "11111010", --  469 - 0x1d5  :  250 - 0xfa
    "11111010", --  470 - 0x1d6  :  250 - 0xfa
    "11111010", --  471 - 0x1d7  :  250 - 0xfa
    "11111001", --  472 - 0x1d8  :  249 - 0xf9
    "11111010", --  473 - 0x1d9  :  250 - 0xfa
    "11111010", --  474 - 0x1da  :  250 - 0xfa
    "11111010", --  475 - 0x1db  :  250 - 0xfa
    "11111010", --  476 - 0x1dc  :  250 - 0xfa
    "11111010", --  477 - 0x1dd  :  250 - 0xfa
    "11111010", --  478 - 0x1de  :  250 - 0xfa
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11111010", --  480 - 0x1e0  :  250 - 0xfa -- line 0xf
    "11111010", --  481 - 0x1e1  :  250 - 0xfa
    "11111010", --  482 - 0x1e2  :  250 - 0xfa
    "11111010", --  483 - 0x1e3  :  250 - 0xfa
    "11111010", --  484 - 0x1e4  :  250 - 0xfa
    "11111010", --  485 - 0x1e5  :  250 - 0xfa
    "11111010", --  486 - 0x1e6  :  250 - 0xfa
    "11111010", --  487 - 0x1e7  :  250 - 0xfa
    "11111010", --  488 - 0x1e8  :  250 - 0xfa
    "11111010", --  489 - 0x1e9  :  250 - 0xfa
    "11111010", --  490 - 0x1ea  :  250 - 0xfa
    "11111010", --  491 - 0x1eb  :  250 - 0xfa
    "11111010", --  492 - 0x1ec  :  250 - 0xfa
    "11111010", --  493 - 0x1ed  :  250 - 0xfa
    "11111010", --  494 - 0x1ee  :  250 - 0xfa
    "11111010", --  495 - 0x1ef  :  250 - 0xfa
    "11111010", --  496 - 0x1f0  :  250 - 0xfa
    "11111010", --  497 - 0x1f1  :  250 - 0xfa
    "11111010", --  498 - 0x1f2  :  250 - 0xfa
    "11111010", --  499 - 0x1f3  :  250 - 0xfa
    "11111010", --  500 - 0x1f4  :  250 - 0xfa
    "11111010", --  501 - 0x1f5  :  250 - 0xfa
    "11111010", --  502 - 0x1f6  :  250 - 0xfa
    "11111010", --  503 - 0x1f7  :  250 - 0xfa
    "11111010", --  504 - 0x1f8  :  250 - 0xfa
    "11111010", --  505 - 0x1f9  :  250 - 0xfa
    "11111010", --  506 - 0x1fa  :  250 - 0xfa
    "11111010", --  507 - 0x1fb  :  250 - 0xfa
    "11111010", --  508 - 0x1fc  :  250 - 0xfa
    "11111010", --  509 - 0x1fd  :  250 - 0xfa
    "11111010", --  510 - 0x1fe  :  250 - 0xfa
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111010", --  513 - 0x201  :  250 - 0xfa
    "11111010", --  514 - 0x202  :  250 - 0xfa
    "11111010", --  515 - 0x203  :  250 - 0xfa
    "11111010", --  516 - 0x204  :  250 - 0xfa
    "11111010", --  517 - 0x205  :  250 - 0xfa
    "11111010", --  518 - 0x206  :  250 - 0xfa
    "11111010", --  519 - 0x207  :  250 - 0xfa
    "11111010", --  520 - 0x208  :  250 - 0xfa
    "11111010", --  521 - 0x209  :  250 - 0xfa
    "11111010", --  522 - 0x20a  :  250 - 0xfa
    "11111010", --  523 - 0x20b  :  250 - 0xfa
    "11111010", --  524 - 0x20c  :  250 - 0xfa
    "11111010", --  525 - 0x20d  :  250 - 0xfa
    "11111010", --  526 - 0x20e  :  250 - 0xfa
    "11111010", --  527 - 0x20f  :  250 - 0xfa
    "11111010", --  528 - 0x210  :  250 - 0xfa
    "11111010", --  529 - 0x211  :  250 - 0xfa
    "11111010", --  530 - 0x212  :  250 - 0xfa
    "11111010", --  531 - 0x213  :  250 - 0xfa
    "11111010", --  532 - 0x214  :  250 - 0xfa
    "11111010", --  533 - 0x215  :  250 - 0xfa
    "11111010", --  534 - 0x216  :  250 - 0xfa
    "11111010", --  535 - 0x217  :  250 - 0xfa
    "11101001", --  536 - 0x218  :  233 - 0xe9
    "11111010", --  537 - 0x219  :  250 - 0xfa
    "11111010", --  538 - 0x21a  :  250 - 0xfa
    "11111001", --  539 - 0x21b  :  249 - 0xf9
    "11111010", --  540 - 0x21c  :  250 - 0xfa
    "11111010", --  541 - 0x21d  :  250 - 0xfa
    "11111010", --  542 - 0x21e  :  250 - 0xfa
    "11111010", --  543 - 0x21f  :  250 - 0xfa
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111010", --  545 - 0x221  :  250 - 0xfa
    "11111010", --  546 - 0x222  :  250 - 0xfa
    "11111010", --  547 - 0x223  :  250 - 0xfa
    "11111001", --  548 - 0x224  :  249 - 0xf9
    "11111010", --  549 - 0x225  :  250 - 0xfa
    "00101100", --  550 - 0x226  :   44 - 0x2c
    "00100100", --  551 - 0x227  :   36 - 0x24
    "00100010", --  552 - 0x228  :   34 - 0x22
    "00010001", --  553 - 0x229  :   17 - 0x11
    "00010011", --  554 - 0x22a  :   19 - 0x13
    "00011011", --  555 - 0x22b  :   27 - 0x1b
    "00101101", --  556 - 0x22c  :   45 - 0x2d
    "11111010", --  557 - 0x22d  :  250 - 0xfa
    "11111001", --  558 - 0x22e  :  249 - 0xf9
    "11111010", --  559 - 0x22f  :  250 - 0xfa
    "11111010", --  560 - 0x230  :  250 - 0xfa
    "11111010", --  561 - 0x231  :  250 - 0xfa
    "11111010", --  562 - 0x232  :  250 - 0xfa
    "00000001", --  563 - 0x233  :    1 - 0x1
    "11111010", --  564 - 0x234  :  250 - 0xfa
    "11111010", --  565 - 0x235  :  250 - 0xfa
    "11111010", --  566 - 0x236  :  250 - 0xfa
    "11111010", --  567 - 0x237  :  250 - 0xfa
    "11111010", --  568 - 0x238  :  250 - 0xfa
    "11111010", --  569 - 0x239  :  250 - 0xfa
    "11111010", --  570 - 0x23a  :  250 - 0xfa
    "11111010", --  571 - 0x23b  :  250 - 0xfa
    "11111010", --  572 - 0x23c  :  250 - 0xfa
    "11111010", --  573 - 0x23d  :  250 - 0xfa
    "11111010", --  574 - 0x23e  :  250 - 0xfa
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111010", --  577 - 0x241  :  250 - 0xfa
    "11111010", --  578 - 0x242  :  250 - 0xfa
    "11111010", --  579 - 0x243  :  250 - 0xfa
    "11111010", --  580 - 0x244  :  250 - 0xfa
    "11111010", --  581 - 0x245  :  250 - 0xfa
    "11101001", --  582 - 0x246  :  233 - 0xe9
    "11111010", --  583 - 0x247  :  250 - 0xfa
    "11111010", --  584 - 0x248  :  250 - 0xfa
    "11111001", --  585 - 0x249  :  249 - 0xf9
    "11111010", --  586 - 0x24a  :  250 - 0xfa
    "11111010", --  587 - 0x24b  :  250 - 0xfa
    "11111010", --  588 - 0x24c  :  250 - 0xfa
    "11111010", --  589 - 0x24d  :  250 - 0xfa
    "11111010", --  590 - 0x24e  :  250 - 0xfa
    "11111010", --  591 - 0x24f  :  250 - 0xfa
    "11111010", --  592 - 0x250  :  250 - 0xfa
    "11111010", --  593 - 0x251  :  250 - 0xfa
    "11111010", --  594 - 0x252  :  250 - 0xfa
    "11111010", --  595 - 0x253  :  250 - 0xfa
    "11111010", --  596 - 0x254  :  250 - 0xfa
    "11111010", --  597 - 0x255  :  250 - 0xfa
    "11111010", --  598 - 0x256  :  250 - 0xfa
    "11111010", --  599 - 0x257  :  250 - 0xfa
    "11111010", --  600 - 0x258  :  250 - 0xfa
    "11111010", --  601 - 0x259  :  250 - 0xfa
    "11111010", --  602 - 0x25a  :  250 - 0xfa
    "11111010", --  603 - 0x25b  :  250 - 0xfa
    "11111010", --  604 - 0x25c  :  250 - 0xfa
    "11111010", --  605 - 0x25d  :  250 - 0xfa
    "11111010", --  606 - 0x25e  :  250 - 0xfa
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa -- line 0x13
    "11111010", --  609 - 0x261  :  250 - 0xfa
    "11111010", --  610 - 0x262  :  250 - 0xfa
    "11111010", --  611 - 0x263  :  250 - 0xfa
    "11111010", --  612 - 0x264  :  250 - 0xfa
    "11111010", --  613 - 0x265  :  250 - 0xfa
    "11111010", --  614 - 0x266  :  250 - 0xfa
    "00010100", --  615 - 0x267  :   20 - 0x14
    "00011001", --  616 - 0x268  :   25 - 0x19
    "00010110", --  617 - 0x269  :   22 - 0x16
    "00010110", --  618 - 0x26a  :   22 - 0x16
    "00011001", --  619 - 0x26b  :   25 - 0x19
    "00010011", --  620 - 0x26c  :   19 - 0x13
    "00100101", --  621 - 0x26d  :   37 - 0x25
    "00011100", --  622 - 0x26e  :   28 - 0x1c
    "00100100", --  623 - 0x26f  :   36 - 0x24
    "00101001", --  624 - 0x270  :   41 - 0x29
    "00101101", --  625 - 0x271  :   45 - 0x2d
    "11111010", --  626 - 0x272  :  250 - 0xfa
    "00011000", --  627 - 0x273  :   24 - 0x18
    "00010001", --  628 - 0x274  :   17 - 0x11
    "00100010", --  629 - 0x275  :   34 - 0x22
    "00010100", --  630 - 0x276  :   20 - 0x14
    "11111010", --  631 - 0x277  :  250 - 0xfa
    "11111010", --  632 - 0x278  :  250 - 0xfa
    "11111010", --  633 - 0x279  :  250 - 0xfa
    "11111010", --  634 - 0x27a  :  250 - 0xfa
    "11111010", --  635 - 0x27b  :  250 - 0xfa
    "11111010", --  636 - 0x27c  :  250 - 0xfa
    "11111010", --  637 - 0x27d  :  250 - 0xfa
    "11111001", --  638 - 0x27e  :  249 - 0xf9
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111010", --  641 - 0x281  :  250 - 0xfa
    "11101001", --  642 - 0x282  :  233 - 0xe9
    "11111010", --  643 - 0x283  :  250 - 0xfa
    "11111010", --  644 - 0x284  :  250 - 0xfa
    "11111010", --  645 - 0x285  :  250 - 0xfa
    "11111010", --  646 - 0x286  :  250 - 0xfa
    "11111001", --  647 - 0x287  :  249 - 0xf9
    "11111001", --  648 - 0x288  :  249 - 0xf9
    "11111010", --  649 - 0x289  :  250 - 0xfa
    "11111010", --  650 - 0x28a  :  250 - 0xfa
    "11111010", --  651 - 0x28b  :  250 - 0xfa
    "11111010", --  652 - 0x28c  :  250 - 0xfa
    "11111010", --  653 - 0x28d  :  250 - 0xfa
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "11111010", --  655 - 0x28f  :  250 - 0xfa
    "11111010", --  656 - 0x290  :  250 - 0xfa
    "11111010", --  657 - 0x291  :  250 - 0xfa
    "11111010", --  658 - 0x292  :  250 - 0xfa
    "11101001", --  659 - 0x293  :  233 - 0xe9
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "11111010", --  661 - 0x295  :  250 - 0xfa
    "11111010", --  662 - 0x296  :  250 - 0xfa
    "11111010", --  663 - 0x297  :  250 - 0xfa
    "11101010", --  664 - 0x298  :  234 - 0xea
    "11111010", --  665 - 0x299  :  250 - 0xfa
    "11111010", --  666 - 0x29a  :  250 - 0xfa
    "11111010", --  667 - 0x29b  :  250 - 0xfa
    "11111010", --  668 - 0x29c  :  250 - 0xfa
    "11111010", --  669 - 0x29d  :  250 - 0xfa
    "11111010", --  670 - 0x29e  :  250 - 0xfa
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111010", --  673 - 0x2a1  :  250 - 0xfa
    "11111010", --  674 - 0x2a2  :  250 - 0xfa
    "11111010", --  675 - 0x2a3  :  250 - 0xfa
    "11111010", --  676 - 0x2a4  :  250 - 0xfa
    "11111010", --  677 - 0x2a5  :  250 - 0xfa
    "11111010", --  678 - 0x2a6  :  250 - 0xfa
    "00011100", --  679 - 0x2a7  :   28 - 0x1c
    "00010001", --  680 - 0x2a8  :   17 - 0x11
    "00100000", --  681 - 0x2a9  :   32 - 0x20
    "00100011", --  682 - 0x2aa  :   35 - 0x23
    "00101101", --  683 - 0x2ab  :   45 - 0x2d
    "11111010", --  684 - 0x2ac  :  250 - 0xfa
    "11111010", --  685 - 0x2ad  :  250 - 0xfa
    "11111010", --  686 - 0x2ae  :  250 - 0xfa
    "11101010", --  687 - 0x2af  :  234 - 0xea
    "11111010", --  688 - 0x2b0  :  250 - 0xfa
    "11111010", --  689 - 0x2b1  :  250 - 0xfa
    "11111010", --  690 - 0x2b2  :  250 - 0xfa
    "00000011", --  691 - 0x2b3  :    3 - 0x3
    "11111010", --  692 - 0x2b4  :  250 - 0xfa
    "11111010", --  693 - 0x2b5  :  250 - 0xfa
    "11111010", --  694 - 0x2b6  :  250 - 0xfa
    "11111010", --  695 - 0x2b7  :  250 - 0xfa
    "11111010", --  696 - 0x2b8  :  250 - 0xfa
    "11111010", --  697 - 0x2b9  :  250 - 0xfa
    "11111010", --  698 - 0x2ba  :  250 - 0xfa
    "11111010", --  699 - 0x2bb  :  250 - 0xfa
    "11111010", --  700 - 0x2bc  :  250 - 0xfa
    "11111010", --  701 - 0x2bd  :  250 - 0xfa
    "11111010", --  702 - 0x2be  :  250 - 0xfa
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111010", --  705 - 0x2c1  :  250 - 0xfa
    "11111010", --  706 - 0x2c2  :  250 - 0xfa
    "11111010", --  707 - 0x2c3  :  250 - 0xfa
    "11111010", --  708 - 0x2c4  :  250 - 0xfa
    "11111010", --  709 - 0x2c5  :  250 - 0xfa
    "11111010", --  710 - 0x2c6  :  250 - 0xfa
    "11111010", --  711 - 0x2c7  :  250 - 0xfa
    "11111010", --  712 - 0x2c8  :  250 - 0xfa
    "11111010", --  713 - 0x2c9  :  250 - 0xfa
    "11111010", --  714 - 0x2ca  :  250 - 0xfa
    "11111010", --  715 - 0x2cb  :  250 - 0xfa
    "11111010", --  716 - 0x2cc  :  250 - 0xfa
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11111010", --  718 - 0x2ce  :  250 - 0xfa
    "11111010", --  719 - 0x2cf  :  250 - 0xfa
    "11111010", --  720 - 0x2d0  :  250 - 0xfa
    "11111010", --  721 - 0x2d1  :  250 - 0xfa
    "11111010", --  722 - 0x2d2  :  250 - 0xfa
    "11111010", --  723 - 0x2d3  :  250 - 0xfa
    "11111010", --  724 - 0x2d4  :  250 - 0xfa
    "11111010", --  725 - 0x2d5  :  250 - 0xfa
    "11111010", --  726 - 0x2d6  :  250 - 0xfa
    "11111010", --  727 - 0x2d7  :  250 - 0xfa
    "11111010", --  728 - 0x2d8  :  250 - 0xfa
    "11111010", --  729 - 0x2d9  :  250 - 0xfa
    "11111010", --  730 - 0x2da  :  250 - 0xfa
    "11111010", --  731 - 0x2db  :  250 - 0xfa
    "11111010", --  732 - 0x2dc  :  250 - 0xfa
    "11101010", --  733 - 0x2dd  :  234 - 0xea
    "11111010", --  734 - 0x2de  :  250 - 0xfa
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111011", --  736 - 0x2e0  :  251 - 0xfb -- line 0x17
    "11111011", --  737 - 0x2e1  :  251 - 0xfb
    "11111011", --  738 - 0x2e2  :  251 - 0xfb
    "11111011", --  739 - 0x2e3  :  251 - 0xfb
    "11111011", --  740 - 0x2e4  :  251 - 0xfb
    "11111011", --  741 - 0x2e5  :  251 - 0xfb
    "11111011", --  742 - 0x2e6  :  251 - 0xfb
    "11111011", --  743 - 0x2e7  :  251 - 0xfb
    "11111011", --  744 - 0x2e8  :  251 - 0xfb
    "11111011", --  745 - 0x2e9  :  251 - 0xfb
    "11111011", --  746 - 0x2ea  :  251 - 0xfb
    "11111011", --  747 - 0x2eb  :  251 - 0xfb
    "11111011", --  748 - 0x2ec  :  251 - 0xfb
    "11111011", --  749 - 0x2ed  :  251 - 0xfb
    "11111011", --  750 - 0x2ee  :  251 - 0xfb
    "11111011", --  751 - 0x2ef  :  251 - 0xfb
    "11111011", --  752 - 0x2f0  :  251 - 0xfb
    "11111011", --  753 - 0x2f1  :  251 - 0xfb
    "11111011", --  754 - 0x2f2  :  251 - 0xfb
    "11111011", --  755 - 0x2f3  :  251 - 0xfb
    "11111011", --  756 - 0x2f4  :  251 - 0xfb
    "11111011", --  757 - 0x2f5  :  251 - 0xfb
    "11111011", --  758 - 0x2f6  :  251 - 0xfb
    "11111011", --  759 - 0x2f7  :  251 - 0xfb
    "11111011", --  760 - 0x2f8  :  251 - 0xfb
    "11111011", --  761 - 0x2f9  :  251 - 0xfb
    "11111011", --  762 - 0x2fa  :  251 - 0xfb
    "11111011", --  763 - 0x2fb  :  251 - 0xfb
    "11111011", --  764 - 0x2fc  :  251 - 0xfb
    "11111011", --  765 - 0x2fd  :  251 - 0xfb
    "11111011", --  766 - 0x2fe  :  251 - 0xfb
    "11111011", --  767 - 0x2ff  :  251 - 0xfb
    "11111111", --  768 - 0x300  :  255 - 0xff -- line 0x18
    "11111111", --  769 - 0x301  :  255 - 0xff
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11111111", --  772 - 0x304  :  255 - 0xff
    "11111111", --  773 - 0x305  :  255 - 0xff
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff
    "11111111", --  793 - 0x319  :  255 - 0xff
    "11111111", --  794 - 0x31a  :  255 - 0xff
    "11111111", --  795 - 0x31b  :  255 - 0xff
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11111111", --  798 - 0x31e  :  255 - 0xff
    "11111111", --  799 - 0x31f  :  255 - 0xff
    "11111111", --  800 - 0x320  :  255 - 0xff -- line 0x19
    "11111101", --  801 - 0x321  :  253 - 0xfd
    "11111111", --  802 - 0x322  :  255 - 0xff
    "11111101", --  803 - 0x323  :  253 - 0xfd
    "11111111", --  804 - 0x324  :  255 - 0xff
    "11111101", --  805 - 0x325  :  253 - 0xfd
    "11111111", --  806 - 0x326  :  255 - 0xff
    "11111101", --  807 - 0x327  :  253 - 0xfd
    "11111111", --  808 - 0x328  :  255 - 0xff
    "11111101", --  809 - 0x329  :  253 - 0xfd
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "11111101", --  811 - 0x32b  :  253 - 0xfd
    "11111111", --  812 - 0x32c  :  255 - 0xff
    "11111101", --  813 - 0x32d  :  253 - 0xfd
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111101", --  815 - 0x32f  :  253 - 0xfd
    "11111111", --  816 - 0x330  :  255 - 0xff
    "11111101", --  817 - 0x331  :  253 - 0xfd
    "11111111", --  818 - 0x332  :  255 - 0xff
    "11111101", --  819 - 0x333  :  253 - 0xfd
    "11111111", --  820 - 0x334  :  255 - 0xff
    "11111101", --  821 - 0x335  :  253 - 0xfd
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111101", --  823 - 0x337  :  253 - 0xfd
    "11111111", --  824 - 0x338  :  255 - 0xff
    "11111101", --  825 - 0x339  :  253 - 0xfd
    "11111111", --  826 - 0x33a  :  255 - 0xff
    "11111101", --  827 - 0x33b  :  253 - 0xfd
    "11111111", --  828 - 0x33c  :  255 - 0xff
    "11111101", --  829 - 0x33d  :  253 - 0xfd
    "11111111", --  830 - 0x33e  :  255 - 0xff
    "11111101", --  831 - 0x33f  :  253 - 0xfd
    "11111111", --  832 - 0x340  :  255 - 0xff -- line 0x1a
    "11111101", --  833 - 0x341  :  253 - 0xfd
    "11111111", --  834 - 0x342  :  255 - 0xff
    "11111101", --  835 - 0x343  :  253 - 0xfd
    "11111111", --  836 - 0x344  :  255 - 0xff
    "11111101", --  837 - 0x345  :  253 - 0xfd
    "11111111", --  838 - 0x346  :  255 - 0xff
    "11111101", --  839 - 0x347  :  253 - 0xfd
    "11111111", --  840 - 0x348  :  255 - 0xff
    "11111101", --  841 - 0x349  :  253 - 0xfd
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111101", --  843 - 0x34b  :  253 - 0xfd
    "11111111", --  844 - 0x34c  :  255 - 0xff
    "11111101", --  845 - 0x34d  :  253 - 0xfd
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111101", --  847 - 0x34f  :  253 - 0xfd
    "11111111", --  848 - 0x350  :  255 - 0xff
    "11111101", --  849 - 0x351  :  253 - 0xfd
    "11111111", --  850 - 0x352  :  255 - 0xff
    "11111101", --  851 - 0x353  :  253 - 0xfd
    "11111111", --  852 - 0x354  :  255 - 0xff
    "11111101", --  853 - 0x355  :  253 - 0xfd
    "11111111", --  854 - 0x356  :  255 - 0xff
    "11111101", --  855 - 0x357  :  253 - 0xfd
    "11111111", --  856 - 0x358  :  255 - 0xff
    "11111101", --  857 - 0x359  :  253 - 0xfd
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111101", --  859 - 0x35b  :  253 - 0xfd
    "11111111", --  860 - 0x35c  :  255 - 0xff
    "11111101", --  861 - 0x35d  :  253 - 0xfd
    "11111111", --  862 - 0x35e  :  255 - 0xff
    "11111101", --  863 - 0x35f  :  253 - 0xfd
    "11111111", --  864 - 0x360  :  255 - 0xff -- line 0x1b
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111111", --  870 - 0x366  :  255 - 0xff
    "11111111", --  871 - 0x367  :  255 - 0xff
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11111111", --  882 - 0x372  :  255 - 0xff
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11111111", --  892 - 0x37c  :  255 - 0xff
    "11111111", --  893 - 0x37d  :  255 - 0xff
    "11111111", --  894 - 0x37e  :  255 - 0xff
    "11111111", --  895 - 0x37f  :  255 - 0xff
    "11101011", --  896 - 0x380  :  235 - 0xeb -- line 0x1c
    "11101011", --  897 - 0x381  :  235 - 0xeb
    "11101011", --  898 - 0x382  :  235 - 0xeb
    "11101011", --  899 - 0x383  :  235 - 0xeb
    "11101011", --  900 - 0x384  :  235 - 0xeb
    "11101011", --  901 - 0x385  :  235 - 0xeb
    "11101011", --  902 - 0x386  :  235 - 0xeb
    "11101011", --  903 - 0x387  :  235 - 0xeb
    "11101011", --  904 - 0x388  :  235 - 0xeb
    "11101011", --  905 - 0x389  :  235 - 0xeb
    "11101011", --  906 - 0x38a  :  235 - 0xeb
    "11101011", --  907 - 0x38b  :  235 - 0xeb
    "11101011", --  908 - 0x38c  :  235 - 0xeb
    "11101011", --  909 - 0x38d  :  235 - 0xeb
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11101011", --  922 - 0x39a  :  235 - 0xeb
    "11101011", --  923 - 0x39b  :  235 - 0xeb
    "11101011", --  924 - 0x39c  :  235 - 0xeb
    "11101011", --  925 - 0x39d  :  235 - 0xeb
    "11101011", --  926 - 0x39e  :  235 - 0xeb
    "11101011", --  927 - 0x39f  :  235 - 0xeb
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111010", --  929 - 0x3a1  :  250 - 0xfa
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11101010", --  943 - 0x3af  :  234 - 0xea
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11111010", --  949 - 0x3b5  :  250 - 0xfa
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11111010", --  956 - 0x3bc  :  250 - 0xfa
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111001", --  959 - 0x3bf  :  249 - 0xf9
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "01010101", --  961 - 0x3c1  :   85 - 0x55
    "01010101", --  962 - 0x3c2  :   85 - 0x55
    "01010101", --  963 - 0x3c3  :   85 - 0x55
    "01010101", --  964 - 0x3c4  :   85 - 0x55
    "01010101", --  965 - 0x3c5  :   85 - 0x55
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "01010101", --  968 - 0x3c8  :   85 - 0x55
    "01010101", --  969 - 0x3c9  :   85 - 0x55
    "01010101", --  970 - 0x3ca  :   85 - 0x55
    "01010101", --  971 - 0x3cb  :   85 - 0x55
    "01010101", --  972 - 0x3cc  :   85 - 0x55
    "01010101", --  973 - 0x3cd  :   85 - 0x55
    "01010101", --  974 - 0x3ce  :   85 - 0x55
    "01010101", --  975 - 0x3cf  :   85 - 0x55
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "01010101", --  977 - 0x3d1  :   85 - 0x55
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "01010101", --  982 - 0x3d6  :   85 - 0x55
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "01010101", --  990 - 0x3de  :   85 - 0x55
    "01010101", --  991 - 0x3df  :   85 - 0x55
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "01010101", --  997 - 0x3e5  :   85 - 0x55
    "01010101", --  998 - 0x3e6  :   85 - 0x55
    "01010101", --  999 - 0x3e7  :   85 - 0x55
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "01010101", -- 1002 - 0x3ea  :   85 - 0x55
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "01010101", -- 1005 - 0x3ed  :   85 - 0x55
    "01010101", -- 1006 - 0x3ee  :   85 - 0x55
    "01010101", -- 1007 - 0x3ef  :   85 - 0x55
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
