--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_racet3.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_RACE3 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_RACE3;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_RACE3 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11101001", --   22 - 0x16  :  233 - 0xe9
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11101010", --   28 - 0x1c  :  234 - 0xea
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11111010", --   33 - 0x21  :  250 - 0xfa
    "11111010", --   34 - 0x22  :  250 - 0xfa
    "11100111", --   35 - 0x23  :  231 - 0xe7
    "11111011", --   36 - 0x24  :  251 - 0xfb
    "11111011", --   37 - 0x25  :  251 - 0xfb
    "11111011", --   38 - 0x26  :  251 - 0xfb
    "11111011", --   39 - 0x27  :  251 - 0xfb
    "11111011", --   40 - 0x28  :  251 - 0xfb
    "11111011", --   41 - 0x29  :  251 - 0xfb
    "11111011", --   42 - 0x2a  :  251 - 0xfb
    "11111011", --   43 - 0x2b  :  251 - 0xfb
    "11111011", --   44 - 0x2c  :  251 - 0xfb
    "11111011", --   45 - 0x2d  :  251 - 0xfb
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111011", --   47 - 0x2f  :  251 - 0xfb
    "11101000", --   48 - 0x30  :  232 - 0xe8
    "11111010", --   49 - 0x31  :  250 - 0xfa
    "11101010", --   50 - 0x32  :  234 - 0xea
    "11111010", --   51 - 0x33  :  250 - 0xfa
    "11111010", --   52 - 0x34  :  250 - 0xfa
    "11111010", --   53 - 0x35  :  250 - 0xfa
    "11111010", --   54 - 0x36  :  250 - 0xfa
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11111001", --   57 - 0x39  :  249 - 0xf9
    "11111010", --   58 - 0x3a  :  250 - 0xfa
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11101010", --   63 - 0x3f  :  234 - 0xea
    "11101010", --   64 - 0x40  :  234 - 0xea -- line 0x2
    "11111010", --   65 - 0x41  :  250 - 0xfa
    "11111010", --   66 - 0x42  :  250 - 0xfa
    "11111100", --   67 - 0x43  :  252 - 0xfc
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11111111", --   70 - 0x46  :  255 - 0xff
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11101100", --   80 - 0x50  :  236 - 0xec
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111001", --   83 - 0x53  :  249 - 0xf9
    "11111010", --   84 - 0x54  :  250 - 0xfa
    "11111010", --   85 - 0x55  :  250 - 0xfa
    "11101001", --   86 - 0x56  :  233 - 0xe9
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11101010", --   91 - 0x5b  :  234 - 0xea
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11101001", --   93 - 0x5d  :  233 - 0xe9
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11100111", --   97 - 0x61  :  231 - 0xe7
    "11111011", --   98 - 0x62  :  251 - 0xfb
    "11110110", --   99 - 0x63  :  246 - 0xf6
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111101", --  102 - 0x66  :  253 - 0xfd
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11111101", --  104 - 0x68  :  253 - 0xfd
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111101", --  106 - 0x6a  :  253 - 0xfd
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111101", --  108 - 0x6c  :  253 - 0xfd
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11111111", --  110 - 0x6e  :  255 - 0xff
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11101100", --  112 - 0x70  :  236 - 0xec
    "11111010", --  113 - 0x71  :  250 - 0xfa
    "11111010", --  114 - 0x72  :  250 - 0xfa
    "11111010", --  115 - 0x73  :  250 - 0xfa
    "11111010", --  116 - 0x74  :  250 - 0xfa
    "11111010", --  117 - 0x75  :  250 - 0xfa
    "11111010", --  118 - 0x76  :  250 - 0xfa
    "11111010", --  119 - 0x77  :  250 - 0xfa
    "11101001", --  120 - 0x78  :  233 - 0xe9
    "11111010", --  121 - 0x79  :  250 - 0xfa
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11101001", --  128 - 0x80  :  233 - 0xe9 -- line 0x4
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111111", --  130 - 0x82  :  255 - 0xff
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111101", --  134 - 0x86  :  253 - 0xfd
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111101", --  136 - 0x88  :  253 - 0xfd
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11111101", --  138 - 0x8a  :  253 - 0xfd
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111101", --  140 - 0x8c  :  253 - 0xfd
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11111111", --  142 - 0x8e  :  255 - 0xff
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11101100", --  144 - 0x90  :  236 - 0xec
    "11111010", --  145 - 0x91  :  250 - 0xfa
    "11111010", --  146 - 0x92  :  250 - 0xfa
    "11101001", --  147 - 0x93  :  233 - 0xe9
    "11111010", --  148 - 0x94  :  250 - 0xfa
    "11111010", --  149 - 0x95  :  250 - 0xfa
    "11111010", --  150 - 0x96  :  250 - 0xfa
    "11111010", --  151 - 0x97  :  250 - 0xfa
    "11111010", --  152 - 0x98  :  250 - 0xfa
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11111010", --  154 - 0x9a  :  250 - 0xfa
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111010", --  156 - 0x9c  :  250 - 0xfa
    "11111010", --  157 - 0x9d  :  250 - 0xfa
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111100", --  161 - 0xa1  :  252 - 0xfc
    "11111111", --  162 - 0xa2  :  255 - 0xff
    "11111111", --  163 - 0xa3  :  255 - 0xff
    "11111111", --  164 - 0xa4  :  255 - 0xff
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11111111", --  175 - 0xaf  :  255 - 0xff
    "11101100", --  176 - 0xb0  :  236 - 0xec
    "11111010", --  177 - 0xb1  :  250 - 0xfa
    "11111010", --  178 - 0xb2  :  250 - 0xfa
    "11111010", --  179 - 0xb3  :  250 - 0xfa
    "11111010", --  180 - 0xb4  :  250 - 0xfa
    "11111010", --  181 - 0xb5  :  250 - 0xfa
    "11101010", --  182 - 0xb6  :  234 - 0xea
    "11111010", --  183 - 0xb7  :  250 - 0xfa
    "11111001", --  184 - 0xb8  :  249 - 0xf9
    "11111010", --  185 - 0xb9  :  250 - 0xfa
    "11111010", --  186 - 0xba  :  250 - 0xfa
    "11101001", --  187 - 0xbb  :  233 - 0xe9
    "11111010", --  188 - 0xbc  :  250 - 0xfa
    "11111010", --  189 - 0xbd  :  250 - 0xfa
    "11111010", --  190 - 0xbe  :  250 - 0xfa
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa -- line 0x6
    "11111100", --  193 - 0xc1  :  252 - 0xfc
    "11111111", --  194 - 0xc2  :  255 - 0xff
    "11111110", --  195 - 0xc3  :  254 - 0xfe
    "11111110", --  196 - 0xc4  :  254 - 0xfe
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11100101", --  198 - 0xc6  :  229 - 0xe5
    "11101011", --  199 - 0xc7  :  235 - 0xeb
    "11101011", --  200 - 0xc8  :  235 - 0xeb
    "11101011", --  201 - 0xc9  :  235 - 0xeb
    "11101011", --  202 - 0xca  :  235 - 0xeb
    "11100110", --  203 - 0xcb  :  230 - 0xe6
    "11111111", --  204 - 0xcc  :  255 - 0xff
    "11111110", --  205 - 0xcd  :  254 - 0xfe
    "11111110", --  206 - 0xce  :  254 - 0xfe
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "11101100", --  208 - 0xd0  :  236 - 0xec
    "11111010", --  209 - 0xd1  :  250 - 0xfa
    "11111001", --  210 - 0xd2  :  249 - 0xf9
    "11111010", --  211 - 0xd3  :  250 - 0xfa
    "11111010", --  212 - 0xd4  :  250 - 0xfa
    "11111010", --  213 - 0xd5  :  250 - 0xfa
    "11111010", --  214 - 0xd6  :  250 - 0xfa
    "11111010", --  215 - 0xd7  :  250 - 0xfa
    "11111010", --  216 - 0xd8  :  250 - 0xfa
    "11111001", --  217 - 0xd9  :  249 - 0xf9
    "11111010", --  218 - 0xda  :  250 - 0xfa
    "11111010", --  219 - 0xdb  :  250 - 0xfa
    "11111010", --  220 - 0xdc  :  250 - 0xfa
    "11111010", --  221 - 0xdd  :  250 - 0xfa
    "11111010", --  222 - 0xde  :  250 - 0xfa
    "11101010", --  223 - 0xdf  :  234 - 0xea
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111100", --  225 - 0xe1  :  252 - 0xfc
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111111", --  227 - 0xe3  :  255 - 0xff
    "11111111", --  228 - 0xe4  :  255 - 0xff
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11101100", --  230 - 0xe6  :  236 - 0xec
    "11111010", --  231 - 0xe7  :  250 - 0xfa
    "11111010", --  232 - 0xe8  :  250 - 0xfa
    "11111010", --  233 - 0xe9  :  250 - 0xfa
    "11111010", --  234 - 0xea  :  250 - 0xfa
    "11111100", --  235 - 0xeb  :  252 - 0xfc
    "11111111", --  236 - 0xec  :  255 - 0xff
    "11111111", --  237 - 0xed  :  255 - 0xff
    "11111111", --  238 - 0xee  :  255 - 0xff
    "11111111", --  239 - 0xef  :  255 - 0xff
    "11101100", --  240 - 0xf0  :  236 - 0xec
    "11111010", --  241 - 0xf1  :  250 - 0xfa
    "11111010", --  242 - 0xf2  :  250 - 0xfa
    "11111010", --  243 - 0xf3  :  250 - 0xfa
    "11111010", --  244 - 0xf4  :  250 - 0xfa
    "11111010", --  245 - 0xf5  :  250 - 0xfa
    "11111010", --  246 - 0xf6  :  250 - 0xfa
    "11111010", --  247 - 0xf7  :  250 - 0xfa
    "11111010", --  248 - 0xf8  :  250 - 0xfa
    "11111010", --  249 - 0xf9  :  250 - 0xfa
    "11101010", --  250 - 0xfa  :  234 - 0xea
    "11111010", --  251 - 0xfb  :  250 - 0xfa
    "11111001", --  252 - 0xfc  :  249 - 0xf9
    "11111010", --  253 - 0xfd  :  250 - 0xfa
    "11111010", --  254 - 0xfe  :  250 - 0xfa
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111100", --  257 - 0x101  :  252 - 0xfc
    "11111111", --  258 - 0x102  :  255 - 0xff
    "11111110", --  259 - 0x103  :  254 - 0xfe
    "11111110", --  260 - 0x104  :  254 - 0xfe
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11101100", --  262 - 0x106  :  236 - 0xec
    "11111010", --  263 - 0x107  :  250 - 0xfa
    "11111001", --  264 - 0x108  :  249 - 0xf9
    "11111010", --  265 - 0x109  :  250 - 0xfa
    "11111010", --  266 - 0x10a  :  250 - 0xfa
    "11111100", --  267 - 0x10b  :  252 - 0xfc
    "11111111", --  268 - 0x10c  :  255 - 0xff
    "11111110", --  269 - 0x10d  :  254 - 0xfe
    "11111110", --  270 - 0x10e  :  254 - 0xfe
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "11101100", --  272 - 0x110  :  236 - 0xec
    "11111010", --  273 - 0x111  :  250 - 0xfa
    "11111010", --  274 - 0x112  :  250 - 0xfa
    "11101001", --  275 - 0x113  :  233 - 0xe9
    "11111010", --  276 - 0x114  :  250 - 0xfa
    "11101010", --  277 - 0x115  :  234 - 0xea
    "11111010", --  278 - 0x116  :  250 - 0xfa
    "11111010", --  279 - 0x117  :  250 - 0xfa
    "11101001", --  280 - 0x118  :  233 - 0xe9
    "11111010", --  281 - 0x119  :  250 - 0xfa
    "11111010", --  282 - 0x11a  :  250 - 0xfa
    "11101010", --  283 - 0x11b  :  234 - 0xea
    "11111010", --  284 - 0x11c  :  250 - 0xfa
    "11111010", --  285 - 0x11d  :  250 - 0xfa
    "11101001", --  286 - 0x11e  :  233 - 0xe9
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111100", --  289 - 0x121  :  252 - 0xfc
    "11111111", --  290 - 0x122  :  255 - 0xff
    "11111111", --  291 - 0x123  :  255 - 0xff
    "11111111", --  292 - 0x124  :  255 - 0xff
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11101100", --  294 - 0x126  :  236 - 0xec
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11101001", --  296 - 0x128  :  233 - 0xe9
    "11111010", --  297 - 0x129  :  250 - 0xfa
    "11101010", --  298 - 0x12a  :  234 - 0xea
    "11111100", --  299 - 0x12b  :  252 - 0xfc
    "11111111", --  300 - 0x12c  :  255 - 0xff
    "11111111", --  301 - 0x12d  :  255 - 0xff
    "11111111", --  302 - 0x12e  :  255 - 0xff
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "11101100", --  304 - 0x130  :  236 - 0xec
    "11111010", --  305 - 0x131  :  250 - 0xfa
    "11111010", --  306 - 0x132  :  250 - 0xfa
    "11111010", --  307 - 0x133  :  250 - 0xfa
    "11111010", --  308 - 0x134  :  250 - 0xfa
    "11111010", --  309 - 0x135  :  250 - 0xfa
    "11111010", --  310 - 0x136  :  250 - 0xfa
    "11111010", --  311 - 0x137  :  250 - 0xfa
    "11111010", --  312 - 0x138  :  250 - 0xfa
    "11111010", --  313 - 0x139  :  250 - 0xfa
    "11111010", --  314 - 0x13a  :  250 - 0xfa
    "11111010", --  315 - 0x13b  :  250 - 0xfa
    "11111010", --  316 - 0x13c  :  250 - 0xfa
    "11111010", --  317 - 0x13d  :  250 - 0xfa
    "11111010", --  318 - 0x13e  :  250 - 0xfa
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111100", --  321 - 0x141  :  252 - 0xfc
    "11111111", --  322 - 0x142  :  255 - 0xff
    "11111110", --  323 - 0x143  :  254 - 0xfe
    "11111110", --  324 - 0x144  :  254 - 0xfe
    "11111111", --  325 - 0x145  :  255 - 0xff
    "11101100", --  326 - 0x146  :  236 - 0xec
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "11111010", --  330 - 0x14a  :  250 - 0xfa
    "11111100", --  331 - 0x14b  :  252 - 0xfc
    "11111111", --  332 - 0x14c  :  255 - 0xff
    "11111110", --  333 - 0x14d  :  254 - 0xfe
    "11111110", --  334 - 0x14e  :  254 - 0xfe
    "11111111", --  335 - 0x14f  :  255 - 0xff
    "11101100", --  336 - 0x150  :  236 - 0xec
    "11101001", --  337 - 0x151  :  233 - 0xe9
    "11111010", --  338 - 0x152  :  250 - 0xfa
    "11111010", --  339 - 0x153  :  250 - 0xfa
    "11111010", --  340 - 0x154  :  250 - 0xfa
    "11111010", --  341 - 0x155  :  250 - 0xfa
    "11111010", --  342 - 0x156  :  250 - 0xfa
    "11111001", --  343 - 0x157  :  249 - 0xf9
    "11111001", --  344 - 0x158  :  249 - 0xf9
    "11111001", --  345 - 0x159  :  249 - 0xf9
    "11111010", --  346 - 0x15a  :  250 - 0xfa
    "11111010", --  347 - 0x15b  :  250 - 0xfa
    "11111010", --  348 - 0x15c  :  250 - 0xfa
    "11111010", --  349 - 0x15d  :  250 - 0xfa
    "11111010", --  350 - 0x15e  :  250 - 0xfa
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111100", --  353 - 0x161  :  252 - 0xfc
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111111", --  355 - 0x163  :  255 - 0xff
    "11111111", --  356 - 0x164  :  255 - 0xff
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11101100", --  358 - 0x166  :  236 - 0xec
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11101010", --  360 - 0x168  :  234 - 0xea
    "11111010", --  361 - 0x169  :  250 - 0xfa
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111100", --  363 - 0x16b  :  252 - 0xfc
    "11111111", --  364 - 0x16c  :  255 - 0xff
    "11111111", --  365 - 0x16d  :  255 - 0xff
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "11110101", --  368 - 0x170  :  245 - 0xf5
    "11111011", --  369 - 0x171  :  251 - 0xfb
    "11101000", --  370 - 0x172  :  232 - 0xe8
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111001", --  372 - 0x174  :  249 - 0xf9
    "11101001", --  373 - 0x175  :  233 - 0xe9
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11111001", --  375 - 0x177  :  249 - 0xf9
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111010", --  377 - 0x179  :  250 - 0xfa
    "11111010", --  378 - 0x17a  :  250 - 0xfa
    "11101001", --  379 - 0x17b  :  233 - 0xe9
    "11111010", --  380 - 0x17c  :  250 - 0xfa
    "11101010", --  381 - 0x17d  :  234 - 0xea
    "11111010", --  382 - 0x17e  :  250 - 0xfa
    "11101001", --  383 - 0x17f  :  233 - 0xe9
    "11101001", --  384 - 0x180  :  233 - 0xe9 -- line 0xc
    "11111100", --  385 - 0x181  :  252 - 0xfc
    "11111111", --  386 - 0x182  :  255 - 0xff
    "11111110", --  387 - 0x183  :  254 - 0xfe
    "11111110", --  388 - 0x184  :  254 - 0xfe
    "11111111", --  389 - 0x185  :  255 - 0xff
    "11101100", --  390 - 0x186  :  236 - 0xec
    "11101010", --  391 - 0x187  :  234 - 0xea
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11101010", --  393 - 0x189  :  234 - 0xea
    "11111010", --  394 - 0x18a  :  250 - 0xfa
    "11111100", --  395 - 0x18b  :  252 - 0xfc
    "11111111", --  396 - 0x18c  :  255 - 0xff
    "11111110", --  397 - 0x18d  :  254 - 0xfe
    "11111110", --  398 - 0x18e  :  254 - 0xfe
    "11111111", --  399 - 0x18f  :  255 - 0xff
    "11111111", --  400 - 0x190  :  255 - 0xff
    "11111111", --  401 - 0x191  :  255 - 0xff
    "11101100", --  402 - 0x192  :  236 - 0xec
    "11111010", --  403 - 0x193  :  250 - 0xfa
    "11111010", --  404 - 0x194  :  250 - 0xfa
    "11111010", --  405 - 0x195  :  250 - 0xfa
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11101010", --  409 - 0x199  :  234 - 0xea
    "11111010", --  410 - 0x19a  :  250 - 0xfa
    "11111010", --  411 - 0x19b  :  250 - 0xfa
    "11111010", --  412 - 0x19c  :  250 - 0xfa
    "11111010", --  413 - 0x19d  :  250 - 0xfa
    "11111010", --  414 - 0x19e  :  250 - 0xfa
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111100", --  417 - 0x1a1  :  252 - 0xfc
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111111", --  419 - 0x1a3  :  255 - 0xff
    "11111111", --  420 - 0x1a4  :  255 - 0xff
    "11111111", --  421 - 0x1a5  :  255 - 0xff
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111010", --  424 - 0x1a8  :  250 - 0xfa
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11111100", --  427 - 0x1ab  :  252 - 0xfc
    "11111111", --  428 - 0x1ac  :  255 - 0xff
    "11111111", --  429 - 0x1ad  :  255 - 0xff
    "11111111", --  430 - 0x1ae  :  255 - 0xff
    "11111111", --  431 - 0x1af  :  255 - 0xff
    "11111111", --  432 - 0x1b0  :  255 - 0xff
    "11111111", --  433 - 0x1b1  :  255 - 0xff
    "11110101", --  434 - 0x1b2  :  245 - 0xf5
    "11111011", --  435 - 0x1b3  :  251 - 0xfb
    "11111011", --  436 - 0x1b4  :  251 - 0xfb
    "11111011", --  437 - 0x1b5  :  251 - 0xfb
    "11111011", --  438 - 0x1b6  :  251 - 0xfb
    "11111011", --  439 - 0x1b7  :  251 - 0xfb
    "11111011", --  440 - 0x1b8  :  251 - 0xfb
    "11111011", --  441 - 0x1b9  :  251 - 0xfb
    "11111011", --  442 - 0x1ba  :  251 - 0xfb
    "11111011", --  443 - 0x1bb  :  251 - 0xfb
    "11111011", --  444 - 0x1bc  :  251 - 0xfb
    "11111011", --  445 - 0x1bd  :  251 - 0xfb
    "11101000", --  446 - 0x1be  :  232 - 0xe8
    "11101001", --  447 - 0x1bf  :  233 - 0xe9
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111100", --  449 - 0x1c1  :  252 - 0xfc
    "11111111", --  450 - 0x1c2  :  255 - 0xff
    "11111110", --  451 - 0x1c3  :  254 - 0xfe
    "11111110", --  452 - 0x1c4  :  254 - 0xfe
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11101100", --  454 - 0x1c6  :  236 - 0xec
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111010", --  456 - 0x1c8  :  250 - 0xfa
    "11111001", --  457 - 0x1c9  :  249 - 0xf9
    "11111010", --  458 - 0x1ca  :  250 - 0xfa
    "11111100", --  459 - 0x1cb  :  252 - 0xfc
    "11111111", --  460 - 0x1cc  :  255 - 0xff
    "11111111", --  461 - 0x1cd  :  255 - 0xff
    "11111111", --  462 - 0x1ce  :  255 - 0xff
    "11111110", --  463 - 0x1cf  :  254 - 0xfe
    "11111111", --  464 - 0x1d0  :  255 - 0xff
    "11111111", --  465 - 0x1d1  :  255 - 0xff
    "11111111", --  466 - 0x1d2  :  255 - 0xff
    "11111111", --  467 - 0x1d3  :  255 - 0xff
    "11111111", --  468 - 0x1d4  :  255 - 0xff
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "11111111", --  470 - 0x1d6  :  255 - 0xff
    "11101111", --  471 - 0x1d7  :  239 - 0xef
    "11111111", --  472 - 0x1d8  :  255 - 0xff
    "11111111", --  473 - 0x1d9  :  255 - 0xff
    "11111111", --  474 - 0x1da  :  255 - 0xff
    "11111111", --  475 - 0x1db  :  255 - 0xff
    "11111111", --  476 - 0x1dc  :  255 - 0xff
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11101100", --  478 - 0x1de  :  236 - 0xec
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11101010", --  480 - 0x1e0  :  234 - 0xea -- line 0xf
    "11111100", --  481 - 0x1e1  :  252 - 0xfc
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11101100", --  486 - 0x1e6  :  236 - 0xec
    "11111010", --  487 - 0x1e7  :  250 - 0xfa
    "11111010", --  488 - 0x1e8  :  250 - 0xfa
    "11111010", --  489 - 0x1e9  :  250 - 0xfa
    "11111010", --  490 - 0x1ea  :  250 - 0xfa
    "11111100", --  491 - 0x1eb  :  252 - 0xfc
    "11111111", --  492 - 0x1ec  :  255 - 0xff
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "11111111", --  494 - 0x1ee  :  255 - 0xff
    "11111111", --  495 - 0x1ef  :  255 - 0xff
    "11111111", --  496 - 0x1f0  :  255 - 0xff
    "11111101", --  497 - 0x1f1  :  253 - 0xfd
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111101", --  499 - 0x1f3  :  253 - 0xfd
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111101", --  501 - 0x1f5  :  253 - 0xfd
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11101111", --  503 - 0x1f7  :  239 - 0xef
    "11111111", --  504 - 0x1f8  :  255 - 0xff
    "11111101", --  505 - 0x1f9  :  253 - 0xfd
    "11111111", --  506 - 0x1fa  :  255 - 0xff
    "11111111", --  507 - 0x1fb  :  255 - 0xff
    "11111111", --  508 - 0x1fc  :  255 - 0xff
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "11101100", --  510 - 0x1fe  :  236 - 0xec
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111100", --  513 - 0x201  :  252 - 0xfc
    "11111111", --  514 - 0x202  :  255 - 0xff
    "11111110", --  515 - 0x203  :  254 - 0xfe
    "11111110", --  516 - 0x204  :  254 - 0xfe
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11101100", --  518 - 0x206  :  236 - 0xec
    "11101001", --  519 - 0x207  :  233 - 0xe9
    "11111010", --  520 - 0x208  :  250 - 0xfa
    "11111010", --  521 - 0x209  :  250 - 0xfa
    "11111010", --  522 - 0x20a  :  250 - 0xfa
    "11110111", --  523 - 0x20b  :  247 - 0xf7
    "11101011", --  524 - 0x20c  :  235 - 0xeb
    "11100110", --  525 - 0x20d  :  230 - 0xe6
    "11111111", --  526 - 0x20e  :  255 - 0xff
    "11111111", --  527 - 0x20f  :  255 - 0xff
    "11111111", --  528 - 0x210  :  255 - 0xff
    "11111101", --  529 - 0x211  :  253 - 0xfd
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11111101", --  531 - 0x213  :  253 - 0xfd
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111101", --  533 - 0x215  :  253 - 0xfd
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11101111", --  535 - 0x217  :  239 - 0xef
    "11111111", --  536 - 0x218  :  255 - 0xff
    "11111101", --  537 - 0x219  :  253 - 0xfd
    "11111111", --  538 - 0x21a  :  255 - 0xff
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11101100", --  542 - 0x21e  :  236 - 0xec
    "11101010", --  543 - 0x21f  :  234 - 0xea
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111100", --  545 - 0x221  :  252 - 0xfc
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111111", --  547 - 0x223  :  255 - 0xff
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11101100", --  550 - 0x226  :  236 - 0xec
    "11111010", --  551 - 0x227  :  250 - 0xfa
    "11111010", --  552 - 0x228  :  250 - 0xfa
    "11111010", --  553 - 0x229  :  250 - 0xfa
    "11101010", --  554 - 0x22a  :  234 - 0xea
    "11111010", --  555 - 0x22b  :  250 - 0xfa
    "11111010", --  556 - 0x22c  :  250 - 0xfa
    "11111100", --  557 - 0x22d  :  252 - 0xfc
    "11111111", --  558 - 0x22e  :  255 - 0xff
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "11111111", --  560 - 0x230  :  255 - 0xff
    "11111111", --  561 - 0x231  :  255 - 0xff
    "11111111", --  562 - 0x232  :  255 - 0xff
    "11111111", --  563 - 0x233  :  255 - 0xff
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "11101111", --  567 - 0x237  :  239 - 0xef
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111111", --  570 - 0x23a  :  255 - 0xff
    "11111110", --  571 - 0x23b  :  254 - 0xfe
    "11111110", --  572 - 0x23c  :  254 - 0xfe
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111100", --  577 - 0x241  :  252 - 0xfc
    "11111111", --  578 - 0x242  :  255 - 0xff
    "11111110", --  579 - 0x243  :  254 - 0xfe
    "11111110", --  580 - 0x244  :  254 - 0xfe
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11101100", --  582 - 0x246  :  236 - 0xec
    "11111001", --  583 - 0x247  :  249 - 0xf9
    "11111010", --  584 - 0x248  :  250 - 0xfa
    "11111010", --  585 - 0x249  :  250 - 0xfa
    "11111010", --  586 - 0x24a  :  250 - 0xfa
    "11111010", --  587 - 0x24b  :  250 - 0xfa
    "11101010", --  588 - 0x24c  :  234 - 0xea
    "11110111", --  589 - 0x24d  :  247 - 0xf7
    "11101011", --  590 - 0x24e  :  235 - 0xeb
    "11101011", --  591 - 0x24f  :  235 - 0xeb
    "11101011", --  592 - 0x250  :  235 - 0xeb
    "11101011", --  593 - 0x251  :  235 - 0xeb
    "11101011", --  594 - 0x252  :  235 - 0xeb
    "11101011", --  595 - 0x253  :  235 - 0xeb
    "11101011", --  596 - 0x254  :  235 - 0xeb
    "11101011", --  597 - 0x255  :  235 - 0xeb
    "11101011", --  598 - 0x256  :  235 - 0xeb
    "11101011", --  599 - 0x257  :  235 - 0xeb
    "11101011", --  600 - 0x258  :  235 - 0xeb
    "11100110", --  601 - 0x259  :  230 - 0xe6
    "11111111", --  602 - 0x25a  :  255 - 0xff
    "11111111", --  603 - 0x25b  :  255 - 0xff
    "11111111", --  604 - 0x25c  :  255 - 0xff
    "11111111", --  605 - 0x25d  :  255 - 0xff
    "11101100", --  606 - 0x25e  :  236 - 0xec
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111001", --  608 - 0x260  :  249 - 0xf9 -- line 0x13
    "11111100", --  609 - 0x261  :  252 - 0xfc
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11110101", --  614 - 0x266  :  245 - 0xf5
    "11111011", --  615 - 0x267  :  251 - 0xfb
    "11111011", --  616 - 0x268  :  251 - 0xfb
    "11111011", --  617 - 0x269  :  251 - 0xfb
    "11111011", --  618 - 0x26a  :  251 - 0xfb
    "11111011", --  619 - 0x26b  :  251 - 0xfb
    "11111011", --  620 - 0x26c  :  251 - 0xfb
    "11111011", --  621 - 0x26d  :  251 - 0xfb
    "11111011", --  622 - 0x26e  :  251 - 0xfb
    "11111011", --  623 - 0x26f  :  251 - 0xfb
    "11111011", --  624 - 0x270  :  251 - 0xfb
    "11111011", --  625 - 0x271  :  251 - 0xfb
    "11101000", --  626 - 0x272  :  232 - 0xe8
    "11111010", --  627 - 0x273  :  250 - 0xfa
    "11111010", --  628 - 0x274  :  250 - 0xfa
    "11101010", --  629 - 0x275  :  234 - 0xea
    "11111010", --  630 - 0x276  :  250 - 0xfa
    "11111010", --  631 - 0x277  :  250 - 0xfa
    "11101001", --  632 - 0x278  :  233 - 0xe9
    "11111100", --  633 - 0x279  :  252 - 0xfc
    "11111111", --  634 - 0x27a  :  255 - 0xff
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "11111110", --  636 - 0x27c  :  254 - 0xfe
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11101100", --  638 - 0x27e  :  236 - 0xec
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111100", --  641 - 0x281  :  252 - 0xfc
    "11111111", --  642 - 0x282  :  255 - 0xff
    "11111110", --  643 - 0x283  :  254 - 0xfe
    "11111110", --  644 - 0x284  :  254 - 0xfe
    "11111111", --  645 - 0x285  :  255 - 0xff
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111101", --  647 - 0x287  :  253 - 0xfd
    "11111111", --  648 - 0x288  :  255 - 0xff
    "11111101", --  649 - 0x289  :  253 - 0xfd
    "11111111", --  650 - 0x28a  :  255 - 0xff
    "11111101", --  651 - 0x28b  :  253 - 0xfd
    "11111111", --  652 - 0x28c  :  255 - 0xff
    "11111101", --  653 - 0x28d  :  253 - 0xfd
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111101", --  655 - 0x28f  :  253 - 0xfd
    "11111111", --  656 - 0x290  :  255 - 0xff
    "11111111", --  657 - 0x291  :  255 - 0xff
    "11101100", --  658 - 0x292  :  236 - 0xec
    "11101001", --  659 - 0x293  :  233 - 0xe9
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "11111010", --  661 - 0x295  :  250 - 0xfa
    "11101010", --  662 - 0x296  :  234 - 0xea
    "11111010", --  663 - 0x297  :  250 - 0xfa
    "11111010", --  664 - 0x298  :  250 - 0xfa
    "11111100", --  665 - 0x299  :  252 - 0xfc
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111111", --  668 - 0x29c  :  255 - 0xff
    "11111111", --  669 - 0x29d  :  255 - 0xff
    "11101100", --  670 - 0x29e  :  236 - 0xec
    "11101010", --  671 - 0x29f  :  234 - 0xea
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111100", --  673 - 0x2a1  :  252 - 0xfc
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111101", --  679 - 0x2a7  :  253 - 0xfd
    "11111111", --  680 - 0x2a8  :  255 - 0xff
    "11111101", --  681 - 0x2a9  :  253 - 0xfd
    "11111111", --  682 - 0x2aa  :  255 - 0xff
    "11111101", --  683 - 0x2ab  :  253 - 0xfd
    "11111111", --  684 - 0x2ac  :  255 - 0xff
    "11111101", --  685 - 0x2ad  :  253 - 0xfd
    "11111111", --  686 - 0x2ae  :  255 - 0xff
    "11111101", --  687 - 0x2af  :  253 - 0xfd
    "11111111", --  688 - 0x2b0  :  255 - 0xff
    "11111111", --  689 - 0x2b1  :  255 - 0xff
    "11101100", --  690 - 0x2b2  :  236 - 0xec
    "11100111", --  691 - 0x2b3  :  231 - 0xe7
    "11111011", --  692 - 0x2b4  :  251 - 0xfb
    "11111011", --  693 - 0x2b5  :  251 - 0xfb
    "11111011", --  694 - 0x2b6  :  251 - 0xfb
    "11111011", --  695 - 0x2b7  :  251 - 0xfb
    "11111011", --  696 - 0x2b8  :  251 - 0xfb
    "11110110", --  697 - 0x2b9  :  246 - 0xf6
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111110", --  699 - 0x2bb  :  254 - 0xfe
    "11111110", --  700 - 0x2bc  :  254 - 0xfe
    "11111111", --  701 - 0x2bd  :  255 - 0xff
    "11101100", --  702 - 0x2be  :  236 - 0xec
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111100", --  705 - 0x2c1  :  252 - 0xfc
    "11111111", --  706 - 0x2c2  :  255 - 0xff
    "11111110", --  707 - 0x2c3  :  254 - 0xfe
    "11111110", --  708 - 0x2c4  :  254 - 0xfe
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11100101", --  710 - 0x2c6  :  229 - 0xe5
    "11101011", --  711 - 0x2c7  :  235 - 0xeb
    "11101011", --  712 - 0x2c8  :  235 - 0xeb
    "11101011", --  713 - 0x2c9  :  235 - 0xeb
    "11101011", --  714 - 0x2ca  :  235 - 0xeb
    "11101011", --  715 - 0x2cb  :  235 - 0xeb
    "11101011", --  716 - 0x2cc  :  235 - 0xeb
    "11101011", --  717 - 0x2cd  :  235 - 0xeb
    "11101011", --  718 - 0x2ce  :  235 - 0xeb
    "11100110", --  719 - 0x2cf  :  230 - 0xe6
    "11111111", --  720 - 0x2d0  :  255 - 0xff
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11101100", --  722 - 0x2d2  :  236 - 0xec
    "11111100", --  723 - 0x2d3  :  252 - 0xfc
    "11111111", --  724 - 0x2d4  :  255 - 0xff
    "11111111", --  725 - 0x2d5  :  255 - 0xff
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "11111111", --  728 - 0x2d8  :  255 - 0xff
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11101100", --  734 - 0x2de  :  236 - 0xec
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa -- line 0x17
    "11111100", --  737 - 0x2e1  :  252 - 0xfc
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11110101", --  742 - 0x2e6  :  245 - 0xf5
    "11111011", --  743 - 0x2e7  :  251 - 0xfb
    "11111011", --  744 - 0x2e8  :  251 - 0xfb
    "11111011", --  745 - 0x2e9  :  251 - 0xfb
    "11111011", --  746 - 0x2ea  :  251 - 0xfb
    "11111011", --  747 - 0x2eb  :  251 - 0xfb
    "11111011", --  748 - 0x2ec  :  251 - 0xfb
    "11111011", --  749 - 0x2ed  :  251 - 0xfb
    "11111011", --  750 - 0x2ee  :  251 - 0xfb
    "11110110", --  751 - 0x2ef  :  246 - 0xf6
    "11111111", --  752 - 0x2f0  :  255 - 0xff
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "11110101", --  754 - 0x2f2  :  245 - 0xf5
    "11110110", --  755 - 0x2f3  :  246 - 0xf6
    "11111111", --  756 - 0x2f4  :  255 - 0xff
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "11111111", --  760 - 0x2f8  :  255 - 0xff
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111110", --  763 - 0x2fb  :  254 - 0xfe
    "11111110", --  764 - 0x2fc  :  254 - 0xfe
    "11111111", --  765 - 0x2fd  :  255 - 0xff
    "11101100", --  766 - 0x2fe  :  236 - 0xec
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa -- line 0x18
    "11111100", --  769 - 0x301  :  252 - 0xfc
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111110", --  771 - 0x303  :  254 - 0xfe
    "11111110", --  772 - 0x304  :  254 - 0xfe
    "11111111", --  773 - 0x305  :  255 - 0xff
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111101", --  789 - 0x315  :  253 - 0xfd
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111101", --  791 - 0x317  :  253 - 0xfd
    "11111111", --  792 - 0x318  :  255 - 0xff
    "11111101", --  793 - 0x319  :  253 - 0xfd
    "11111111", --  794 - 0x31a  :  255 - 0xff
    "11111111", --  795 - 0x31b  :  255 - 0xff
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11101100", --  798 - 0x31e  :  236 - 0xec
    "11101001", --  799 - 0x31f  :  233 - 0xe9
    "11101010", --  800 - 0x320  :  234 - 0xea -- line 0x19
    "11111100", --  801 - 0x321  :  252 - 0xfc
    "11111111", --  802 - 0x322  :  255 - 0xff
    "11111111", --  803 - 0x323  :  255 - 0xff
    "11111111", --  804 - 0x324  :  255 - 0xff
    "11111111", --  805 - 0x325  :  255 - 0xff
    "11111111", --  806 - 0x326  :  255 - 0xff
    "11111101", --  807 - 0x327  :  253 - 0xfd
    "11111111", --  808 - 0x328  :  255 - 0xff
    "11111101", --  809 - 0x329  :  253 - 0xfd
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "11111101", --  811 - 0x32b  :  253 - 0xfd
    "11111111", --  812 - 0x32c  :  255 - 0xff
    "11111101", --  813 - 0x32d  :  253 - 0xfd
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111101", --  815 - 0x32f  :  253 - 0xfd
    "11111111", --  816 - 0x330  :  255 - 0xff
    "11111101", --  817 - 0x331  :  253 - 0xfd
    "11111111", --  818 - 0x332  :  255 - 0xff
    "11111101", --  819 - 0x333  :  253 - 0xfd
    "11111111", --  820 - 0x334  :  255 - 0xff
    "11111101", --  821 - 0x335  :  253 - 0xfd
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111101", --  823 - 0x337  :  253 - 0xfd
    "11111111", --  824 - 0x338  :  255 - 0xff
    "11111101", --  825 - 0x339  :  253 - 0xfd
    "11111111", --  826 - 0x33a  :  255 - 0xff
    "11111111", --  827 - 0x33b  :  255 - 0xff
    "11111111", --  828 - 0x33c  :  255 - 0xff
    "11111111", --  829 - 0x33d  :  255 - 0xff
    "11101100", --  830 - 0x33e  :  236 - 0xec
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11110111", --  833 - 0x341  :  247 - 0xf7
    "11101011", --  834 - 0x342  :  235 - 0xeb
    "11100110", --  835 - 0x343  :  230 - 0xe6
    "11111111", --  836 - 0x344  :  255 - 0xff
    "11111111", --  837 - 0x345  :  255 - 0xff
    "11111111", --  838 - 0x346  :  255 - 0xff
    "11111101", --  839 - 0x347  :  253 - 0xfd
    "11111111", --  840 - 0x348  :  255 - 0xff
    "11111101", --  841 - 0x349  :  253 - 0xfd
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111101", --  843 - 0x34b  :  253 - 0xfd
    "11111111", --  844 - 0x34c  :  255 - 0xff
    "11111101", --  845 - 0x34d  :  253 - 0xfd
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111101", --  847 - 0x34f  :  253 - 0xfd
    "11111111", --  848 - 0x350  :  255 - 0xff
    "11111101", --  849 - 0x351  :  253 - 0xfd
    "11111111", --  850 - 0x352  :  255 - 0xff
    "11111101", --  851 - 0x353  :  253 - 0xfd
    "11111111", --  852 - 0x354  :  255 - 0xff
    "11111111", --  853 - 0x355  :  255 - 0xff
    "11111111", --  854 - 0x356  :  255 - 0xff
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11111111", --  856 - 0x358  :  255 - 0xff
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "11100101", --  860 - 0x35c  :  229 - 0xe5
    "11101011", --  861 - 0x35d  :  235 - 0xeb
    "11111000", --  862 - 0x35e  :  248 - 0xf8
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "11111010", --  865 - 0x361  :  250 - 0xfa
    "11111010", --  866 - 0x362  :  250 - 0xfa
    "11111100", --  867 - 0x363  :  252 - 0xfc
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111111", --  870 - 0x366  :  255 - 0xff
    "11111111", --  871 - 0x367  :  255 - 0xff
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11111111", --  882 - 0x372  :  255 - 0xff
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11101100", --  892 - 0x37c  :  236 - 0xec
    "11111010", --  893 - 0x37d  :  250 - 0xfa
    "11111010", --  894 - 0x37e  :  250 - 0xfa
    "11111001", --  895 - 0x37f  :  249 - 0xf9
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111010", --  898 - 0x382  :  250 - 0xfa
    "11110111", --  899 - 0x383  :  247 - 0xf7
    "11101011", --  900 - 0x384  :  235 - 0xeb
    "11101011", --  901 - 0x385  :  235 - 0xeb
    "11101011", --  902 - 0x386  :  235 - 0xeb
    "11101011", --  903 - 0x387  :  235 - 0xeb
    "11101011", --  904 - 0x388  :  235 - 0xeb
    "11101011", --  905 - 0x389  :  235 - 0xeb
    "11101011", --  906 - 0x38a  :  235 - 0xeb
    "11101011", --  907 - 0x38b  :  235 - 0xeb
    "11101011", --  908 - 0x38c  :  235 - 0xeb
    "11101011", --  909 - 0x38d  :  235 - 0xeb
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11101011", --  922 - 0x39a  :  235 - 0xeb
    "11101011", --  923 - 0x39b  :  235 - 0xeb
    "11111000", --  924 - 0x39c  :  248 - 0xf8
    "11111010", --  925 - 0x39d  :  250 - 0xfa
    "11111010", --  926 - 0x39e  :  250 - 0xfa
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11101001", --  949 - 0x3b5  :  233 - 0xe9
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11101010", --  956 - 0x3bc  :  234 - 0xea
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "00000101", --  961 - 0x3c1  :    5 - 0x5
    "00000101", --  962 - 0x3c2  :    5 - 0x5
    "00000101", --  963 - 0x3c3  :    5 - 0x5
    "01010101", --  964 - 0x3c4  :   85 - 0x55
    "01010101", --  965 - 0x3c5  :   85 - 0x55
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "00010001", --  968 - 0x3c8  :   17 - 0x11
    "01000000", --  969 - 0x3c9  :   64 - 0x40
    "01010000", --  970 - 0x3ca  :   80 - 0x50
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "01010101", --  972 - 0x3cc  :   85 - 0x55
    "01010101", --  973 - 0x3cd  :   85 - 0x55
    "01010101", --  974 - 0x3ce  :   85 - 0x55
    "01010101", --  975 - 0x3cf  :   85 - 0x55
    "00010001", --  976 - 0x3d0  :   17 - 0x11
    "01000100", --  977 - 0x3d1  :   68 - 0x44
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "01010101", --  982 - 0x3d6  :   85 - 0x55
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "00010001", --  984 - 0x3d8  :   17 - 0x11
    "01000100", --  985 - 0x3d9  :   68 - 0x44
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000100", --  988 - 0x3dc  :    4 - 0x4
    "00000101", --  989 - 0x3dd  :    5 - 0x5
    "00000101", --  990 - 0x3de  :    5 - 0x5
    "01000101", --  991 - 0x3df  :   69 - 0x45
    "00010001", --  992 - 0x3e0  :   17 - 0x11
    "01000100", --  993 - 0x3e1  :   68 - 0x44
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010001", --  995 - 0x3e3  :   81 - 0x51
    "01010000", --  996 - 0x3e4  :   80 - 0x50
    "01010000", --  997 - 0x3e5  :   80 - 0x50
    "00010000", --  998 - 0x3e6  :   16 - 0x10
    "01000100", --  999 - 0x3e7  :   68 - 0x44
    "00010001", -- 1000 - 0x3e8  :   17 - 0x11
    "01000000", -- 1001 - 0x3e9  :   64 - 0x40
    "01010000", -- 1002 - 0x3ea  :   80 - 0x50
    "01010000", -- 1003 - 0x3eb  :   80 - 0x50
    "01000100", -- 1004 - 0x3ec  :   68 - 0x44
    "00000101", -- 1005 - 0x3ed  :    5 - 0x5
    "00000001", -- 1006 - 0x3ee  :    1 - 0x1
    "01000100", -- 1007 - 0x3ef  :   68 - 0x44
    "01010001", -- 1008 - 0x3f0  :   81 - 0x51
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "01010100", -- 1015 - 0x3f7  :   84 - 0x54
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
