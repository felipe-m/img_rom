//-   Sprites Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_LAWN_SPR_PLN1
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 1
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      11'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      11'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      11'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      11'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      11'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      11'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      11'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      11'hD: dout  = 8'b00000111; //   13 :   7 - 0x7
      11'hE: dout  = 8'b00000111; //   14 :   7 - 0x7
      11'hF: dout  = 8'b00000110; //   15 :   6 - 0x6
      11'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      11'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      11'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      11'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      11'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      11'h15: dout  = 8'b11111111; //   21 : 255 - 0xff
      11'h16: dout  = 8'b11111111; //   22 : 255 - 0xff
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      11'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      11'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      11'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      11'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      11'h1D: dout  = 8'b11100000; //   29 : 224 - 0xe0
      11'h1E: dout  = 8'b11100000; //   30 : 224 - 0xe0
      11'h1F: dout  = 8'b01100000; //   31 :  96 - 0x60
      11'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x4
      11'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      11'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      11'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      11'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      11'h25: dout  = 8'b00011111; //   37 :  31 - 0x1f
      11'h26: dout  = 8'b01111111; //   38 : 127 - 0x7f
      11'h27: dout  = 8'b11110000; //   39 : 240 - 0xf0
      11'h28: dout  = 8'b00000000; //   40 :   0 - 0x0 -- Sprite 0x5
      11'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      11'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      11'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      11'h2D: dout  = 8'b11111000; //   45 : 248 - 0xf8
      11'h2E: dout  = 8'b11111110; //   46 : 254 - 0xfe
      11'h2F: dout  = 8'b00001111; //   47 :  15 - 0xf
      11'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      11'h31: dout  = 8'b00000000; //   49 :   0 - 0x0
      11'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      11'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      11'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      11'h35: dout  = 8'b11100111; //   53 : 231 - 0xe7
      11'h36: dout  = 8'b11100111; //   54 : 231 - 0xe7
      11'h37: dout  = 8'b01100110; //   55 : 102 - 0x66
      11'h38: dout  = 8'b00000000; //   56 :   0 - 0x0 -- Sprite 0x7
      11'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      11'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      11'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      11'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout  = 8'b11000111; //   61 : 199 - 0xc7
      11'h3E: dout  = 8'b11000111; //   62 : 199 - 0xc7
      11'h3F: dout  = 8'b01100110; //   63 : 102 - 0x66
      11'h40: dout  = 8'b00000110; //   64 :   6 - 0x6 -- Sprite 0x8
      11'h41: dout  = 8'b00000110; //   65 :   6 - 0x6
      11'h42: dout  = 8'b00000110; //   66 :   6 - 0x6
      11'h43: dout  = 8'b00000110; //   67 :   6 - 0x6
      11'h44: dout  = 8'b00000110; //   68 :   6 - 0x6
      11'h45: dout  = 8'b00000110; //   69 :   6 - 0x6
      11'h46: dout  = 8'b00000110; //   70 :   6 - 0x6
      11'h47: dout  = 8'b00000110; //   71 :   6 - 0x6
      11'h48: dout  = 8'b11111111; //   72 : 255 - 0xff -- Sprite 0x9
      11'h49: dout  = 8'b11111111; //   73 : 255 - 0xff
      11'h4A: dout  = 8'b11111111; //   74 : 255 - 0xff
      11'h4B: dout  = 8'b11111111; //   75 : 255 - 0xff
      11'h4C: dout  = 8'b11111111; //   76 : 255 - 0xff
      11'h4D: dout  = 8'b11111111; //   77 : 255 - 0xff
      11'h4E: dout  = 8'b11111111; //   78 : 255 - 0xff
      11'h4F: dout  = 8'b11111111; //   79 : 255 - 0xff
      11'h50: dout  = 8'b01100000; //   80 :  96 - 0x60 -- Sprite 0xa
      11'h51: dout  = 8'b01100000; //   81 :  96 - 0x60
      11'h52: dout  = 8'b01100000; //   82 :  96 - 0x60
      11'h53: dout  = 8'b01100000; //   83 :  96 - 0x60
      11'h54: dout  = 8'b01100000; //   84 :  96 - 0x60
      11'h55: dout  = 8'b01100000; //   85 :  96 - 0x60
      11'h56: dout  = 8'b01100000; //   86 :  96 - 0x60
      11'h57: dout  = 8'b01100000; //   87 :  96 - 0x60
      11'h58: dout  = 8'b00000001; //   88 :   1 - 0x1 -- Sprite 0xb
      11'h59: dout  = 8'b00000011; //   89 :   3 - 0x3
      11'h5A: dout  = 8'b00000011; //   90 :   3 - 0x3
      11'h5B: dout  = 8'b00000111; //   91 :   7 - 0x7
      11'h5C: dout  = 8'b00000110; //   92 :   6 - 0x6
      11'h5D: dout  = 8'b00000110; //   93 :   6 - 0x6
      11'h5E: dout  = 8'b00000110; //   94 :   6 - 0x6
      11'h5F: dout  = 8'b00000110; //   95 :   6 - 0x6
      11'h60: dout  = 8'b11000111; //   96 : 199 - 0xc7 -- Sprite 0xc
      11'h61: dout  = 8'b10011111; //   97 : 159 - 0x9f
      11'h62: dout  = 8'b00111111; //   98 :  63 - 0x3f
      11'h63: dout  = 8'b01111111; //   99 : 127 - 0x7f
      11'h64: dout  = 8'b01111111; //  100 : 127 - 0x7f
      11'h65: dout  = 8'b11111111; //  101 : 255 - 0xff
      11'h66: dout  = 8'b11111111; //  102 : 255 - 0xff
      11'h67: dout  = 8'b11111111; //  103 : 255 - 0xff
      11'h68: dout  = 8'b11100011; //  104 : 227 - 0xe3 -- Sprite 0xd
      11'h69: dout  = 8'b11111001; //  105 : 249 - 0xf9
      11'h6A: dout  = 8'b11111100; //  106 : 252 - 0xfc
      11'h6B: dout  = 8'b11111110; //  107 : 254 - 0xfe
      11'h6C: dout  = 8'b11111110; //  108 : 254 - 0xfe
      11'h6D: dout  = 8'b11111111; //  109 : 255 - 0xff
      11'h6E: dout  = 8'b11111111; //  110 : 255 - 0xff
      11'h6F: dout  = 8'b11111111; //  111 : 255 - 0xff
      11'h70: dout  = 8'b10000110; //  112 : 134 - 0x86 -- Sprite 0xe
      11'h71: dout  = 8'b11000110; //  113 : 198 - 0xc6
      11'h72: dout  = 8'b11000110; //  114 : 198 - 0xc6
      11'h73: dout  = 8'b11100110; //  115 : 230 - 0xe6
      11'h74: dout  = 8'b01100110; //  116 : 102 - 0x66
      11'h75: dout  = 8'b01100110; //  117 : 102 - 0x66
      11'h76: dout  = 8'b01100110; //  118 : 102 - 0x66
      11'h77: dout  = 8'b01100110; //  119 : 102 - 0x66
      11'h78: dout  = 8'b01100110; //  120 : 102 - 0x66 -- Sprite 0xf
      11'h79: dout  = 8'b01100110; //  121 : 102 - 0x66
      11'h7A: dout  = 8'b01100110; //  122 : 102 - 0x66
      11'h7B: dout  = 8'b01100110; //  123 : 102 - 0x66
      11'h7C: dout  = 8'b01100110; //  124 : 102 - 0x66
      11'h7D: dout  = 8'b01100110; //  125 : 102 - 0x66
      11'h7E: dout  = 8'b01100110; //  126 : 102 - 0x66
      11'h7F: dout  = 8'b01100110; //  127 : 102 - 0x66
      11'h80: dout  = 8'b01100110; //  128 : 102 - 0x66 -- Sprite 0x10
      11'h81: dout  = 8'b00110110; //  129 :  54 - 0x36
      11'h82: dout  = 8'b10110110; //  130 : 182 - 0xb6
      11'h83: dout  = 8'b10011110; //  131 : 158 - 0x9e
      11'h84: dout  = 8'b11011110; //  132 : 222 - 0xde
      11'h85: dout  = 8'b11001110; //  133 : 206 - 0xce
      11'h86: dout  = 8'b11101110; //  134 : 238 - 0xee
      11'h87: dout  = 8'b11100110; //  135 : 230 - 0xe6
      11'h88: dout  = 8'b10000001; //  136 : 129 - 0x81 -- Sprite 0x11
      11'h89: dout  = 8'b00111100; //  137 :  60 - 0x3c
      11'h8A: dout  = 8'b01111110; //  138 : 126 - 0x7e
      11'h8B: dout  = 8'b01100110; //  139 : 102 - 0x66
      11'h8C: dout  = 8'b01100110; //  140 : 102 - 0x66
      11'h8D: dout  = 8'b01100110; //  141 : 102 - 0x66
      11'h8E: dout  = 8'b01100110; //  142 : 102 - 0x66
      11'h8F: dout  = 8'b01100110; //  143 : 102 - 0x66
      11'h90: dout  = 8'b11110110; //  144 : 246 - 0xf6 -- Sprite 0x12
      11'h91: dout  = 8'b11110010; //  145 : 242 - 0xf2
      11'h92: dout  = 8'b11111010; //  146 : 250 - 0xfa
      11'h93: dout  = 8'b11111000; //  147 : 248 - 0xf8
      11'h94: dout  = 8'b11111100; //  148 : 252 - 0xfc
      11'h95: dout  = 8'b11111100; //  149 : 252 - 0xfc
      11'h96: dout  = 8'b11111110; //  150 : 254 - 0xfe
      11'h97: dout  = 8'b11111110; //  151 : 254 - 0xfe
      11'h98: dout  = 8'b01100110; //  152 : 102 - 0x66 -- Sprite 0x13
      11'h99: dout  = 8'b01100110; //  153 : 102 - 0x66
      11'h9A: dout  = 8'b01100110; //  154 : 102 - 0x66
      11'h9B: dout  = 8'b01100110; //  155 : 102 - 0x66
      11'h9C: dout  = 8'b01100110; //  156 : 102 - 0x66
      11'h9D: dout  = 8'b01100110; //  157 : 102 - 0x66
      11'h9E: dout  = 8'b01100110; //  158 : 102 - 0x66
      11'h9F: dout  = 8'b01111110; //  159 : 126 - 0x7e
      11'hA0: dout  = 8'b11111111; //  160 : 255 - 0xff -- Sprite 0x14
      11'hA1: dout  = 8'b01111111; //  161 : 127 - 0x7f
      11'hA2: dout  = 8'b01111111; //  162 : 127 - 0x7f
      11'hA3: dout  = 8'b00111111; //  163 :  63 - 0x3f
      11'hA4: dout  = 8'b00111111; //  164 :  63 - 0x3f
      11'hA5: dout  = 8'b00011111; //  165 :  31 - 0x1f
      11'hA6: dout  = 8'b01011111; //  166 :  95 - 0x5f
      11'hA7: dout  = 8'b01001111; //  167 :  79 - 0x4f
      11'hA8: dout  = 8'b01100110; //  168 : 102 - 0x66 -- Sprite 0x15
      11'hA9: dout  = 8'b01100110; //  169 : 102 - 0x66
      11'hAA: dout  = 8'b01100110; //  170 : 102 - 0x66
      11'hAB: dout  = 8'b01100110; //  171 : 102 - 0x66
      11'hAC: dout  = 8'b01100110; //  172 : 102 - 0x66
      11'hAD: dout  = 8'b01111110; //  173 : 126 - 0x7e
      11'hAE: dout  = 8'b01111110; //  174 : 126 - 0x7e
      11'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout  = 8'b01111110; //  176 : 126 - 0x7e -- Sprite 0x16
      11'hB1: dout  = 8'b01100110; //  177 : 102 - 0x66
      11'hB2: dout  = 8'b01000010; //  178 :  66 - 0x42
      11'hB3: dout  = 8'b00011000; //  179 :  24 - 0x18
      11'hB4: dout  = 8'b00111100; //  180 :  60 - 0x3c
      11'hB5: dout  = 8'b01111110; //  181 : 126 - 0x7e
      11'hB6: dout  = 8'b11111111; //  182 : 255 - 0xff
      11'hB7: dout  = 8'b11111111; //  183 : 255 - 0xff
      11'hB8: dout  = 8'b01101111; //  184 : 111 - 0x6f -- Sprite 0x17
      11'hB9: dout  = 8'b01100111; //  185 : 103 - 0x67
      11'hBA: dout  = 8'b01110111; //  186 : 119 - 0x77
      11'hBB: dout  = 8'b01110011; //  187 : 115 - 0x73
      11'hBC: dout  = 8'b01111011; //  188 : 123 - 0x7b
      11'hBD: dout  = 8'b01111001; //  189 : 121 - 0x79
      11'hBE: dout  = 8'b01101101; //  190 : 109 - 0x6d
      11'hBF: dout  = 8'b01101100; //  191 : 108 - 0x6c
      11'hC0: dout  = 8'b01100000; //  192 :  96 - 0x60 -- Sprite 0x18
      11'hC1: dout  = 8'b01100000; //  193 :  96 - 0x60
      11'hC2: dout  = 8'b01100000; //  194 :  96 - 0x60
      11'hC3: dout  = 8'b01100000; //  195 :  96 - 0x60
      11'hC4: dout  = 8'b01100000; //  196 :  96 - 0x60
      11'hC5: dout  = 8'b01111111; //  197 : 127 - 0x7f
      11'hC6: dout  = 8'b01111111; //  198 : 127 - 0x7f
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b00000110; //  200 :   6 - 0x6 -- Sprite 0x19
      11'hC9: dout  = 8'b00000110; //  201 :   6 - 0x6
      11'hCA: dout  = 8'b00000110; //  202 :   6 - 0x6
      11'hCB: dout  = 8'b00000110; //  203 :   6 - 0x6
      11'hCC: dout  = 8'b00000110; //  204 :   6 - 0x6
      11'hCD: dout  = 8'b11100110; //  205 : 230 - 0xe6
      11'hCE: dout  = 8'b11100110; //  206 : 230 - 0xe6
      11'hCF: dout  = 8'b01100110; //  207 : 102 - 0x66
      11'hD0: dout  = 8'b11111111; //  208 : 255 - 0xff -- Sprite 0x1a
      11'hD1: dout  = 8'b11111111; //  209 : 255 - 0xff
      11'hD2: dout  = 8'b11111111; //  210 : 255 - 0xff
      11'hD3: dout  = 8'b11111111; //  211 : 255 - 0xff
      11'hD4: dout  = 8'b11100111; //  212 : 231 - 0xe7
      11'hD5: dout  = 8'b11000011; //  213 : 195 - 0xc3
      11'hD6: dout  = 8'b10011001; //  214 : 153 - 0x99
      11'hD7: dout  = 8'b00111100; //  215 :  60 - 0x3c
      11'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      11'hD9: dout  = 8'b01111110; //  217 : 126 - 0x7e
      11'hDA: dout  = 8'b01111110; //  218 : 126 - 0x7e
      11'hDB: dout  = 8'b01100110; //  219 : 102 - 0x66
      11'hDC: dout  = 8'b01100110; //  220 : 102 - 0x66
      11'hDD: dout  = 8'b01100110; //  221 : 102 - 0x66
      11'hDE: dout  = 8'b01100110; //  222 : 102 - 0x66
      11'hDF: dout  = 8'b01100110; //  223 : 102 - 0x66
      11'hE0: dout  = 8'b11111110; //  224 : 254 - 0xfe -- Sprite 0x1c
      11'hE1: dout  = 8'b11111100; //  225 : 252 - 0xfc
      11'hE2: dout  = 8'b11111001; //  226 : 249 - 0xf9
      11'hE3: dout  = 8'b11110011; //  227 : 243 - 0xf3
      11'hE4: dout  = 8'b11100111; //  228 : 231 - 0xe7
      11'hE5: dout  = 8'b11001110; //  229 : 206 - 0xce
      11'hE6: dout  = 8'b10011100; //  230 : 156 - 0x9c
      11'hE7: dout  = 8'b00111000; //  231 :  56 - 0x38
      11'hE8: dout  = 8'b01111110; //  232 : 126 - 0x7e -- Sprite 0x1d
      11'hE9: dout  = 8'b11100111; //  233 : 231 - 0xe7
      11'hEA: dout  = 8'b11000011; //  234 : 195 - 0xc3
      11'hEB: dout  = 8'b10000001; //  235 : 129 - 0x81
      11'hEC: dout  = 8'b00000000; //  236 :   0 - 0x0
      11'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      11'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b01111111; //  240 : 127 - 0x7f -- Sprite 0x1e
      11'hF1: dout  = 8'b00111111; //  241 :  63 - 0x3f
      11'hF2: dout  = 8'b10011111; //  242 : 159 - 0x9f
      11'hF3: dout  = 8'b11001111; //  243 : 207 - 0xcf
      11'hF4: dout  = 8'b11100111; //  244 : 231 - 0xe7
      11'hF5: dout  = 8'b01110011; //  245 : 115 - 0x73
      11'hF6: dout  = 8'b00111001; //  246 :  57 - 0x39
      11'hF7: dout  = 8'b00011100; //  247 :  28 - 0x1c
      11'hF8: dout  = 8'b00000110; //  248 :   6 - 0x6 -- Sprite 0x1f
      11'hF9: dout  = 8'b00000111; //  249 :   7 - 0x7
      11'hFA: dout  = 8'b00000111; //  250 :   7 - 0x7
      11'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      11'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      11'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      11'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      11'h101: dout  = 8'b11111111; //  257 : 255 - 0xff
      11'h102: dout  = 8'b11111111; //  258 : 255 - 0xff
      11'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b01100110; //  264 : 102 - 0x66 -- Sprite 0x21
      11'h109: dout  = 8'b11100111; //  265 : 231 - 0xe7
      11'h10A: dout  = 8'b11100111; //  266 : 231 - 0xe7
      11'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      11'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      11'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      11'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b01110000; //  272 : 112 - 0x70 -- Sprite 0x22
      11'h111: dout  = 8'b11100000; //  273 : 224 - 0xe0
      11'h112: dout  = 8'b11000000; //  274 : 192 - 0xc0
      11'h113: dout  = 8'b00000000; //  275 :   0 - 0x0
      11'h114: dout  = 8'b00000000; //  276 :   0 - 0x0
      11'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      11'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b00001110; //  280 :  14 - 0xe -- Sprite 0x23
      11'h119: dout  = 8'b00000111; //  281 :   7 - 0x7
      11'h11A: dout  = 8'b00000011; //  282 :   3 - 0x3
      11'h11B: dout  = 8'b00000000; //  283 :   0 - 0x0
      11'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      11'h11D: dout  = 8'b00000000; //  285 :   0 - 0x0
      11'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b01100000; //  288 :  96 - 0x60 -- Sprite 0x24
      11'h121: dout  = 8'b11100000; //  289 : 224 - 0xe0
      11'h122: dout  = 8'b11100000; //  290 : 224 - 0xe0
      11'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b00000000; //  296 :   0 - 0x0 -- Sprite 0x25
      11'h129: dout  = 8'b00000000; //  297 :   0 - 0x0
      11'h12A: dout  = 8'b00000000; //  298 :   0 - 0x0
      11'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      11'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      11'h12D: dout  = 8'b11000000; //  301 : 192 - 0xc0
      11'h12E: dout  = 8'b11100000; //  302 : 224 - 0xe0
      11'h12F: dout  = 8'b01110000; //  303 : 112 - 0x70
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      11'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      11'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout  = 8'b00000011; //  309 :   3 - 0x3
      11'h136: dout  = 8'b00000111; //  310 :   7 - 0x7
      11'h137: dout  = 8'b00001110; //  311 :  14 - 0xe
      11'h138: dout  = 8'b00111000; //  312 :  56 - 0x38 -- Sprite 0x27
      11'h139: dout  = 8'b10011100; //  313 : 156 - 0x9c
      11'h13A: dout  = 8'b11001110; //  314 : 206 - 0xce
      11'h13B: dout  = 8'b11100111; //  315 : 231 - 0xe7
      11'h13C: dout  = 8'b11110011; //  316 : 243 - 0xf3
      11'h13D: dout  = 8'b11111001; //  317 : 249 - 0xf9
      11'h13E: dout  = 8'b11111100; //  318 : 252 - 0xfc
      11'h13F: dout  = 8'b11111110; //  319 : 254 - 0xfe
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      11'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout  = 8'b10000001; //  324 : 129 - 0x81
      11'h145: dout  = 8'b11000011; //  325 : 195 - 0xc3
      11'h146: dout  = 8'b11100111; //  326 : 231 - 0xe7
      11'h147: dout  = 8'b01111110; //  327 : 126 - 0x7e
      11'h148: dout  = 8'b00011100; //  328 :  28 - 0x1c -- Sprite 0x29
      11'h149: dout  = 8'b00111001; //  329 :  57 - 0x39
      11'h14A: dout  = 8'b01110011; //  330 : 115 - 0x73
      11'h14B: dout  = 8'b11100111; //  331 : 231 - 0xe7
      11'h14C: dout  = 8'b11001111; //  332 : 207 - 0xcf
      11'h14D: dout  = 8'b10011111; //  333 : 159 - 0x9f
      11'h14E: dout  = 8'b00111111; //  334 :  63 - 0x3f
      11'h14F: dout  = 8'b01111111; //  335 : 127 - 0x7f
      11'h150: dout  = 8'b01100001; //  336 :  97 - 0x61 -- Sprite 0x2a
      11'h151: dout  = 8'b01100011; //  337 :  99 - 0x63
      11'h152: dout  = 8'b01100011; //  338 :  99 - 0x63
      11'h153: dout  = 8'b01100111; //  339 : 103 - 0x67
      11'h154: dout  = 8'b01100110; //  340 : 102 - 0x66
      11'h155: dout  = 8'b01100110; //  341 : 102 - 0x66
      11'h156: dout  = 8'b01100110; //  342 : 102 - 0x66
      11'h157: dout  = 8'b01100110; //  343 : 102 - 0x66
      11'h158: dout  = 8'b10000000; //  344 : 128 - 0x80 -- Sprite 0x2b
      11'h159: dout  = 8'b11000000; //  345 : 192 - 0xc0
      11'h15A: dout  = 8'b11000000; //  346 : 192 - 0xc0
      11'h15B: dout  = 8'b11100000; //  347 : 224 - 0xe0
      11'h15C: dout  = 8'b01100000; //  348 :  96 - 0x60
      11'h15D: dout  = 8'b01100000; //  349 :  96 - 0x60
      11'h15E: dout  = 8'b01100000; //  350 :  96 - 0x60
      11'h15F: dout  = 8'b01100000; //  351 :  96 - 0x60
      11'h160: dout  = 8'b00111100; //  352 :  60 - 0x3c -- Sprite 0x2c
      11'h161: dout  = 8'b10011001; //  353 : 153 - 0x99
      11'h162: dout  = 8'b11000011; //  354 : 195 - 0xc3
      11'h163: dout  = 8'b11100111; //  355 : 231 - 0xe7
      11'h164: dout  = 8'b11111111; //  356 : 255 - 0xff
      11'h165: dout  = 8'b11111111; //  357 : 255 - 0xff
      11'h166: dout  = 8'b11111111; //  358 : 255 - 0xff
      11'h167: dout  = 8'b11111111; //  359 : 255 - 0xff
      11'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      11'h169: dout  = 8'b01111111; //  361 : 127 - 0x7f
      11'h16A: dout  = 8'b01111111; //  362 : 127 - 0x7f
      11'h16B: dout  = 8'b01100000; //  363 :  96 - 0x60
      11'h16C: dout  = 8'b01100000; //  364 :  96 - 0x60
      11'h16D: dout  = 8'b01100000; //  365 :  96 - 0x60
      11'h16E: dout  = 8'b01100000; //  366 :  96 - 0x60
      11'h16F: dout  = 8'b01100000; //  367 :  96 - 0x60
      11'h170: dout  = 8'b01100110; //  368 : 102 - 0x66 -- Sprite 0x2e
      11'h171: dout  = 8'b11100110; //  369 : 230 - 0xe6
      11'h172: dout  = 8'b11100110; //  370 : 230 - 0xe6
      11'h173: dout  = 8'b00000110; //  371 :   6 - 0x6
      11'h174: dout  = 8'b00000110; //  372 :   6 - 0x6
      11'h175: dout  = 8'b00000110; //  373 :   6 - 0x6
      11'h176: dout  = 8'b00000110; //  374 :   6 - 0x6
      11'h177: dout  = 8'b00000110; //  375 :   6 - 0x6
      11'h178: dout  = 8'b00000001; //  376 :   1 - 0x1 -- Sprite 0x2f
      11'h179: dout  = 8'b01111100; //  377 : 124 - 0x7c
      11'h17A: dout  = 8'b01111110; //  378 : 126 - 0x7e
      11'h17B: dout  = 8'b01100110; //  379 : 102 - 0x66
      11'h17C: dout  = 8'b01100110; //  380 : 102 - 0x66
      11'h17D: dout  = 8'b01100110; //  381 : 102 - 0x66
      11'h17E: dout  = 8'b01100110; //  382 : 102 - 0x66
      11'h17F: dout  = 8'b01100110; //  383 : 102 - 0x66
      11'h180: dout  = 8'b11111111; //  384 : 255 - 0xff -- Sprite 0x30
      11'h181: dout  = 8'b11111111; //  385 : 255 - 0xff
      11'h182: dout  = 8'b01111110; //  386 : 126 - 0x7e
      11'h183: dout  = 8'b00111100; //  387 :  60 - 0x3c
      11'h184: dout  = 8'b00011000; //  388 :  24 - 0x18
      11'h185: dout  = 8'b01000010; //  389 :  66 - 0x42
      11'h186: dout  = 8'b01100110; //  390 : 102 - 0x66
      11'h187: dout  = 8'b01111110; //  391 : 126 - 0x7e
      11'h188: dout  = 8'b01100000; //  392 :  96 - 0x60 -- Sprite 0x31
      11'h189: dout  = 8'b01111111; //  393 : 127 - 0x7f
      11'h18A: dout  = 8'b01111111; //  394 : 127 - 0x7f
      11'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout  = 8'b11111111; //  396 : 255 - 0xff
      11'h18D: dout  = 8'b11111111; //  397 : 255 - 0xff
      11'h18E: dout  = 8'b11111111; //  398 : 255 - 0xff
      11'h18F: dout  = 8'b11111111; //  399 : 255 - 0xff
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout  = 8'b11111111; //  401 : 255 - 0xff
      11'h192: dout  = 8'b11111111; //  402 : 255 - 0xff
      11'h193: dout  = 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout  = 8'b11111111; //  404 : 255 - 0xff
      11'h195: dout  = 8'b11111111; //  405 : 255 - 0xff
      11'h196: dout  = 8'b11111111; //  406 : 255 - 0xff
      11'h197: dout  = 8'b11111111; //  407 : 255 - 0xff
      11'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      11'h199: dout  = 8'b11100000; //  409 : 224 - 0xe0
      11'h19A: dout  = 8'b11100000; //  410 : 224 - 0xe0
      11'h19B: dout  = 8'b01100000; //  411 :  96 - 0x60
      11'h19C: dout  = 8'b01100000; //  412 :  96 - 0x60
      11'h19D: dout  = 8'b01100000; //  413 :  96 - 0x60
      11'h19E: dout  = 8'b01100000; //  414 :  96 - 0x60
      11'h19F: dout  = 8'b01100000; //  415 :  96 - 0x60
      11'h1A0: dout  = 8'b01111110; //  416 : 126 - 0x7e -- Sprite 0x34
      11'h1A1: dout  = 8'b01100110; //  417 : 102 - 0x66
      11'h1A2: dout  = 8'b01100110; //  418 : 102 - 0x66
      11'h1A3: dout  = 8'b01100110; //  419 : 102 - 0x66
      11'h1A4: dout  = 8'b01100110; //  420 : 102 - 0x66
      11'h1A5: dout  = 8'b01100110; //  421 : 102 - 0x66
      11'h1A6: dout  = 8'b01100110; //  422 : 102 - 0x66
      11'h1A7: dout  = 8'b01100110; //  423 : 102 - 0x66
      11'h1A8: dout  = 8'b11111111; //  424 : 255 - 0xff -- Sprite 0x35
      11'h1A9: dout  = 8'b11111111; //  425 : 255 - 0xff
      11'h1AA: dout  = 8'b11111111; //  426 : 255 - 0xff
      11'h1AB: dout  = 8'b11111111; //  427 : 255 - 0xff
      11'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout  = 8'b01111111; //  429 : 127 - 0x7f
      11'h1AE: dout  = 8'b01111111; //  430 : 127 - 0x7f
      11'h1AF: dout  = 8'b01100000; //  431 :  96 - 0x60
      11'h1B0: dout  = 8'b11111111; //  432 : 255 - 0xff -- Sprite 0x36
      11'h1B1: dout  = 8'b11111111; //  433 : 255 - 0xff
      11'h1B2: dout  = 8'b11111111; //  434 : 255 - 0xff
      11'h1B3: dout  = 8'b11111111; //  435 : 255 - 0xff
      11'h1B4: dout  = 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout  = 8'b11111111; //  437 : 255 - 0xff
      11'h1B6: dout  = 8'b11111111; //  438 : 255 - 0xff
      11'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout  = 8'b01100000; //  440 :  96 - 0x60 -- Sprite 0x37
      11'h1B9: dout  = 8'b01100000; //  441 :  96 - 0x60
      11'h1BA: dout  = 8'b01100000; //  442 :  96 - 0x60
      11'h1BB: dout  = 8'b01100000; //  443 :  96 - 0x60
      11'h1BC: dout  = 8'b01100000; //  444 :  96 - 0x60
      11'h1BD: dout  = 8'b11100000; //  445 : 224 - 0xe0
      11'h1BE: dout  = 8'b11100000; //  446 : 224 - 0xe0
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b01100110; //  448 : 102 - 0x66 -- Sprite 0x38
      11'h1C1: dout  = 8'b01100110; //  449 : 102 - 0x66
      11'h1C2: dout  = 8'b01100110; //  450 : 102 - 0x66
      11'h1C3: dout  = 8'b01100110; //  451 : 102 - 0x66
      11'h1C4: dout  = 8'b01100110; //  452 : 102 - 0x66
      11'h1C5: dout  = 8'b01111110; //  453 : 126 - 0x7e
      11'h1C6: dout  = 8'b01111100; //  454 : 124 - 0x7c
      11'h1C7: dout  = 8'b00000001; //  455 :   1 - 0x1
      11'h1C8: dout  = 8'b11111111; //  456 : 255 - 0xff -- Sprite 0x39
      11'h1C9: dout  = 8'b11111111; //  457 : 255 - 0xff
      11'h1CA: dout  = 8'b11111111; //  458 : 255 - 0xff
      11'h1CB: dout  = 8'b11111111; //  459 : 255 - 0xff
      11'h1CC: dout  = 8'b11111111; //  460 : 255 - 0xff
      11'h1CD: dout  = 8'b11111111; //  461 : 255 - 0xff
      11'h1CE: dout  = 8'b11111111; //  462 : 255 - 0xff
      11'h1CF: dout  = 8'b11111110; //  463 : 254 - 0xfe
      11'h1D0: dout  = 8'b01100110; //  464 : 102 - 0x66 -- Sprite 0x3a
      11'h1D1: dout  = 8'b01100110; //  465 : 102 - 0x66
      11'h1D2: dout  = 8'b01100110; //  466 : 102 - 0x66
      11'h1D3: dout  = 8'b01100110; //  467 : 102 - 0x66
      11'h1D4: dout  = 8'b01100110; //  468 : 102 - 0x66
      11'h1D5: dout  = 8'b01111110; //  469 : 126 - 0x7e
      11'h1D6: dout  = 8'b00111100; //  470 :  60 - 0x3c
      11'h1D7: dout  = 8'b10000001; //  471 : 129 - 0x81
      11'h1D8: dout  = 8'b01100000; //  472 :  96 - 0x60 -- Sprite 0x3b
      11'h1D9: dout  = 8'b01100000; //  473 :  96 - 0x60
      11'h1DA: dout  = 8'b01100000; //  474 :  96 - 0x60
      11'h1DB: dout  = 8'b01100000; //  475 :  96 - 0x60
      11'h1DC: dout  = 8'b01100000; //  476 :  96 - 0x60
      11'h1DD: dout  = 8'b01111111; //  477 : 127 - 0x7f
      11'h1DE: dout  = 8'b01111111; //  478 : 127 - 0x7f
      11'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout  = 8'b11111111; //  485 : 255 - 0xff
      11'h1E6: dout  = 8'b11111111; //  486 : 255 - 0xff
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      11'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout  = 8'b11111111; //  493 : 255 - 0xff
      11'h1EE: dout  = 8'b11111111; //  494 : 255 - 0xff
      11'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout  = 8'b11111110; //  496 : 254 - 0xfe -- Sprite 0x3e
      11'h1F1: dout  = 8'b11111100; //  497 : 252 - 0xfc
      11'h1F2: dout  = 8'b11111001; //  498 : 249 - 0xf9
      11'h1F3: dout  = 8'b11110011; //  499 : 243 - 0xf3
      11'h1F4: dout  = 8'b11110011; //  500 : 243 - 0xf3
      11'h1F5: dout  = 8'b11111001; //  501 : 249 - 0xf9
      11'h1F6: dout  = 8'b11111100; //  502 : 252 - 0xfc
      11'h1F7: dout  = 8'b11111110; //  503 : 254 - 0xfe
      11'h1F8: dout  = 8'b11100000; //  504 : 224 - 0xe0 -- Sprite 0x3f
      11'h1F9: dout  = 8'b11000000; //  505 : 192 - 0xc0
      11'h1FA: dout  = 8'b11000000; //  506 : 192 - 0xc0
      11'h1FB: dout  = 8'b10000000; //  507 : 128 - 0x80
      11'h1FC: dout  = 8'b10000000; //  508 : 128 - 0x80
      11'h1FD: dout  = 8'b11000000; //  509 : 192 - 0xc0
      11'h1FE: dout  = 8'b11000000; //  510 : 192 - 0xc0
      11'h1FF: dout  = 8'b11100000; //  511 : 224 - 0xe0
      11'h200: dout  = 8'b01100110; //  512 : 102 - 0x66 -- Sprite 0x40
      11'h201: dout  = 8'b01100110; //  513 : 102 - 0x66
      11'h202: dout  = 8'b01100110; //  514 : 102 - 0x66
      11'h203: dout  = 8'b01100110; //  515 : 102 - 0x66
      11'h204: dout  = 8'b01100111; //  516 : 103 - 0x67
      11'h205: dout  = 8'b01100011; //  517 :  99 - 0x63
      11'h206: dout  = 8'b01100011; //  518 :  99 - 0x63
      11'h207: dout  = 8'b01100001; //  519 :  97 - 0x61
      11'h208: dout  = 8'b11111111; //  520 : 255 - 0xff -- Sprite 0x41
      11'h209: dout  = 8'b11111111; //  521 : 255 - 0xff
      11'h20A: dout  = 8'b11111111; //  522 : 255 - 0xff
      11'h20B: dout  = 8'b01111111; //  523 : 127 - 0x7f
      11'h20C: dout  = 8'b01111111; //  524 : 127 - 0x7f
      11'h20D: dout  = 8'b00111111; //  525 :  63 - 0x3f
      11'h20E: dout  = 8'b10011111; //  526 : 159 - 0x9f
      11'h20F: dout  = 8'b11000111; //  527 : 199 - 0xc7
      11'h210: dout  = 8'b11111111; //  528 : 255 - 0xff -- Sprite 0x42
      11'h211: dout  = 8'b11111111; //  529 : 255 - 0xff
      11'h212: dout  = 8'b11111111; //  530 : 255 - 0xff
      11'h213: dout  = 8'b11111110; //  531 : 254 - 0xfe
      11'h214: dout  = 8'b11111110; //  532 : 254 - 0xfe
      11'h215: dout  = 8'b11111100; //  533 : 252 - 0xfc
      11'h216: dout  = 8'b11111001; //  534 : 249 - 0xf9
      11'h217: dout  = 8'b11100011; //  535 : 227 - 0xe3
      11'h218: dout  = 8'b01100110; //  536 : 102 - 0x66 -- Sprite 0x43
      11'h219: dout  = 8'b01100110; //  537 : 102 - 0x66
      11'h21A: dout  = 8'b01100110; //  538 : 102 - 0x66
      11'h21B: dout  = 8'b01100110; //  539 : 102 - 0x66
      11'h21C: dout  = 8'b11100110; //  540 : 230 - 0xe6
      11'h21D: dout  = 8'b11000110; //  541 : 198 - 0xc6
      11'h21E: dout  = 8'b11000110; //  542 : 198 - 0xc6
      11'h21F: dout  = 8'b10000110; //  543 : 134 - 0x86
      11'h220: dout  = 8'b11111110; //  544 : 254 - 0xfe -- Sprite 0x44
      11'h221: dout  = 8'b11111111; //  545 : 255 - 0xff
      11'h222: dout  = 8'b11111111; //  546 : 255 - 0xff
      11'h223: dout  = 8'b11111111; //  547 : 255 - 0xff
      11'h224: dout  = 8'b11111111; //  548 : 255 - 0xff
      11'h225: dout  = 8'b11111111; //  549 : 255 - 0xff
      11'h226: dout  = 8'b11111111; //  550 : 255 - 0xff
      11'h227: dout  = 8'b11111111; //  551 : 255 - 0xff
      11'h228: dout  = 8'b01100000; //  552 :  96 - 0x60 -- Sprite 0x45
      11'h229: dout  = 8'b01100000; //  553 :  96 - 0x60
      11'h22A: dout  = 8'b01100000; //  554 :  96 - 0x60
      11'h22B: dout  = 8'b01100000; //  555 :  96 - 0x60
      11'h22C: dout  = 8'b01100000; //  556 :  96 - 0x60
      11'h22D: dout  = 8'b01100000; //  557 :  96 - 0x60
      11'h22E: dout  = 8'b01100000; //  558 :  96 - 0x60
      11'h22F: dout  = 8'b01100000; //  559 :  96 - 0x60
      11'h230: dout  = 8'b11110000; //  560 : 240 - 0xf0 -- Sprite 0x46
      11'h231: dout  = 8'b01111111; //  561 : 127 - 0x7f
      11'h232: dout  = 8'b00011111; //  562 :  31 - 0x1f
      11'h233: dout  = 8'b00000000; //  563 :   0 - 0x0
      11'h234: dout  = 8'b00000000; //  564 :   0 - 0x0
      11'h235: dout  = 8'b00000000; //  565 :   0 - 0x0
      11'h236: dout  = 8'b00000000; //  566 :   0 - 0x0
      11'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout  = 8'b00001111; //  568 :  15 - 0xf -- Sprite 0x47
      11'h239: dout  = 8'b11111110; //  569 : 254 - 0xfe
      11'h23A: dout  = 8'b11111000; //  570 : 248 - 0xf8
      11'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00000110; //  576 :   6 - 0x6 -- Sprite 0x48
      11'h241: dout  = 8'b00000111; //  577 :   7 - 0x7
      11'h242: dout  = 8'b00000111; //  578 :   7 - 0x7
      11'h243: dout  = 8'b00000000; //  579 :   0 - 0x0
      11'h244: dout  = 8'b00000000; //  580 :   0 - 0x0
      11'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      11'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b00000000; //  584 :   0 - 0x0 -- Sprite 0x49
      11'h249: dout  = 8'b00000000; //  585 :   0 - 0x0
      11'h24A: dout  = 8'b00000000; //  586 :   0 - 0x0
      11'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      11'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      11'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      11'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x4a
      11'h251: dout  = 8'b01110110; //  593 : 118 - 0x76
      11'h252: dout  = 8'b01010111; //  594 :  87 - 0x57
      11'h253: dout  = 8'b01010101; //  595 :  85 - 0x55
      11'h254: dout  = 8'b01010101; //  596 :  85 - 0x55
      11'h255: dout  = 8'b01110101; //  597 : 117 - 0x75
      11'h256: dout  = 8'b01000111; //  598 :  71 - 0x47
      11'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout  = 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      11'h259: dout  = 8'b01110111; //  601 : 119 - 0x77
      11'h25A: dout  = 8'b00010101; //  602 :  21 - 0x15
      11'h25B: dout  = 8'b01110101; //  603 : 117 - 0x75
      11'h25C: dout  = 8'b01000101; //  604 :  69 - 0x45
      11'h25D: dout  = 8'b01000101; //  605 :  69 - 0x45
      11'h25E: dout  = 8'b01110111; //  606 : 119 - 0x77
      11'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      11'h261: dout  = 8'b00100100; //  609 :  36 - 0x24
      11'h262: dout  = 8'b01101100; //  610 : 108 - 0x6c
      11'h263: dout  = 8'b00100100; //  611 :  36 - 0x24
      11'h264: dout  = 8'b00100100; //  612 :  36 - 0x24
      11'h265: dout  = 8'b00100100; //  613 :  36 - 0x24
      11'h266: dout  = 8'b00100101; //  614 :  37 - 0x25
      11'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      11'h268: dout  = 8'b00000000; //  616 :   0 - 0x0 -- Sprite 0x4d
      11'h269: dout  = 8'b01110100; //  617 : 116 - 0x74
      11'h26A: dout  = 8'b01000111; //  618 :  71 - 0x47
      11'h26B: dout  = 8'b01110101; //  619 : 117 - 0x75
      11'h26C: dout  = 8'b00010101; //  620 :  21 - 0x15
      11'h26D: dout  = 8'b00010101; //  621 :  21 - 0x15
      11'h26E: dout  = 8'b01110101; //  622 : 117 - 0x75
      11'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      11'h271: dout  = 8'b01000000; //  625 :  64 - 0x40
      11'h272: dout  = 8'b00011101; //  626 :  29 - 0x1d
      11'h273: dout  = 8'b01010101; //  627 :  85 - 0x55
      11'h274: dout  = 8'b01010001; //  628 :  81 - 0x51
      11'h275: dout  = 8'b01010001; //  629 :  81 - 0x51
      11'h276: dout  = 8'b01010001; //  630 :  81 - 0x51
      11'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      11'h278: dout  = 8'b00000000; //  632 :   0 - 0x0 -- Sprite 0x4f
      11'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      11'h27A: dout  = 8'b01001000; //  634 :  72 - 0x48
      11'h27B: dout  = 8'b01000001; //  635 :  65 - 0x41
      11'h27C: dout  = 8'b01000100; //  636 :  68 - 0x44
      11'h27D: dout  = 8'b01000000; //  637 :  64 - 0x40
      11'h27E: dout  = 8'b11010000; //  638 : 208 - 0xd0
      11'h27F: dout  = 8'b00000010; //  639 :   2 - 0x2
      11'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      11'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      11'h282: dout  = 8'b11111100; //  642 : 252 - 0xfc
      11'h283: dout  = 8'b11111110; //  643 : 254 - 0xfe
      11'h284: dout  = 8'b11101110; //  644 : 238 - 0xee
      11'h285: dout  = 8'b11101110; //  645 : 238 - 0xee
      11'h286: dout  = 8'b11101110; //  646 : 238 - 0xee
      11'h287: dout  = 8'b11101110; //  647 : 238 - 0xee
      11'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      11'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      11'h28A: dout  = 8'b11111100; //  650 : 252 - 0xfc
      11'h28B: dout  = 8'b11111110; //  651 : 254 - 0xfe
      11'h28C: dout  = 8'b11101110; //  652 : 238 - 0xee
      11'h28D: dout  = 8'b11101110; //  653 : 238 - 0xee
      11'h28E: dout  = 8'b11101110; //  654 : 238 - 0xee
      11'h28F: dout  = 8'b11101110; //  655 : 238 - 0xee
      11'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      11'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      11'h292: dout  = 8'b11111110; //  658 : 254 - 0xfe
      11'h293: dout  = 8'b11111110; //  659 : 254 - 0xfe
      11'h294: dout  = 8'b11100000; //  660 : 224 - 0xe0
      11'h295: dout  = 8'b11100000; //  661 : 224 - 0xe0
      11'h296: dout  = 8'b11111000; //  662 : 248 - 0xf8
      11'h297: dout  = 8'b11111000; //  663 : 248 - 0xf8
      11'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      11'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      11'h29A: dout  = 8'b01111100; //  666 : 124 - 0x7c
      11'h29B: dout  = 8'b11111110; //  667 : 254 - 0xfe
      11'h29C: dout  = 8'b11101110; //  668 : 238 - 0xee
      11'h29D: dout  = 8'b11100000; //  669 : 224 - 0xe0
      11'h29E: dout  = 8'b11111100; //  670 : 252 - 0xfc
      11'h29F: dout  = 8'b01111110; //  671 : 126 - 0x7e
      11'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x54
      11'h2A1: dout  = 8'b00000000; //  673 :   0 - 0x0
      11'h2A2: dout  = 8'b11111110; //  674 : 254 - 0xfe
      11'h2A3: dout  = 8'b11111110; //  675 : 254 - 0xfe
      11'h2A4: dout  = 8'b00111000; //  676 :  56 - 0x38
      11'h2A5: dout  = 8'b00111000; //  677 :  56 - 0x38
      11'h2A6: dout  = 8'b00111000; //  678 :  56 - 0x38
      11'h2A7: dout  = 8'b00111000; //  679 :  56 - 0x38
      11'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      11'h2AA: dout  = 8'b01111100; //  682 : 124 - 0x7c
      11'h2AB: dout  = 8'b11111110; //  683 : 254 - 0xfe
      11'h2AC: dout  = 8'b11101110; //  684 : 238 - 0xee
      11'h2AD: dout  = 8'b11101110; //  685 : 238 - 0xee
      11'h2AE: dout  = 8'b11101110; //  686 : 238 - 0xee
      11'h2AF: dout  = 8'b11101110; //  687 : 238 - 0xee
      11'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x56
      11'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      11'h2B2: dout  = 8'b11100000; //  690 : 224 - 0xe0
      11'h2B3: dout  = 8'b11100000; //  691 : 224 - 0xe0
      11'h2B4: dout  = 8'b11100000; //  692 : 224 - 0xe0
      11'h2B5: dout  = 8'b11100000; //  693 : 224 - 0xe0
      11'h2B6: dout  = 8'b11100000; //  694 : 224 - 0xe0
      11'h2B7: dout  = 8'b11100000; //  695 : 224 - 0xe0
      11'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      11'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      11'h2BA: dout  = 8'b11101110; //  698 : 238 - 0xee
      11'h2BB: dout  = 8'b11101110; //  699 : 238 - 0xee
      11'h2BC: dout  = 8'b11101110; //  700 : 238 - 0xee
      11'h2BD: dout  = 8'b11101110; //  701 : 238 - 0xee
      11'h2BE: dout  = 8'b11101110; //  702 : 238 - 0xee
      11'h2BF: dout  = 8'b11101110; //  703 : 238 - 0xee
      11'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x58
      11'h2C1: dout  = 8'b00000000; //  705 :   0 - 0x0
      11'h2C2: dout  = 8'b10001110; //  706 : 142 - 0x8e
      11'h2C3: dout  = 8'b11001110; //  707 : 206 - 0xce
      11'h2C4: dout  = 8'b11101110; //  708 : 238 - 0xee
      11'h2C5: dout  = 8'b11111110; //  709 : 254 - 0xfe
      11'h2C6: dout  = 8'b11111110; //  710 : 254 - 0xfe
      11'h2C7: dout  = 8'b11101110; //  711 : 238 - 0xee
      11'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0 -- Sprite 0x59
      11'h2C9: dout  = 8'b00000000; //  713 :   0 - 0x0
      11'h2CA: dout  = 8'b11111100; //  714 : 252 - 0xfc
      11'h2CB: dout  = 8'b11111110; //  715 : 254 - 0xfe
      11'h2CC: dout  = 8'b11101110; //  716 : 238 - 0xee
      11'h2CD: dout  = 8'b11101110; //  717 : 238 - 0xee
      11'h2CE: dout  = 8'b11101110; //  718 : 238 - 0xee
      11'h2CF: dout  = 8'b11101110; //  719 : 238 - 0xee
      11'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      11'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      11'h2D2: dout  = 8'b01111100; //  722 : 124 - 0x7c
      11'h2D3: dout  = 8'b11111110; //  723 : 254 - 0xfe
      11'h2D4: dout  = 8'b11101110; //  724 : 238 - 0xee
      11'h2D5: dout  = 8'b11101110; //  725 : 238 - 0xee
      11'h2D6: dout  = 8'b11101110; //  726 : 238 - 0xee
      11'h2D7: dout  = 8'b11101110; //  727 : 238 - 0xee
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b11111110; //  730 : 254 - 0xfe
      11'h2DB: dout  = 8'b11111110; //  731 : 254 - 0xfe
      11'h2DC: dout  = 8'b11100000; //  732 : 224 - 0xe0
      11'h2DD: dout  = 8'b11100000; //  733 : 224 - 0xe0
      11'h2DE: dout  = 8'b11111000; //  734 : 248 - 0xf8
      11'h2DF: dout  = 8'b11111000; //  735 : 248 - 0xf8
      11'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      11'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      11'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      11'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      11'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      11'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      11'h2E6: dout  = 8'b11001100; //  742 : 204 - 0xcc
      11'h2E7: dout  = 8'b11001100; //  743 : 204 - 0xcc
      11'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      11'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      11'h2EA: dout  = 8'b11111110; //  746 : 254 - 0xfe
      11'h2EB: dout  = 8'b11111110; //  747 : 254 - 0xfe
      11'h2EC: dout  = 8'b11100000; //  748 : 224 - 0xe0
      11'h2ED: dout  = 8'b11100000; //  749 : 224 - 0xe0
      11'h2EE: dout  = 8'b11111000; //  750 : 248 - 0xf8
      11'h2EF: dout  = 8'b11111000; //  751 : 248 - 0xf8
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      11'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      11'h2F2: dout  = 8'b11101110; //  754 : 238 - 0xee
      11'h2F3: dout  = 8'b11101110; //  755 : 238 - 0xee
      11'h2F4: dout  = 8'b11101110; //  756 : 238 - 0xee
      11'h2F5: dout  = 8'b11101110; //  757 : 238 - 0xee
      11'h2F6: dout  = 8'b11101110; //  758 : 238 - 0xee
      11'h2F7: dout  = 8'b11101110; //  759 : 238 - 0xee
      11'h2F8: dout  = 8'b01111110; //  760 : 126 - 0x7e -- Sprite 0x5f
      11'h2F9: dout  = 8'b01111110; //  761 : 126 - 0x7e
      11'h2FA: dout  = 8'b01111110; //  762 : 126 - 0x7e
      11'h2FB: dout  = 8'b01111110; //  763 : 126 - 0x7e
      11'h2FC: dout  = 8'b01111110; //  764 : 126 - 0x7e
      11'h2FD: dout  = 8'b01111110; //  765 : 126 - 0x7e
      11'h2FE: dout  = 8'b01111110; //  766 : 126 - 0x7e
      11'h2FF: dout  = 8'b01111110; //  767 : 126 - 0x7e
      11'h300: dout  = 8'b11101110; //  768 : 238 - 0xee -- Sprite 0x60
      11'h301: dout  = 8'b11101110; //  769 : 238 - 0xee
      11'h302: dout  = 8'b11111110; //  770 : 254 - 0xfe
      11'h303: dout  = 8'b11111100; //  771 : 252 - 0xfc
      11'h304: dout  = 8'b11100000; //  772 : 224 - 0xe0
      11'h305: dout  = 8'b11100000; //  773 : 224 - 0xe0
      11'h306: dout  = 8'b00000000; //  774 :   0 - 0x0
      11'h307: dout  = 8'b00000000; //  775 :   0 - 0x0
      11'h308: dout  = 8'b11101110; //  776 : 238 - 0xee -- Sprite 0x61
      11'h309: dout  = 8'b11101110; //  777 : 238 - 0xee
      11'h30A: dout  = 8'b11111100; //  778 : 252 - 0xfc
      11'h30B: dout  = 8'b11111100; //  779 : 252 - 0xfc
      11'h30C: dout  = 8'b11101110; //  780 : 238 - 0xee
      11'h30D: dout  = 8'b11101110; //  781 : 238 - 0xee
      11'h30E: dout  = 8'b00000000; //  782 :   0 - 0x0
      11'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      11'h310: dout  = 8'b11100000; //  784 : 224 - 0xe0 -- Sprite 0x62
      11'h311: dout  = 8'b11100000; //  785 : 224 - 0xe0
      11'h312: dout  = 8'b11100000; //  786 : 224 - 0xe0
      11'h313: dout  = 8'b11100000; //  787 : 224 - 0xe0
      11'h314: dout  = 8'b11111110; //  788 : 254 - 0xfe
      11'h315: dout  = 8'b11111110; //  789 : 254 - 0xfe
      11'h316: dout  = 8'b00000000; //  790 :   0 - 0x0
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b00001110; //  792 :  14 - 0xe -- Sprite 0x63
      11'h319: dout  = 8'b00001110; //  793 :  14 - 0xe
      11'h31A: dout  = 8'b00001110; //  794 :  14 - 0xe
      11'h31B: dout  = 8'b11101110; //  795 : 238 - 0xee
      11'h31C: dout  = 8'b11111110; //  796 : 254 - 0xfe
      11'h31D: dout  = 8'b01111100; //  797 : 124 - 0x7c
      11'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      11'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout  = 8'b00111000; //  800 :  56 - 0x38 -- Sprite 0x64
      11'h321: dout  = 8'b00111000; //  801 :  56 - 0x38
      11'h322: dout  = 8'b00111000; //  802 :  56 - 0x38
      11'h323: dout  = 8'b00111000; //  803 :  56 - 0x38
      11'h324: dout  = 8'b00111000; //  804 :  56 - 0x38
      11'h325: dout  = 8'b00111000; //  805 :  56 - 0x38
      11'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      11'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      11'h328: dout  = 8'b11101110; //  808 : 238 - 0xee -- Sprite 0x65
      11'h329: dout  = 8'b11101110; //  809 : 238 - 0xee
      11'h32A: dout  = 8'b11111110; //  810 : 254 - 0xfe
      11'h32B: dout  = 8'b11111110; //  811 : 254 - 0xfe
      11'h32C: dout  = 8'b11101110; //  812 : 238 - 0xee
      11'h32D: dout  = 8'b11101110; //  813 : 238 - 0xee
      11'h32E: dout  = 8'b00000000; //  814 :   0 - 0x0
      11'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout  = 8'b11100000; //  816 : 224 - 0xe0 -- Sprite 0x66
      11'h331: dout  = 8'b11100000; //  817 : 224 - 0xe0
      11'h332: dout  = 8'b11100000; //  818 : 224 - 0xe0
      11'h333: dout  = 8'b11101110; //  819 : 238 - 0xee
      11'h334: dout  = 8'b11111110; //  820 : 254 - 0xfe
      11'h335: dout  = 8'b11111110; //  821 : 254 - 0xfe
      11'h336: dout  = 8'b00000000; //  822 :   0 - 0x0
      11'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      11'h338: dout  = 8'b11101110; //  824 : 238 - 0xee -- Sprite 0x67
      11'h339: dout  = 8'b11101110; //  825 : 238 - 0xee
      11'h33A: dout  = 8'b11111110; //  826 : 254 - 0xfe
      11'h33B: dout  = 8'b11111110; //  827 : 254 - 0xfe
      11'h33C: dout  = 8'b11101110; //  828 : 238 - 0xee
      11'h33D: dout  = 8'b11000110; //  829 : 198 - 0xc6
      11'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout  = 8'b11101110; //  832 : 238 - 0xee -- Sprite 0x68
      11'h341: dout  = 8'b11101110; //  833 : 238 - 0xee
      11'h342: dout  = 8'b11101110; //  834 : 238 - 0xee
      11'h343: dout  = 8'b11101110; //  835 : 238 - 0xee
      11'h344: dout  = 8'b11101110; //  836 : 238 - 0xee
      11'h345: dout  = 8'b11101110; //  837 : 238 - 0xee
      11'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout  = 8'b11101110; //  840 : 238 - 0xee -- Sprite 0x69
      11'h349: dout  = 8'b11101110; //  841 : 238 - 0xee
      11'h34A: dout  = 8'b11101110; //  842 : 238 - 0xee
      11'h34B: dout  = 8'b11101110; //  843 : 238 - 0xee
      11'h34C: dout  = 8'b11111110; //  844 : 254 - 0xfe
      11'h34D: dout  = 8'b11111100; //  845 : 252 - 0xfc
      11'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout  = 8'b11101110; //  848 : 238 - 0xee -- Sprite 0x6a
      11'h351: dout  = 8'b11101110; //  849 : 238 - 0xee
      11'h352: dout  = 8'b11101110; //  850 : 238 - 0xee
      11'h353: dout  = 8'b11101110; //  851 : 238 - 0xee
      11'h354: dout  = 8'b11111110; //  852 : 254 - 0xfe
      11'h355: dout  = 8'b01111100; //  853 : 124 - 0x7c
      11'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout  = 8'b11100000; //  856 : 224 - 0xe0 -- Sprite 0x6b
      11'h359: dout  = 8'b11100000; //  857 : 224 - 0xe0
      11'h35A: dout  = 8'b11100000; //  858 : 224 - 0xe0
      11'h35B: dout  = 8'b11100000; //  859 : 224 - 0xe0
      11'h35C: dout  = 8'b11111110; //  860 : 254 - 0xfe
      11'h35D: dout  = 8'b11111110; //  861 : 254 - 0xfe
      11'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout  = 8'b00011000; //  864 :  24 - 0x18 -- Sprite 0x6c
      11'h361: dout  = 8'b00011000; //  865 :  24 - 0x18
      11'h362: dout  = 8'b00110000; //  866 :  48 - 0x30
      11'h363: dout  = 8'b00110000; //  867 :  48 - 0x30
      11'h364: dout  = 8'b01100110; //  868 : 102 - 0x66
      11'h365: dout  = 8'b01100110; //  869 : 102 - 0x66
      11'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      11'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      11'h368: dout  = 8'b11100000; //  872 : 224 - 0xe0 -- Sprite 0x6d
      11'h369: dout  = 8'b11100000; //  873 : 224 - 0xe0
      11'h36A: dout  = 8'b11100000; //  874 : 224 - 0xe0
      11'h36B: dout  = 8'b11100000; //  875 : 224 - 0xe0
      11'h36C: dout  = 8'b11100000; //  876 : 224 - 0xe0
      11'h36D: dout  = 8'b11100000; //  877 : 224 - 0xe0
      11'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout  = 8'b11101110; //  880 : 238 - 0xee -- Sprite 0x6e
      11'h371: dout  = 8'b11101110; //  881 : 238 - 0xee
      11'h372: dout  = 8'b11101110; //  882 : 238 - 0xee
      11'h373: dout  = 8'b11101110; //  883 : 238 - 0xee
      11'h374: dout  = 8'b11111110; //  884 : 254 - 0xfe
      11'h375: dout  = 8'b01111100; //  885 : 124 - 0x7c
      11'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout  = 8'b01111110; //  888 : 126 - 0x7e -- Sprite 0x6f
      11'h379: dout  = 8'b01111110; //  889 : 126 - 0x7e
      11'h37A: dout  = 8'b01111110; //  890 : 126 - 0x7e
      11'h37B: dout  = 8'b01111110; //  891 : 126 - 0x7e
      11'h37C: dout  = 8'b00111100; //  892 :  60 - 0x3c
      11'h37D: dout  = 8'b00111100; //  893 :  60 - 0x3c
      11'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout  = 8'b00000111; //  896 :   7 - 0x7 -- Sprite 0x70
      11'h381: dout  = 8'b00011111; //  897 :  31 - 0x1f
      11'h382: dout  = 8'b00111111; //  898 :  63 - 0x3f
      11'h383: dout  = 8'b00111111; //  899 :  63 - 0x3f
      11'h384: dout  = 8'b01111111; //  900 : 127 - 0x7f
      11'h385: dout  = 8'b01111111; //  901 : 127 - 0x7f
      11'h386: dout  = 8'b01111111; //  902 : 127 - 0x7f
      11'h387: dout  = 8'b01111110; //  903 : 126 - 0x7e
      11'h388: dout  = 8'b11100000; //  904 : 224 - 0xe0 -- Sprite 0x71
      11'h389: dout  = 8'b11111000; //  905 : 248 - 0xf8
      11'h38A: dout  = 8'b11111100; //  906 : 252 - 0xfc
      11'h38B: dout  = 8'b11111100; //  907 : 252 - 0xfc
      11'h38C: dout  = 8'b11111110; //  908 : 254 - 0xfe
      11'h38D: dout  = 8'b11111110; //  909 : 254 - 0xfe
      11'h38E: dout  = 8'b11111110; //  910 : 254 - 0xfe
      11'h38F: dout  = 8'b01111110; //  911 : 126 - 0x7e
      11'h390: dout  = 8'b01111110; //  912 : 126 - 0x7e -- Sprite 0x72
      11'h391: dout  = 8'b01111110; //  913 : 126 - 0x7e
      11'h392: dout  = 8'b01111110; //  914 : 126 - 0x7e
      11'h393: dout  = 8'b01111110; //  915 : 126 - 0x7e
      11'h394: dout  = 8'b01111110; //  916 : 126 - 0x7e
      11'h395: dout  = 8'b01111110; //  917 : 126 - 0x7e
      11'h396: dout  = 8'b01111110; //  918 : 126 - 0x7e
      11'h397: dout  = 8'b01111110; //  919 : 126 - 0x7e
      11'h398: dout  = 8'b01111110; //  920 : 126 - 0x7e -- Sprite 0x73
      11'h399: dout  = 8'b01111111; //  921 : 127 - 0x7f
      11'h39A: dout  = 8'b01111111; //  922 : 127 - 0x7f
      11'h39B: dout  = 8'b01111111; //  923 : 127 - 0x7f
      11'h39C: dout  = 8'b00111111; //  924 :  63 - 0x3f
      11'h39D: dout  = 8'b00111111; //  925 :  63 - 0x3f
      11'h39E: dout  = 8'b00011111; //  926 :  31 - 0x1f
      11'h39F: dout  = 8'b00000111; //  927 :   7 - 0x7
      11'h3A0: dout  = 8'b01111110; //  928 : 126 - 0x7e -- Sprite 0x74
      11'h3A1: dout  = 8'b11111110; //  929 : 254 - 0xfe
      11'h3A2: dout  = 8'b11111110; //  930 : 254 - 0xfe
      11'h3A3: dout  = 8'b11111110; //  931 : 254 - 0xfe
      11'h3A4: dout  = 8'b11111100; //  932 : 252 - 0xfc
      11'h3A5: dout  = 8'b11111100; //  933 : 252 - 0xfc
      11'h3A6: dout  = 8'b11111000; //  934 : 248 - 0xf8
      11'h3A7: dout  = 8'b11100000; //  935 : 224 - 0xe0
      11'h3A8: dout  = 8'b01111111; //  936 : 127 - 0x7f -- Sprite 0x75
      11'h3A9: dout  = 8'b01111111; //  937 : 127 - 0x7f
      11'h3AA: dout  = 8'b01111111; //  938 : 127 - 0x7f
      11'h3AB: dout  = 8'b01111111; //  939 : 127 - 0x7f
      11'h3AC: dout  = 8'b01111111; //  940 : 127 - 0x7f
      11'h3AD: dout  = 8'b01111111; //  941 : 127 - 0x7f
      11'h3AE: dout  = 8'b00000111; //  942 :   7 - 0x7
      11'h3AF: dout  = 8'b00000111; //  943 :   7 - 0x7
      11'h3B0: dout  = 8'b11111110; //  944 : 254 - 0xfe -- Sprite 0x76
      11'h3B1: dout  = 8'b11111110; //  945 : 254 - 0xfe
      11'h3B2: dout  = 8'b11111110; //  946 : 254 - 0xfe
      11'h3B3: dout  = 8'b11111110; //  947 : 254 - 0xfe
      11'h3B4: dout  = 8'b11111110; //  948 : 254 - 0xfe
      11'h3B5: dout  = 8'b11111110; //  949 : 254 - 0xfe
      11'h3B6: dout  = 8'b11100000; //  950 : 224 - 0xe0
      11'h3B7: dout  = 8'b11100000; //  951 : 224 - 0xe0
      11'h3B8: dout  = 8'b00000111; //  952 :   7 - 0x7 -- Sprite 0x77
      11'h3B9: dout  = 8'b00000111; //  953 :   7 - 0x7
      11'h3BA: dout  = 8'b00000111; //  954 :   7 - 0x7
      11'h3BB: dout  = 8'b00000111; //  955 :   7 - 0x7
      11'h3BC: dout  = 8'b00000111; //  956 :   7 - 0x7
      11'h3BD: dout  = 8'b00000111; //  957 :   7 - 0x7
      11'h3BE: dout  = 8'b00000111; //  958 :   7 - 0x7
      11'h3BF: dout  = 8'b00000111; //  959 :   7 - 0x7
      11'h3C0: dout  = 8'b11100000; //  960 : 224 - 0xe0 -- Sprite 0x78
      11'h3C1: dout  = 8'b11100000; //  961 : 224 - 0xe0
      11'h3C2: dout  = 8'b11100000; //  962 : 224 - 0xe0
      11'h3C3: dout  = 8'b11100000; //  963 : 224 - 0xe0
      11'h3C4: dout  = 8'b11100000; //  964 : 224 - 0xe0
      11'h3C5: dout  = 8'b11100000; //  965 : 224 - 0xe0
      11'h3C6: dout  = 8'b11100000; //  966 : 224 - 0xe0
      11'h3C7: dout  = 8'b11100000; //  967 : 224 - 0xe0
      11'h3C8: dout  = 8'b01111111; //  968 : 127 - 0x7f -- Sprite 0x79
      11'h3C9: dout  = 8'b01111111; //  969 : 127 - 0x7f
      11'h3CA: dout  = 8'b01111111; //  970 : 127 - 0x7f
      11'h3CB: dout  = 8'b01111111; //  971 : 127 - 0x7f
      11'h3CC: dout  = 8'b01111111; //  972 : 127 - 0x7f
      11'h3CD: dout  = 8'b01111111; //  973 : 127 - 0x7f
      11'h3CE: dout  = 8'b01111110; //  974 : 126 - 0x7e
      11'h3CF: dout  = 8'b01111110; //  975 : 126 - 0x7e
      11'h3D0: dout  = 8'b11111110; //  976 : 254 - 0xfe -- Sprite 0x7a
      11'h3D1: dout  = 8'b11111110; //  977 : 254 - 0xfe
      11'h3D2: dout  = 8'b11111110; //  978 : 254 - 0xfe
      11'h3D3: dout  = 8'b11111110; //  979 : 254 - 0xfe
      11'h3D4: dout  = 8'b11111110; //  980 : 254 - 0xfe
      11'h3D5: dout  = 8'b11111110; //  981 : 254 - 0xfe
      11'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout  = 8'b01111110; //  984 : 126 - 0x7e -- Sprite 0x7b
      11'h3D9: dout  = 8'b01111111; //  985 : 127 - 0x7f
      11'h3DA: dout  = 8'b01111111; //  986 : 127 - 0x7f
      11'h3DB: dout  = 8'b01111111; //  987 : 127 - 0x7f
      11'h3DC: dout  = 8'b01111111; //  988 : 127 - 0x7f
      11'h3DD: dout  = 8'b01111111; //  989 : 127 - 0x7f
      11'h3DE: dout  = 8'b01111111; //  990 : 127 - 0x7f
      11'h3DF: dout  = 8'b01111110; //  991 : 126 - 0x7e
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      11'h3E1: dout  = 8'b11110000; //  993 : 240 - 0xf0
      11'h3E2: dout  = 8'b11110000; //  994 : 240 - 0xf0
      11'h3E3: dout  = 8'b11110000; //  995 : 240 - 0xf0
      11'h3E4: dout  = 8'b11110000; //  996 : 240 - 0xf0
      11'h3E5: dout  = 8'b11110000; //  997 : 240 - 0xf0
      11'h3E6: dout  = 8'b11110000; //  998 : 240 - 0xf0
      11'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      11'h3E8: dout  = 8'b01111110; // 1000 : 126 - 0x7e -- Sprite 0x7d
      11'h3E9: dout  = 8'b01111110; // 1001 : 126 - 0x7e
      11'h3EA: dout  = 8'b01111111; // 1002 : 127 - 0x7f
      11'h3EB: dout  = 8'b01111111; // 1003 : 127 - 0x7f
      11'h3EC: dout  = 8'b01111111; // 1004 : 127 - 0x7f
      11'h3ED: dout  = 8'b01111111; // 1005 : 127 - 0x7f
      11'h3EE: dout  = 8'b01111111; // 1006 : 127 - 0x7f
      11'h3EF: dout  = 8'b01111111; // 1007 : 127 - 0x7f
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b11111110; // 1010 : 254 - 0xfe
      11'h3F3: dout  = 8'b11111110; // 1011 : 254 - 0xfe
      11'h3F4: dout  = 8'b11111110; // 1012 : 254 - 0xfe
      11'h3F5: dout  = 8'b11111110; // 1013 : 254 - 0xfe
      11'h3F6: dout  = 8'b11111110; // 1014 : 254 - 0xfe
      11'h3F7: dout  = 8'b11111110; // 1015 : 254 - 0xfe
      11'h3F8: dout  = 8'b01111110; // 1016 : 126 - 0x7e -- Sprite 0x7f
      11'h3F9: dout  = 8'b11111110; // 1017 : 254 - 0xfe
      11'h3FA: dout  = 8'b11111110; // 1018 : 254 - 0xfe
      11'h3FB: dout  = 8'b11111110; // 1019 : 254 - 0xfe
      11'h3FC: dout  = 8'b11111110; // 1020 : 254 - 0xfe
      11'h3FD: dout  = 8'b11111110; // 1021 : 254 - 0xfe
      11'h3FE: dout  = 8'b11111110; // 1022 : 254 - 0xfe
      11'h3FF: dout  = 8'b01111110; // 1023 : 126 - 0x7e
      11'h400: dout  = 8'b01000000; // 1024 :  64 - 0x40 -- Sprite 0x80
      11'h401: dout  = 8'b00001000; // 1025 :   8 - 0x8
      11'h402: dout  = 8'b00000010; // 1026 :   2 - 0x2
      11'h403: dout  = 8'b00100000; // 1027 :  32 - 0x20
      11'h404: dout  = 8'b00000100; // 1028 :   4 - 0x4
      11'h405: dout  = 8'b01000000; // 1029 :  64 - 0x40
      11'h406: dout  = 8'b00000001; // 1030 :   1 - 0x1
      11'h407: dout  = 8'b00010000; // 1031 :  16 - 0x10
      11'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      11'h409: dout  = 8'b00010001; // 1033 :  17 - 0x11
      11'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      11'h40B: dout  = 8'b00100000; // 1035 :  32 - 0x20
      11'h40C: dout  = 8'b10001000; // 1036 : 136 - 0x88
      11'h40D: dout  = 8'b00000010; // 1037 :   2 - 0x2
      11'h40E: dout  = 8'b00100000; // 1038 :  32 - 0x20
      11'h40F: dout  = 8'b01000000; // 1039 :  64 - 0x40
      11'h410: dout  = 8'b00000001; // 1040 :   1 - 0x1 -- Sprite 0x82
      11'h411: dout  = 8'b00010000; // 1041 :  16 - 0x10
      11'h412: dout  = 8'b01000000; // 1042 :  64 - 0x40
      11'h413: dout  = 8'b00001000; // 1043 :   8 - 0x8
      11'h414: dout  = 8'b00000010; // 1044 :   2 - 0x2
      11'h415: dout  = 8'b00100000; // 1045 :  32 - 0x20
      11'h416: dout  = 8'b00000100; // 1046 :   4 - 0x4
      11'h417: dout  = 8'b01000000; // 1047 :  64 - 0x40
      11'h418: dout  = 8'b00010000; // 1048 :  16 - 0x10 -- Sprite 0x83
      11'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout  = 8'b01000100; // 1050 :  68 - 0x44
      11'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      11'h41C: dout  = 8'b00001000; // 1052 :   8 - 0x8
      11'h41D: dout  = 8'b00100010; // 1053 :  34 - 0x22
      11'h41E: dout  = 8'b10000000; // 1054 : 128 - 0x80
      11'h41F: dout  = 8'b00001000; // 1055 :   8 - 0x8
      11'h420: dout  = 8'b00010100; // 1056 :  20 - 0x14 -- Sprite 0x84
      11'h421: dout  = 8'b10110101; // 1057 : 181 - 0xb5
      11'h422: dout  = 8'b01000100; // 1058 :  68 - 0x44
      11'h423: dout  = 8'b01001010; // 1059 :  74 - 0x4a
      11'h424: dout  = 8'b10010010; // 1060 : 146 - 0x92
      11'h425: dout  = 8'b10010010; // 1061 : 146 - 0x92
      11'h426: dout  = 8'b01000100; // 1062 :  68 - 0x44
      11'h427: dout  = 8'b01001001; // 1063 :  73 - 0x49
      11'h428: dout  = 8'b01000010; // 1064 :  66 - 0x42 -- Sprite 0x85
      11'h429: dout  = 8'b01001010; // 1065 :  74 - 0x4a
      11'h42A: dout  = 8'b11001010; // 1066 : 202 - 0xca
      11'h42B: dout  = 8'b00101001; // 1067 :  41 - 0x29
      11'h42C: dout  = 8'b10100110; // 1068 : 166 - 0xa6
      11'h42D: dout  = 8'b10010010; // 1069 : 146 - 0x92
      11'h42E: dout  = 8'b10001001; // 1070 : 137 - 0x89
      11'h42F: dout  = 8'b00101101; // 1071 :  45 - 0x2d
      11'h430: dout  = 8'b10001000; // 1072 : 136 - 0x88 -- Sprite 0x86
      11'h431: dout  = 8'b00101001; // 1073 :  41 - 0x29
      11'h432: dout  = 8'b10000010; // 1074 : 130 - 0x82
      11'h433: dout  = 8'b10110110; // 1075 : 182 - 0xb6
      11'h434: dout  = 8'b10001000; // 1076 : 136 - 0x88
      11'h435: dout  = 8'b01001001; // 1077 :  73 - 0x49
      11'h436: dout  = 8'b01010010; // 1078 :  82 - 0x52
      11'h437: dout  = 8'b01010010; // 1079 :  82 - 0x52
      11'h438: dout  = 8'b10110010; // 1080 : 178 - 0xb2 -- Sprite 0x87
      11'h439: dout  = 8'b01001010; // 1081 :  74 - 0x4a
      11'h43A: dout  = 8'b10101001; // 1082 : 169 - 0xa9
      11'h43B: dout  = 8'b10100100; // 1083 : 164 - 0xa4
      11'h43C: dout  = 8'b01100010; // 1084 :  98 - 0x62
      11'h43D: dout  = 8'b01001011; // 1085 :  75 - 0x4b
      11'h43E: dout  = 8'b10010000; // 1086 : 144 - 0x90
      11'h43F: dout  = 8'b10010010; // 1087 : 146 - 0x92
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      11'h441: dout  = 8'b01100000; // 1089 :  96 - 0x60
      11'h442: dout  = 8'b11111110; // 1090 : 254 - 0xfe
      11'h443: dout  = 8'b11111111; // 1091 : 255 - 0xff
      11'h444: dout  = 8'b01111111; // 1092 : 127 - 0x7f
      11'h445: dout  = 8'b00011111; // 1093 :  31 - 0x1f
      11'h446: dout  = 8'b00001110; // 1094 :  14 - 0xe
      11'h447: dout  = 8'b00000000; // 1095 :   0 - 0x0
      11'h448: dout  = 8'b00110000; // 1096 :  48 - 0x30 -- Sprite 0x89
      11'h449: dout  = 8'b01111000; // 1097 : 120 - 0x78
      11'h44A: dout  = 8'b01111000; // 1098 : 120 - 0x78
      11'h44B: dout  = 8'b00111110; // 1099 :  62 - 0x3e
      11'h44C: dout  = 8'b00011111; // 1100 :  31 - 0x1f
      11'h44D: dout  = 8'b00011111; // 1101 :  31 - 0x1f
      11'h44E: dout  = 8'b00011111; // 1102 :  31 - 0x1f
      11'h44F: dout  = 8'b00001110; // 1103 :  14 - 0xe
      11'h450: dout  = 8'b01000000; // 1104 :  64 - 0x40 -- Sprite 0x8a
      11'h451: dout  = 8'b00001000; // 1105 :   8 - 0x8
      11'h452: dout  = 8'b00000010; // 1106 :   2 - 0x2
      11'h453: dout  = 8'b00101000; // 1107 :  40 - 0x28
      11'h454: dout  = 8'b00010100; // 1108 :  20 - 0x14
      11'h455: dout  = 8'b01010100; // 1109 :  84 - 0x54
      11'h456: dout  = 8'b00000001; // 1110 :   1 - 0x1
      11'h457: dout  = 8'b00010000; // 1111 :  16 - 0x10
      11'h458: dout  = 8'b01000000; // 1112 :  64 - 0x40 -- Sprite 0x8b
      11'h459: dout  = 8'b00000000; // 1113 :   0 - 0x0
      11'h45A: dout  = 8'b10010001; // 1114 : 145 - 0x91
      11'h45B: dout  = 8'b00010100; // 1115 :  20 - 0x14
      11'h45C: dout  = 8'b00101000; // 1116 :  40 - 0x28
      11'h45D: dout  = 8'b10001010; // 1117 : 138 - 0x8a
      11'h45E: dout  = 8'b01000000; // 1118 :  64 - 0x40
      11'h45F: dout  = 8'b00100000; // 1119 :  32 - 0x20
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      11'h461: dout  = 8'b00000111; // 1121 :   7 - 0x7
      11'h462: dout  = 8'b00011111; // 1122 :  31 - 0x1f
      11'h463: dout  = 8'b00111111; // 1123 :  63 - 0x3f
      11'h464: dout  = 8'b00111111; // 1124 :  63 - 0x3f
      11'h465: dout  = 8'b01111111; // 1125 : 127 - 0x7f
      11'h466: dout  = 8'b01111111; // 1126 : 127 - 0x7f
      11'h467: dout  = 8'b01111111; // 1127 : 127 - 0x7f
      11'h468: dout  = 8'b00000000; // 1128 :   0 - 0x0 -- Sprite 0x8d
      11'h469: dout  = 8'b11100000; // 1129 : 224 - 0xe0
      11'h46A: dout  = 8'b11111000; // 1130 : 248 - 0xf8
      11'h46B: dout  = 8'b11111000; // 1131 : 248 - 0xf8
      11'h46C: dout  = 8'b11110000; // 1132 : 240 - 0xf0
      11'h46D: dout  = 8'b11111000; // 1133 : 248 - 0xf8
      11'h46E: dout  = 8'b11110100; // 1134 : 244 - 0xf4
      11'h46F: dout  = 8'b11111000; // 1135 : 248 - 0xf8
      11'h470: dout  = 8'b01111111; // 1136 : 127 - 0x7f -- Sprite 0x8e
      11'h471: dout  = 8'b00111111; // 1137 :  63 - 0x3f
      11'h472: dout  = 8'b00111111; // 1138 :  63 - 0x3f
      11'h473: dout  = 8'b00011111; // 1139 :  31 - 0x1f
      11'h474: dout  = 8'b00011111; // 1140 :  31 - 0x1f
      11'h475: dout  = 8'b00001111; // 1141 :  15 - 0xf
      11'h476: dout  = 8'b00001111; // 1142 :  15 - 0xf
      11'h477: dout  = 8'b00000111; // 1143 :   7 - 0x7
      11'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe -- Sprite 0x8f
      11'h479: dout  = 8'b11111100; // 1145 : 252 - 0xfc
      11'h47A: dout  = 8'b11111100; // 1146 : 252 - 0xfc
      11'h47B: dout  = 8'b11111000; // 1147 : 248 - 0xf8
      11'h47C: dout  = 8'b11111000; // 1148 : 248 - 0xf8
      11'h47D: dout  = 8'b11110000; // 1149 : 240 - 0xf0
      11'h47E: dout  = 8'b11110000; // 1150 : 240 - 0xf0
      11'h47F: dout  = 8'b11100000; // 1151 : 224 - 0xe0
      11'h480: dout  = 8'b01000001; // 1152 :  65 - 0x41 -- Sprite 0x90
      11'h481: dout  = 8'b00001000; // 1153 :   8 - 0x8
      11'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout  = 8'b00100000; // 1155 :  32 - 0x20
      11'h484: dout  = 8'b00000100; // 1156 :   4 - 0x4
      11'h485: dout  = 8'b00000001; // 1157 :   1 - 0x1
      11'h486: dout  = 8'b01000000; // 1158 :  64 - 0x40
      11'h487: dout  = 8'b00001000; // 1159 :   8 - 0x8
      11'h488: dout  = 8'b00010001; // 1160 :  17 - 0x11 -- Sprite 0x91
      11'h489: dout  = 8'b00000000; // 1161 :   0 - 0x0
      11'h48A: dout  = 8'b10000100; // 1162 : 132 - 0x84
      11'h48B: dout  = 8'b00000010; // 1163 :   2 - 0x2
      11'h48C: dout  = 8'b00010000; // 1164 :  16 - 0x10
      11'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      11'h48E: dout  = 8'b01000010; // 1166 :  66 - 0x42
      11'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout  = 8'b00000100; // 1168 :   4 - 0x4 -- Sprite 0x92
      11'h491: dout  = 8'b01000000; // 1169 :  64 - 0x40
      11'h492: dout  = 8'b00010000; // 1170 :  16 - 0x10
      11'h493: dout  = 8'b00000010; // 1171 :   2 - 0x2
      11'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      11'h495: dout  = 8'b01000000; // 1173 :  64 - 0x40
      11'h496: dout  = 8'b00000100; // 1174 :   4 - 0x4
      11'h497: dout  = 8'b00100000; // 1175 :  32 - 0x20
      11'h498: dout  = 8'b01000010; // 1176 :  66 - 0x42 -- Sprite 0x93
      11'h499: dout  = 8'b00000000; // 1177 :   0 - 0x0
      11'h49A: dout  = 8'b10001000; // 1178 : 136 - 0x88
      11'h49B: dout  = 8'b00000001; // 1179 :   1 - 0x1
      11'h49C: dout  = 8'b00100000; // 1180 :  32 - 0x20
      11'h49D: dout  = 8'b00000100; // 1181 :   4 - 0x4
      11'h49E: dout  = 8'b00010000; // 1182 :  16 - 0x10
      11'h49F: dout  = 8'b10000000; // 1183 : 128 - 0x80
      11'h4A0: dout  = 8'b11001000; // 1184 : 200 - 0xc8 -- Sprite 0x94
      11'h4A1: dout  = 8'b00101010; // 1185 :  42 - 0x2a
      11'h4A2: dout  = 8'b10100010; // 1186 : 162 - 0xa2
      11'h4A3: dout  = 8'b10010100; // 1187 : 148 - 0x94
      11'h4A4: dout  = 8'b10010001; // 1188 : 145 - 0x91
      11'h4A5: dout  = 8'b01010101; // 1189 :  85 - 0x55
      11'h4A6: dout  = 8'b01000100; // 1190 :  68 - 0x44
      11'h4A7: dout  = 8'b00010010; // 1191 :  18 - 0x12
      11'h4A8: dout  = 8'b10101010; // 1192 : 170 - 0xaa -- Sprite 0x95
      11'h4A9: dout  = 8'b10100010; // 1193 : 162 - 0xa2
      11'h4AA: dout  = 8'b00010010; // 1194 :  18 - 0x12
      11'h4AB: dout  = 8'b01010011; // 1195 :  83 - 0x53
      11'h4AC: dout  = 8'b01001100; // 1196 :  76 - 0x4c
      11'h4AD: dout  = 8'b01010101; // 1197 :  85 - 0x55
      11'h4AE: dout  = 8'b10010001; // 1198 : 145 - 0x91
      11'h4AF: dout  = 8'b01001000; // 1199 :  72 - 0x48
      11'h4B0: dout  = 8'b01010001; // 1200 :  81 - 0x51 -- Sprite 0x96
      11'h4B1: dout  = 8'b00010101; // 1201 :  21 - 0x15
      11'h4B2: dout  = 8'b10100100; // 1202 : 164 - 0xa4
      11'h4B3: dout  = 8'b10001100; // 1203 : 140 - 0x8c
      11'h4B4: dout  = 8'b10101010; // 1204 : 170 - 0xaa
      11'h4B5: dout  = 8'b00100010; // 1205 :  34 - 0x22
      11'h4B6: dout  = 8'b10010000; // 1206 : 144 - 0x90
      11'h4B7: dout  = 8'b01000110; // 1207 :  70 - 0x46
      11'h4B8: dout  = 8'b00010011; // 1208 :  19 - 0x13 -- Sprite 0x97
      11'h4B9: dout  = 8'b01010101; // 1209 :  85 - 0x55
      11'h4BA: dout  = 8'b01100100; // 1210 : 100 - 0x64
      11'h4BB: dout  = 8'b00010010; // 1211 :  18 - 0x12
      11'h4BC: dout  = 8'b10101010; // 1212 : 170 - 0xaa
      11'h4BD: dout  = 8'b10101000; // 1213 : 168 - 0xa8
      11'h4BE: dout  = 8'b10000100; // 1214 : 132 - 0x84
      11'h4BF: dout  = 8'b11010100; // 1215 : 212 - 0xd4
      11'h4C0: dout  = 8'b00110000; // 1216 :  48 - 0x30 -- Sprite 0x98
      11'h4C1: dout  = 8'b01111000; // 1217 : 120 - 0x78
      11'h4C2: dout  = 8'b01111000; // 1218 : 120 - 0x78
      11'h4C3: dout  = 8'b00111110; // 1219 :  62 - 0x3e
      11'h4C4: dout  = 8'b00011111; // 1220 :  31 - 0x1f
      11'h4C5: dout  = 8'b00011111; // 1221 :  31 - 0x1f
      11'h4C6: dout  = 8'b00011111; // 1222 :  31 - 0x1f
      11'h4C7: dout  = 8'b00001110; // 1223 :  14 - 0xe
      11'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- Sprite 0x99
      11'h4C9: dout  = 8'b01100000; // 1225 :  96 - 0x60
      11'h4CA: dout  = 8'b11111110; // 1226 : 254 - 0xfe
      11'h4CB: dout  = 8'b11111111; // 1227 : 255 - 0xff
      11'h4CC: dout  = 8'b01111111; // 1228 : 127 - 0x7f
      11'h4CD: dout  = 8'b00011111; // 1229 :  31 - 0x1f
      11'h4CE: dout  = 8'b00001110; // 1230 :  14 - 0xe
      11'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout  = 8'b01000000; // 1232 :  64 - 0x40 -- Sprite 0x9a
      11'h4D1: dout  = 8'b00001100; // 1233 :  12 - 0xc
      11'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      11'h4D3: dout  = 8'b00101000; // 1235 :  40 - 0x28
      11'h4D4: dout  = 8'b00101100; // 1236 :  44 - 0x2c
      11'h4D5: dout  = 8'b00010001; // 1237 :  17 - 0x11
      11'h4D6: dout  = 8'b01000000; // 1238 :  64 - 0x40
      11'h4D7: dout  = 8'b00001000; // 1239 :   8 - 0x8
      11'h4D8: dout  = 8'b00100000; // 1240 :  32 - 0x20 -- Sprite 0x9b
      11'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      11'h4DA: dout  = 8'b10010100; // 1242 : 148 - 0x94
      11'h4DB: dout  = 8'b01001000; // 1243 :  72 - 0x48
      11'h4DC: dout  = 8'b00011000; // 1244 :  24 - 0x18
      11'h4DD: dout  = 8'b00000110; // 1245 :   6 - 0x6
      11'h4DE: dout  = 8'b01000000; // 1246 :  64 - 0x40
      11'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout  = 8'b01111111; // 1248 : 127 - 0x7f -- Sprite 0x9c
      11'h4E1: dout  = 8'b01111111; // 1249 : 127 - 0x7f
      11'h4E2: dout  = 8'b01111111; // 1250 : 127 - 0x7f
      11'h4E3: dout  = 8'b00111111; // 1251 :  63 - 0x3f
      11'h4E4: dout  = 8'b00110101; // 1252 :  53 - 0x35
      11'h4E5: dout  = 8'b00000010; // 1253 :   2 - 0x2
      11'h4E6: dout  = 8'b00000000; // 1254 :   0 - 0x0
      11'h4E7: dout  = 8'b00000000; // 1255 :   0 - 0x0
      11'h4E8: dout  = 8'b11110100; // 1256 : 244 - 0xf4 -- Sprite 0x9d
      11'h4E9: dout  = 8'b11111000; // 1257 : 248 - 0xf8
      11'h4EA: dout  = 8'b11110000; // 1258 : 240 - 0xf0
      11'h4EB: dout  = 8'b11101000; // 1259 : 232 - 0xe8
      11'h4EC: dout  = 8'b01010000; // 1260 :  80 - 0x50
      11'h4ED: dout  = 8'b10000000; // 1261 : 128 - 0x80
      11'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      11'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout  = 8'b11111110; // 1264 : 254 - 0xfe -- Sprite 0x9e
      11'h4F1: dout  = 8'b11111100; // 1265 : 252 - 0xfc
      11'h4F2: dout  = 8'b11111100; // 1266 : 252 - 0xfc
      11'h4F3: dout  = 8'b11111000; // 1267 : 248 - 0xf8
      11'h4F4: dout  = 8'b11111000; // 1268 : 248 - 0xf8
      11'h4F5: dout  = 8'b11111100; // 1269 : 252 - 0xfc
      11'h4F6: dout  = 8'b11111100; // 1270 : 252 - 0xfc
      11'h4F7: dout  = 8'b11111110; // 1271 : 254 - 0xfe
      11'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      11'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout  = 8'b01111110; // 1274 : 126 - 0x7e
      11'h4FB: dout  = 8'b01111110; // 1275 : 126 - 0x7e
      11'h4FC: dout  = 8'b01111110; // 1276 : 126 - 0x7e
      11'h4FD: dout  = 8'b01111110; // 1277 : 126 - 0x7e
      11'h4FE: dout  = 8'b01111110; // 1278 : 126 - 0x7e
      11'h4FF: dout  = 8'b01111110; // 1279 : 126 - 0x7e
      11'h500: dout  = 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0xa0
      11'h501: dout  = 8'b00111000; // 1281 :  56 - 0x38
      11'h502: dout  = 8'b01111100; // 1282 : 124 - 0x7c
      11'h503: dout  = 8'b11111000; // 1283 : 248 - 0xf8
      11'h504: dout  = 8'b01110000; // 1284 : 112 - 0x70
      11'h505: dout  = 8'b00100010; // 1285 :  34 - 0x22
      11'h506: dout  = 8'b00000101; // 1286 :   5 - 0x5
      11'h507: dout  = 8'b00000010; // 1287 :   2 - 0x2
      11'h508: dout  = 8'b00010000; // 1288 :  16 - 0x10 -- Sprite 0xa1
      11'h509: dout  = 8'b00111000; // 1289 :  56 - 0x38
      11'h50A: dout  = 8'b01111100; // 1290 : 124 - 0x7c
      11'h50B: dout  = 8'b11100000; // 1291 : 224 - 0xe0
      11'h50C: dout  = 8'b01100000; // 1292 :  96 - 0x60
      11'h50D: dout  = 8'b00100000; // 1293 :  32 - 0x20
      11'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      11'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      11'h510: dout  = 8'b00010000; // 1296 :  16 - 0x10 -- Sprite 0xa2
      11'h511: dout  = 8'b00111000; // 1297 :  56 - 0x38
      11'h512: dout  = 8'b01111100; // 1298 : 124 - 0x7c
      11'h513: dout  = 8'b00000000; // 1299 :   0 - 0x0
      11'h514: dout  = 8'b00000000; // 1300 :   0 - 0x0
      11'h515: dout  = 8'b00000000; // 1301 :   0 - 0x0
      11'h516: dout  = 8'b00000000; // 1302 :   0 - 0x0
      11'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- Sprite 0xa3
      11'h519: dout  = 8'b00100000; // 1305 :  32 - 0x20
      11'h51A: dout  = 8'b01100000; // 1306 :  96 - 0x60
      11'h51B: dout  = 8'b11100000; // 1307 : 224 - 0xe0
      11'h51C: dout  = 8'b01100000; // 1308 :  96 - 0x60
      11'h51D: dout  = 8'b00100000; // 1309 :  32 - 0x20
      11'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      11'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      11'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      11'h521: dout  = 8'b00100000; // 1313 :  32 - 0x20
      11'h522: dout  = 8'b01100011; // 1314 :  99 - 0x63
      11'h523: dout  = 8'b11100111; // 1315 : 231 - 0xe7
      11'h524: dout  = 8'b01100000; // 1316 :  96 - 0x60
      11'h525: dout  = 8'b00100010; // 1317 :  34 - 0x22
      11'h526: dout  = 8'b00000101; // 1318 :   5 - 0x5
      11'h527: dout  = 8'b00000010; // 1319 :   2 - 0x2
      11'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      11'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout  = 8'b11111111; // 1322 : 255 - 0xff
      11'h52B: dout  = 8'b11111111; // 1323 : 255 - 0xff
      11'h52C: dout  = 8'b00000000; // 1324 :   0 - 0x0
      11'h52D: dout  = 8'b00100010; // 1325 :  34 - 0x22
      11'h52E: dout  = 8'b00000101; // 1326 :   5 - 0x5
      11'h52F: dout  = 8'b00000010; // 1327 :   2 - 0x2
      11'h530: dout  = 8'b00010000; // 1328 :  16 - 0x10 -- Sprite 0xa6
      11'h531: dout  = 8'b00111000; // 1329 :  56 - 0x38
      11'h532: dout  = 8'b01111100; // 1330 : 124 - 0x7c
      11'h533: dout  = 8'b00000000; // 1331 :   0 - 0x0
      11'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      11'h535: dout  = 8'b00010010; // 1333 :  18 - 0x12
      11'h536: dout  = 8'b00110101; // 1334 :  53 - 0x35
      11'h537: dout  = 8'b00110010; // 1335 :  50 - 0x32
      11'h538: dout  = 8'b00110000; // 1336 :  48 - 0x30 -- Sprite 0xa7
      11'h539: dout  = 8'b00110000; // 1337 :  48 - 0x30
      11'h53A: dout  = 8'b00110100; // 1338 :  52 - 0x34
      11'h53B: dout  = 8'b00110000; // 1339 :  48 - 0x30
      11'h53C: dout  = 8'b00110000; // 1340 :  48 - 0x30
      11'h53D: dout  = 8'b00110010; // 1341 :  50 - 0x32
      11'h53E: dout  = 8'b00110101; // 1342 :  53 - 0x35
      11'h53F: dout  = 8'b00110010; // 1343 :  50 - 0x32
      11'h540: dout  = 8'b00110000; // 1344 :  48 - 0x30 -- Sprite 0xa8
      11'h541: dout  = 8'b00110000; // 1345 :  48 - 0x30
      11'h542: dout  = 8'b11110100; // 1346 : 244 - 0xf4
      11'h543: dout  = 8'b11110000; // 1347 : 240 - 0xf0
      11'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      11'h545: dout  = 8'b00100010; // 1349 :  34 - 0x22
      11'h546: dout  = 8'b00000101; // 1350 :   5 - 0x5
      11'h547: dout  = 8'b00000010; // 1351 :   2 - 0x2
      11'h548: dout  = 8'b00000000; // 1352 :   0 - 0x0 -- Sprite 0xa9
      11'h549: dout  = 8'b00000000; // 1353 :   0 - 0x0
      11'h54A: dout  = 8'b00000000; // 1354 :   0 - 0x0
      11'h54B: dout  = 8'b00000000; // 1355 :   0 - 0x0
      11'h54C: dout  = 8'b00000000; // 1356 :   0 - 0x0
      11'h54D: dout  = 8'b00000000; // 1357 :   0 - 0x0
      11'h54E: dout  = 8'b00000000; // 1358 :   0 - 0x0
      11'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      11'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      11'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout  = 8'b01010000; // 1362 :  80 - 0x50
      11'h553: dout  = 8'b10101000; // 1363 : 168 - 0xa8
      11'h554: dout  = 8'b01110000; // 1364 : 112 - 0x70
      11'h555: dout  = 8'b00100010; // 1365 :  34 - 0x22
      11'h556: dout  = 8'b00000101; // 1366 :   5 - 0x5
      11'h557: dout  = 8'b00000010; // 1367 :   2 - 0x2
      11'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      11'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout  = 8'b00000000; // 1374 :   0 - 0x0
      11'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout  = 8'b00000000; // 1380 :   0 - 0x0
      11'h565: dout  = 8'b00000000; // 1381 :   0 - 0x0
      11'h566: dout  = 8'b00000000; // 1382 :   0 - 0x0
      11'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      11'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      11'h569: dout  = 8'b00000000; // 1385 :   0 - 0x0
      11'h56A: dout  = 8'b11111111; // 1386 : 255 - 0xff
      11'h56B: dout  = 8'b00000000; // 1387 :   0 - 0x0
      11'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      11'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      11'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      11'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      11'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      11'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      11'h575: dout  = 8'b11111111; // 1397 : 255 - 0xff
      11'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      11'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      11'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      11'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      11'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      11'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      11'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      11'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      11'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      11'h581: dout  = 8'b00011111; // 1409 :  31 - 0x1f
      11'h582: dout  = 8'b00011111; // 1410 :  31 - 0x1f
      11'h583: dout  = 8'b00011111; // 1411 :  31 - 0x1f
      11'h584: dout  = 8'b00011111; // 1412 :  31 - 0x1f
      11'h585: dout  = 8'b00011111; // 1413 :  31 - 0x1f
      11'h586: dout  = 8'b00011111; // 1414 :  31 - 0x1f
      11'h587: dout  = 8'b00011111; // 1415 :  31 - 0x1f
      11'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0 -- Sprite 0xb1
      11'h589: dout  = 8'b11110000; // 1417 : 240 - 0xf0
      11'h58A: dout  = 8'b11110000; // 1418 : 240 - 0xf0
      11'h58B: dout  = 8'b11110000; // 1419 : 240 - 0xf0
      11'h58C: dout  = 8'b11110000; // 1420 : 240 - 0xf0
      11'h58D: dout  = 8'b11110000; // 1421 : 240 - 0xf0
      11'h58E: dout  = 8'b11110000; // 1422 : 240 - 0xf0
      11'h58F: dout  = 8'b11110000; // 1423 : 240 - 0xf0
      11'h590: dout  = 8'b00011111; // 1424 :  31 - 0x1f -- Sprite 0xb2
      11'h591: dout  = 8'b00011111; // 1425 :  31 - 0x1f
      11'h592: dout  = 8'b00011111; // 1426 :  31 - 0x1f
      11'h593: dout  = 8'b00011111; // 1427 :  31 - 0x1f
      11'h594: dout  = 8'b00000000; // 1428 :   0 - 0x0
      11'h595: dout  = 8'b00000000; // 1429 :   0 - 0x0
      11'h596: dout  = 8'b00000000; // 1430 :   0 - 0x0
      11'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout  = 8'b11110000; // 1432 : 240 - 0xf0 -- Sprite 0xb3
      11'h599: dout  = 8'b11110000; // 1433 : 240 - 0xf0
      11'h59A: dout  = 8'b11110000; // 1434 : 240 - 0xf0
      11'h59B: dout  = 8'b11110000; // 1435 : 240 - 0xf0
      11'h59C: dout  = 8'b00000000; // 1436 :   0 - 0x0
      11'h59D: dout  = 8'b00000000; // 1437 :   0 - 0x0
      11'h59E: dout  = 8'b00000000; // 1438 :   0 - 0x0
      11'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      11'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      11'h5A2: dout  = 8'b00111111; // 1442 :  63 - 0x3f
      11'h5A3: dout  = 8'b01111111; // 1443 : 127 - 0x7f
      11'h5A4: dout  = 8'b01111111; // 1444 : 127 - 0x7f
      11'h5A5: dout  = 8'b01111111; // 1445 : 127 - 0x7f
      11'h5A6: dout  = 8'b01111111; // 1446 : 127 - 0x7f
      11'h5A7: dout  = 8'b01111111; // 1447 : 127 - 0x7f
      11'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0 -- Sprite 0xb5
      11'h5A9: dout  = 8'b00000000; // 1449 :   0 - 0x0
      11'h5AA: dout  = 8'b11111000; // 1450 : 248 - 0xf8
      11'h5AB: dout  = 8'b11111000; // 1451 : 248 - 0xf8
      11'h5AC: dout  = 8'b11111000; // 1452 : 248 - 0xf8
      11'h5AD: dout  = 8'b11111000; // 1453 : 248 - 0xf8
      11'h5AE: dout  = 8'b11111000; // 1454 : 248 - 0xf8
      11'h5AF: dout  = 8'b11111000; // 1455 : 248 - 0xf8
      11'h5B0: dout  = 8'b01111111; // 1456 : 127 - 0x7f -- Sprite 0xb6
      11'h5B1: dout  = 8'b01111111; // 1457 : 127 - 0x7f
      11'h5B2: dout  = 8'b01111111; // 1458 : 127 - 0x7f
      11'h5B3: dout  = 8'b01000000; // 1459 :  64 - 0x40
      11'h5B4: dout  = 8'b00000000; // 1460 :   0 - 0x0
      11'h5B5: dout  = 8'b00000000; // 1461 :   0 - 0x0
      11'h5B6: dout  = 8'b00000000; // 1462 :   0 - 0x0
      11'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout  = 8'b11111000; // 1464 : 248 - 0xf8 -- Sprite 0xb7
      11'h5B9: dout  = 8'b11111000; // 1465 : 248 - 0xf8
      11'h5BA: dout  = 8'b11111000; // 1466 : 248 - 0xf8
      11'h5BB: dout  = 8'b00000000; // 1467 :   0 - 0x0
      11'h5BC: dout  = 8'b00000000; // 1468 :   0 - 0x0
      11'h5BD: dout  = 8'b00000000; // 1469 :   0 - 0x0
      11'h5BE: dout  = 8'b00000000; // 1470 :   0 - 0x0
      11'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      11'h5C1: dout  = 8'b00000011; // 1473 :   3 - 0x3
      11'h5C2: dout  = 8'b00000111; // 1474 :   7 - 0x7
      11'h5C3: dout  = 8'b00000111; // 1475 :   7 - 0x7
      11'h5C4: dout  = 8'b00000111; // 1476 :   7 - 0x7
      11'h5C5: dout  = 8'b00000011; // 1477 :   3 - 0x3
      11'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      11'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- Sprite 0xb9
      11'h5C9: dout  = 8'b11000001; // 1481 : 193 - 0xc1
      11'h5CA: dout  = 8'b11100010; // 1482 : 226 - 0xe2
      11'h5CB: dout  = 8'b11001100; // 1483 : 204 - 0xcc
      11'h5CC: dout  = 8'b11000000; // 1484 : 192 - 0xc0
      11'h5CD: dout  = 8'b10000000; // 1485 : 128 - 0x80
      11'h5CE: dout  = 8'b00000001; // 1486 :   1 - 0x1
      11'h5CF: dout  = 8'b00000010; // 1487 :   2 - 0x2
      11'h5D0: dout  = 8'b11110000; // 1488 : 240 - 0xf0 -- Sprite 0xba
      11'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      11'h5D2: dout  = 8'b00100000; // 1490 :  32 - 0x20
      11'h5D3: dout  = 8'b00100000; // 1491 :  32 - 0x20
      11'h5D4: dout  = 8'b00000000; // 1492 :   0 - 0x0
      11'h5D5: dout  = 8'b11110000; // 1493 : 240 - 0xf0
      11'h5D6: dout  = 8'b00000000; // 1494 :   0 - 0x0
      11'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      11'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      11'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      11'h5DD: dout  = 8'b01100000; // 1501 :  96 - 0x60
      11'h5DE: dout  = 8'b01100000; // 1502 :  96 - 0x60
      11'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout  = 8'b00001100; // 1504 :  12 - 0xc -- Sprite 0xbc
      11'h5E1: dout  = 8'b00000000; // 1505 :   0 - 0x0
      11'h5E2: dout  = 8'b00000000; // 1506 :   0 - 0x0
      11'h5E3: dout  = 8'b00000000; // 1507 :   0 - 0x0
      11'h5E4: dout  = 8'b00000000; // 1508 :   0 - 0x0
      11'h5E5: dout  = 8'b00000110; // 1509 :   6 - 0x6
      11'h5E6: dout  = 8'b00000110; // 1510 :   6 - 0x6
      11'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      11'h5E9: dout  = 8'b10000011; // 1513 : 131 - 0x83
      11'h5EA: dout  = 8'b00000111; // 1514 :   7 - 0x7
      11'h5EB: dout  = 8'b00000111; // 1515 :   7 - 0x7
      11'h5EC: dout  = 8'b00000111; // 1516 :   7 - 0x7
      11'h5ED: dout  = 8'b00000011; // 1517 :   3 - 0x3
      11'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      11'h5F1: dout  = 8'b11000100; // 1521 : 196 - 0xc4
      11'h5F2: dout  = 8'b11100000; // 1522 : 224 - 0xe0
      11'h5F3: dout  = 8'b11000000; // 1523 : 192 - 0xc0
      11'h5F4: dout  = 8'b11000000; // 1524 : 192 - 0xc0
      11'h5F5: dout  = 8'b10000000; // 1525 : 128 - 0x80
      11'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      11'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      11'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout  = 8'b00001000; // 1532 :   8 - 0x8
      11'h5FD: dout  = 8'b10001000; // 1533 : 136 - 0x88
      11'h5FE: dout  = 8'b00001011; // 1534 :  11 - 0xb
      11'h5FF: dout  = 8'b00001000; // 1535 :   8 - 0x8
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      11'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout  = 8'b00000000; // 1538 :   0 - 0x0
      11'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout  = 8'b00100000; // 1540 :  32 - 0x20
      11'h605: dout  = 8'b00100100; // 1541 :  36 - 0x24
      11'h606: dout  = 8'b10100000; // 1542 : 160 - 0xa0
      11'h607: dout  = 8'b00100000; // 1543 :  32 - 0x20
      11'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      11'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout  = 8'b00000000; // 1546 :   0 - 0x0
      11'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout  = 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      11'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout  = 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout  = 8'b00000000; // 1556 :   0 - 0x0
      11'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout  = 8'b00000000; // 1558 :   0 - 0x0
      11'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      11'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout  = 8'b00001000; // 1562 :   8 - 0x8
      11'h61B: dout  = 8'b00001011; // 1563 :  11 - 0xb
      11'h61C: dout  = 8'b00001000; // 1564 :   8 - 0x8
      11'h61D: dout  = 8'b00001000; // 1565 :   8 - 0x8
      11'h61E: dout  = 8'b00001000; // 1566 :   8 - 0x8
      11'h61F: dout  = 8'b00001000; // 1567 :   8 - 0x8
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout  = 8'b00100000; // 1570 :  32 - 0x20
      11'h623: dout  = 8'b10100000; // 1571 : 160 - 0xa0
      11'h624: dout  = 8'b00100000; // 1572 :  32 - 0x20
      11'h625: dout  = 8'b00100000; // 1573 :  32 - 0x20
      11'h626: dout  = 8'b00100000; // 1574 :  32 - 0x20
      11'h627: dout  = 8'b00100000; // 1575 :  32 - 0x20
      11'h628: dout  = 8'b00001000; // 1576 :   8 - 0x8 -- Sprite 0xc5
      11'h629: dout  = 8'b11001000; // 1577 : 200 - 0xc8
      11'h62A: dout  = 8'b00000011; // 1578 :   3 - 0x3
      11'h62B: dout  = 8'b00000111; // 1579 :   7 - 0x7
      11'h62C: dout  = 8'b00000111; // 1580 :   7 - 0x7
      11'h62D: dout  = 8'b00000111; // 1581 :   7 - 0x7
      11'h62E: dout  = 8'b00000011; // 1582 :   3 - 0x3
      11'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout  = 8'b00100000; // 1584 :  32 - 0x20 -- Sprite 0xc6
      11'h631: dout  = 8'b00100110; // 1585 :  38 - 0x26
      11'h632: dout  = 8'b11000000; // 1586 : 192 - 0xc0
      11'h633: dout  = 8'b11100000; // 1587 : 224 - 0xe0
      11'h634: dout  = 8'b11000000; // 1588 : 192 - 0xc0
      11'h635: dout  = 8'b11000000; // 1589 : 192 - 0xc0
      11'h636: dout  = 8'b10000000; // 1590 : 128 - 0x80
      11'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- Sprite 0xc7
      11'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      11'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      11'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      11'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      11'h63D: dout  = 8'b11000000; // 1597 : 192 - 0xc0
      11'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      11'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      11'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout  = 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout  = 8'b00000110; // 1605 :   6 - 0x6
      11'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout  = 8'b00001111; // 1608 :  15 - 0xf -- Sprite 0xc9
      11'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      11'h64A: dout  = 8'b00001000; // 1610 :   8 - 0x8
      11'h64B: dout  = 8'b00001000; // 1611 :   8 - 0x8
      11'h64C: dout  = 8'b00000000; // 1612 :   0 - 0x0
      11'h64D: dout  = 8'b00001111; // 1613 :  15 - 0xf
      11'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout  = 8'b10000011; // 1617 : 131 - 0x83
      11'h652: dout  = 8'b01000111; // 1618 :  71 - 0x47
      11'h653: dout  = 8'b00110111; // 1619 :  55 - 0x37
      11'h654: dout  = 8'b00000111; // 1620 :   7 - 0x7
      11'h655: dout  = 8'b00000011; // 1621 :   3 - 0x3
      11'h656: dout  = 8'b10000000; // 1622 : 128 - 0x80
      11'h657: dout  = 8'b01000000; // 1623 :  64 - 0x40
      11'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      11'h659: dout  = 8'b11000000; // 1625 : 192 - 0xc0
      11'h65A: dout  = 8'b11100000; // 1626 : 224 - 0xe0
      11'h65B: dout  = 8'b11000000; // 1627 : 192 - 0xc0
      11'h65C: dout  = 8'b11000000; // 1628 : 192 - 0xc0
      11'h65D: dout  = 8'b10000000; // 1629 : 128 - 0x80
      11'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout  = 8'b00110000; // 1632 :  48 - 0x30 -- Sprite 0xcc
      11'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      11'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      11'h665: dout  = 8'b01100000; // 1637 :  96 - 0x60
      11'h666: dout  = 8'b01100000; // 1638 :  96 - 0x60
      11'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      11'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout  = 8'b00000000; // 1643 :   0 - 0x0
      11'h66C: dout  = 8'b00000000; // 1644 :   0 - 0x0
      11'h66D: dout  = 8'b00000110; // 1645 :   6 - 0x6
      11'h66E: dout  = 8'b00000110; // 1646 :   6 - 0x6
      11'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      11'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      11'h671: dout  = 8'b00000001; // 1649 :   1 - 0x1
      11'h672: dout  = 8'b00011011; // 1650 :  27 - 0x1b
      11'h673: dout  = 8'b00010011; // 1651 :  19 - 0x13
      11'h674: dout  = 8'b00011111; // 1652 :  31 - 0x1f
      11'h675: dout  = 8'b00111111; // 1653 :  63 - 0x3f
      11'h676: dout  = 8'b00111111; // 1654 :  63 - 0x3f
      11'h677: dout  = 8'b00111111; // 1655 :  63 - 0x3f
      11'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      11'h679: dout  = 8'b11111000; // 1657 : 248 - 0xf8
      11'h67A: dout  = 8'b00001000; // 1658 :   8 - 0x8
      11'h67B: dout  = 8'b00001000; // 1659 :   8 - 0x8
      11'h67C: dout  = 8'b00001000; // 1660 :   8 - 0x8
      11'h67D: dout  = 8'b11111000; // 1661 : 248 - 0xf8
      11'h67E: dout  = 8'b11110000; // 1662 : 240 - 0xf0
      11'h67F: dout  = 8'b11010000; // 1663 : 208 - 0xd0
      11'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      11'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout  = 8'b01111100; // 1666 : 124 - 0x7c
      11'h683: dout  = 8'b11111110; // 1667 : 254 - 0xfe
      11'h684: dout  = 8'b11101110; // 1668 : 238 - 0xee
      11'h685: dout  = 8'b11101110; // 1669 : 238 - 0xee
      11'h686: dout  = 8'b11101110; // 1670 : 238 - 0xee
      11'h687: dout  = 8'b11101110; // 1671 : 238 - 0xee
      11'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      11'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout  = 8'b00111000; // 1674 :  56 - 0x38
      11'h68B: dout  = 8'b01111000; // 1675 : 120 - 0x78
      11'h68C: dout  = 8'b01111000; // 1676 : 120 - 0x78
      11'h68D: dout  = 8'b00111000; // 1677 :  56 - 0x38
      11'h68E: dout  = 8'b00111000; // 1678 :  56 - 0x38
      11'h68F: dout  = 8'b00111000; // 1679 :  56 - 0x38
      11'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      11'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout  = 8'b01111100; // 1682 : 124 - 0x7c
      11'h693: dout  = 8'b11111110; // 1683 : 254 - 0xfe
      11'h694: dout  = 8'b11101110; // 1684 : 238 - 0xee
      11'h695: dout  = 8'b00001110; // 1685 :  14 - 0xe
      11'h696: dout  = 8'b00001110; // 1686 :  14 - 0xe
      11'h697: dout  = 8'b01111110; // 1687 : 126 - 0x7e
      11'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0 -- Sprite 0xd3
      11'h699: dout  = 8'b00000000; // 1689 :   0 - 0x0
      11'h69A: dout  = 8'b01111100; // 1690 : 124 - 0x7c
      11'h69B: dout  = 8'b11111110; // 1691 : 254 - 0xfe
      11'h69C: dout  = 8'b11101110; // 1692 : 238 - 0xee
      11'h69D: dout  = 8'b00001110; // 1693 :  14 - 0xe
      11'h69E: dout  = 8'b00111100; // 1694 :  60 - 0x3c
      11'h69F: dout  = 8'b00111100; // 1695 :  60 - 0x3c
      11'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      11'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout  = 8'b00111110; // 1698 :  62 - 0x3e
      11'h6A3: dout  = 8'b01111110; // 1699 : 126 - 0x7e
      11'h6A4: dout  = 8'b11101110; // 1700 : 238 - 0xee
      11'h6A5: dout  = 8'b11101110; // 1701 : 238 - 0xee
      11'h6A6: dout  = 8'b11101110; // 1702 : 238 - 0xee
      11'h6A7: dout  = 8'b11101110; // 1703 : 238 - 0xee
      11'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      11'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      11'h6AA: dout  = 8'b11111100; // 1706 : 252 - 0xfc
      11'h6AB: dout  = 8'b11111100; // 1707 : 252 - 0xfc
      11'h6AC: dout  = 8'b11100000; // 1708 : 224 - 0xe0
      11'h6AD: dout  = 8'b11100000; // 1709 : 224 - 0xe0
      11'h6AE: dout  = 8'b11111100; // 1710 : 252 - 0xfc
      11'h6AF: dout  = 8'b11111110; // 1711 : 254 - 0xfe
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b01111100; // 1714 : 124 - 0x7c
      11'h6B3: dout  = 8'b11111100; // 1715 : 252 - 0xfc
      11'h6B4: dout  = 8'b11100000; // 1716 : 224 - 0xe0
      11'h6B5: dout  = 8'b11100000; // 1717 : 224 - 0xe0
      11'h6B6: dout  = 8'b11111100; // 1718 : 252 - 0xfc
      11'h6B7: dout  = 8'b11111110; // 1719 : 254 - 0xfe
      11'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0 -- Sprite 0xd7
      11'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      11'h6BA: dout  = 8'b11111110; // 1722 : 254 - 0xfe
      11'h6BB: dout  = 8'b11111110; // 1723 : 254 - 0xfe
      11'h6BC: dout  = 8'b11101110; // 1724 : 238 - 0xee
      11'h6BD: dout  = 8'b00001110; // 1725 :  14 - 0xe
      11'h6BE: dout  = 8'b00001110; // 1726 :  14 - 0xe
      11'h6BF: dout  = 8'b00011100; // 1727 :  28 - 0x1c
      11'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      11'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout  = 8'b01111100; // 1730 : 124 - 0x7c
      11'h6C3: dout  = 8'b11111110; // 1731 : 254 - 0xfe
      11'h6C4: dout  = 8'b11101110; // 1732 : 238 - 0xee
      11'h6C5: dout  = 8'b11101110; // 1733 : 238 - 0xee
      11'h6C6: dout  = 8'b01111100; // 1734 : 124 - 0x7c
      11'h6C7: dout  = 8'b11111110; // 1735 : 254 - 0xfe
      11'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      11'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      11'h6CA: dout  = 8'b01111100; // 1738 : 124 - 0x7c
      11'h6CB: dout  = 8'b11111110; // 1739 : 254 - 0xfe
      11'h6CC: dout  = 8'b11101110; // 1740 : 238 - 0xee
      11'h6CD: dout  = 8'b11101110; // 1741 : 238 - 0xee
      11'h6CE: dout  = 8'b11101110; // 1742 : 238 - 0xee
      11'h6CF: dout  = 8'b11101110; // 1743 : 238 - 0xee
      11'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      11'h6D1: dout  = 8'b00100000; // 1745 :  32 - 0x20
      11'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      11'h6D3: dout  = 8'b00000010; // 1747 :   2 - 0x2
      11'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout  = 8'b00100000; // 1749 :  32 - 0x20
      11'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      11'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout  = 8'b00100000; // 1752 :  32 - 0x20 -- Sprite 0xdb
      11'h6D9: dout  = 8'b00000000; // 1753 :   0 - 0x0
      11'h6DA: dout  = 8'b00000000; // 1754 :   0 - 0x0
      11'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      11'h6DC: dout  = 8'b10000000; // 1756 : 128 - 0x80
      11'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      11'h6DE: dout  = 8'b00000100; // 1758 :   4 - 0x4
      11'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      11'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      11'h6E1: dout  = 8'b00001000; // 1761 :   8 - 0x8
      11'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      11'h6E4: dout  = 8'b00000010; // 1764 :   2 - 0x2
      11'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      11'h6E6: dout  = 8'b01000000; // 1766 :  64 - 0x40
      11'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      11'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      11'h6E9: dout  = 8'b01000000; // 1769 :  64 - 0x40
      11'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      11'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      11'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      11'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      11'h6EE: dout  = 8'b00000010; // 1774 :   2 - 0x2
      11'h6EF: dout  = 8'b00100000; // 1775 :  32 - 0x20
      11'h6F0: dout  = 8'b00111110; // 1776 :  62 - 0x3e -- Sprite 0xde
      11'h6F1: dout  = 8'b00111111; // 1777 :  63 - 0x3f
      11'h6F2: dout  = 8'b00111110; // 1778 :  62 - 0x3e
      11'h6F3: dout  = 8'b00111100; // 1779 :  60 - 0x3c
      11'h6F4: dout  = 8'b00111111; // 1780 :  63 - 0x3f
      11'h6F5: dout  = 8'b00110000; // 1781 :  48 - 0x30
      11'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      11'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      11'h6F8: dout  = 8'b00010000; // 1784 :  16 - 0x10 -- Sprite 0xdf
      11'h6F9: dout  = 8'b10110000; // 1785 : 176 - 0xb0
      11'h6FA: dout  = 8'b00110000; // 1786 :  48 - 0x30
      11'h6FB: dout  = 8'b11110000; // 1787 : 240 - 0xf0
      11'h6FC: dout  = 8'b11110000; // 1788 : 240 - 0xf0
      11'h6FD: dout  = 8'b00000000; // 1789 :   0 - 0x0
      11'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      11'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      11'h700: dout  = 8'b11101110; // 1792 : 238 - 0xee -- Sprite 0xe0
      11'h701: dout  = 8'b11101110; // 1793 : 238 - 0xee
      11'h702: dout  = 8'b11101110; // 1794 : 238 - 0xee
      11'h703: dout  = 8'b11101110; // 1795 : 238 - 0xee
      11'h704: dout  = 8'b11111110; // 1796 : 254 - 0xfe
      11'h705: dout  = 8'b01111100; // 1797 : 124 - 0x7c
      11'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      11'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout  = 8'b00111000; // 1800 :  56 - 0x38 -- Sprite 0xe1
      11'h709: dout  = 8'b00111000; // 1801 :  56 - 0x38
      11'h70A: dout  = 8'b00111000; // 1802 :  56 - 0x38
      11'h70B: dout  = 8'b00111000; // 1803 :  56 - 0x38
      11'h70C: dout  = 8'b01111100; // 1804 : 124 - 0x7c
      11'h70D: dout  = 8'b01111100; // 1805 : 124 - 0x7c
      11'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout  = 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      11'h711: dout  = 8'b11100000; // 1809 : 224 - 0xe0
      11'h712: dout  = 8'b11100000; // 1810 : 224 - 0xe0
      11'h713: dout  = 8'b11100000; // 1811 : 224 - 0xe0
      11'h714: dout  = 8'b11111110; // 1812 : 254 - 0xfe
      11'h715: dout  = 8'b11111110; // 1813 : 254 - 0xfe
      11'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout  = 8'b00001110; // 1816 :  14 - 0xe -- Sprite 0xe3
      11'h719: dout  = 8'b00001110; // 1817 :  14 - 0xe
      11'h71A: dout  = 8'b00001110; // 1818 :  14 - 0xe
      11'h71B: dout  = 8'b11101110; // 1819 : 238 - 0xee
      11'h71C: dout  = 8'b11111110; // 1820 : 254 - 0xfe
      11'h71D: dout  = 8'b01111100; // 1821 : 124 - 0x7c
      11'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      11'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      11'h720: dout  = 8'b11101110; // 1824 : 238 - 0xee -- Sprite 0xe4
      11'h721: dout  = 8'b11101110; // 1825 : 238 - 0xee
      11'h722: dout  = 8'b11111110; // 1826 : 254 - 0xfe
      11'h723: dout  = 8'b11111110; // 1827 : 254 - 0xfe
      11'h724: dout  = 8'b00001110; // 1828 :  14 - 0xe
      11'h725: dout  = 8'b00001110; // 1829 :  14 - 0xe
      11'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      11'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      11'h728: dout  = 8'b00001110; // 1832 :  14 - 0xe -- Sprite 0xe5
      11'h729: dout  = 8'b00001110; // 1833 :  14 - 0xe
      11'h72A: dout  = 8'b00001110; // 1834 :  14 - 0xe
      11'h72B: dout  = 8'b11101110; // 1835 : 238 - 0xee
      11'h72C: dout  = 8'b11111110; // 1836 : 254 - 0xfe
      11'h72D: dout  = 8'b01111100; // 1837 : 124 - 0x7c
      11'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      11'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      11'h730: dout  = 8'b11101110; // 1840 : 238 - 0xee -- Sprite 0xe6
      11'h731: dout  = 8'b11101110; // 1841 : 238 - 0xee
      11'h732: dout  = 8'b11101110; // 1842 : 238 - 0xee
      11'h733: dout  = 8'b11101110; // 1843 : 238 - 0xee
      11'h734: dout  = 8'b11111110; // 1844 : 254 - 0xfe
      11'h735: dout  = 8'b01111100; // 1845 : 124 - 0x7c
      11'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      11'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout  = 8'b00011100; // 1848 :  28 - 0x1c -- Sprite 0xe7
      11'h739: dout  = 8'b00011100; // 1849 :  28 - 0x1c
      11'h73A: dout  = 8'b00111000; // 1850 :  56 - 0x38
      11'h73B: dout  = 8'b00111000; // 1851 :  56 - 0x38
      11'h73C: dout  = 8'b00111000; // 1852 :  56 - 0x38
      11'h73D: dout  = 8'b00111000; // 1853 :  56 - 0x38
      11'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      11'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      11'h740: dout  = 8'b11101110; // 1856 : 238 - 0xee -- Sprite 0xe8
      11'h741: dout  = 8'b11101110; // 1857 : 238 - 0xee
      11'h742: dout  = 8'b11101110; // 1858 : 238 - 0xee
      11'h743: dout  = 8'b11101110; // 1859 : 238 - 0xee
      11'h744: dout  = 8'b11111110; // 1860 : 254 - 0xfe
      11'h745: dout  = 8'b01111100; // 1861 : 124 - 0x7c
      11'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout  = 8'b11111110; // 1864 : 254 - 0xfe -- Sprite 0xe9
      11'h749: dout  = 8'b01111110; // 1865 : 126 - 0x7e
      11'h74A: dout  = 8'b00001110; // 1866 :  14 - 0xe
      11'h74B: dout  = 8'b00001110; // 1867 :  14 - 0xe
      11'h74C: dout  = 8'b01111110; // 1868 : 126 - 0x7e
      11'h74D: dout  = 8'b01111100; // 1869 : 124 - 0x7c
      11'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      11'h751: dout  = 8'b01110000; // 1873 : 112 - 0x70
      11'h752: dout  = 8'b00111000; // 1874 :  56 - 0x38
      11'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout  = 8'b00000010; // 1876 :   2 - 0x2
      11'h755: dout  = 8'b00000111; // 1877 :   7 - 0x7
      11'h756: dout  = 8'b00000011; // 1878 :   3 - 0x3
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      11'h759: dout  = 8'b00001100; // 1881 :  12 - 0xc
      11'h75A: dout  = 8'b00000110; // 1882 :   6 - 0x6
      11'h75B: dout  = 8'b00000110; // 1883 :   6 - 0x6
      11'h75C: dout  = 8'b01100000; // 1884 :  96 - 0x60
      11'h75D: dout  = 8'b01110000; // 1885 : 112 - 0x70
      11'h75E: dout  = 8'b00110000; // 1886 :  48 - 0x30
      11'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout  = 8'b11000000; // 1889 : 192 - 0xc0
      11'h762: dout  = 8'b11100000; // 1890 : 224 - 0xe0
      11'h763: dout  = 8'b01100000; // 1891 :  96 - 0x60
      11'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout  = 8'b00001100; // 1893 :  12 - 0xc
      11'h766: dout  = 8'b00001110; // 1894 :  14 - 0xe
      11'h767: dout  = 8'b00000110; // 1895 :   6 - 0x6
      11'h768: dout  = 8'b01100000; // 1896 :  96 - 0x60 -- Sprite 0xed
      11'h769: dout  = 8'b01110000; // 1897 : 112 - 0x70
      11'h76A: dout  = 8'b00110000; // 1898 :  48 - 0x30
      11'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout  = 8'b00001100; // 1901 :  12 - 0xc
      11'h76E: dout  = 8'b00001110; // 1902 :  14 - 0xe
      11'h76F: dout  = 8'b00000110; // 1903 :   6 - 0x6
      11'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      11'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout  = 8'b01000010; // 1906 :  66 - 0x42
      11'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout  = 8'b00000100; // 1909 :   4 - 0x4
      11'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      11'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      11'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout  = 8'b00000100; // 1914 :   4 - 0x4
      11'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout  = 8'b00100000; // 1916 :  32 - 0x20
      11'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      11'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      11'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      11'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout  = 8'b10000000; // 1928 : 128 - 0x80 -- Sprite 0xf1
      11'h789: dout  = 8'b10000000; // 1929 : 128 - 0x80
      11'h78A: dout  = 8'b10000000; // 1930 : 128 - 0x80
      11'h78B: dout  = 8'b10000000; // 1931 : 128 - 0x80
      11'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      11'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      11'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout  = 8'b11000000; // 1936 : 192 - 0xc0 -- Sprite 0xf2
      11'h791: dout  = 8'b11000000; // 1937 : 192 - 0xc0
      11'h792: dout  = 8'b11000000; // 1938 : 192 - 0xc0
      11'h793: dout  = 8'b11000000; // 1939 : 192 - 0xc0
      11'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      11'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      11'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      11'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      11'h798: dout  = 8'b11100000; // 1944 : 224 - 0xe0 -- Sprite 0xf3
      11'h799: dout  = 8'b11100000; // 1945 : 224 - 0xe0
      11'h79A: dout  = 8'b11100000; // 1946 : 224 - 0xe0
      11'h79B: dout  = 8'b11100000; // 1947 : 224 - 0xe0
      11'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      11'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout  = 8'b11110000; // 1952 : 240 - 0xf0 -- Sprite 0xf4
      11'h7A1: dout  = 8'b11110000; // 1953 : 240 - 0xf0
      11'h7A2: dout  = 8'b11110000; // 1954 : 240 - 0xf0
      11'h7A3: dout  = 8'b11110000; // 1955 : 240 - 0xf0
      11'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      11'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      11'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout  = 8'b11111000; // 1960 : 248 - 0xf8 -- Sprite 0xf5
      11'h7A9: dout  = 8'b11111000; // 1961 : 248 - 0xf8
      11'h7AA: dout  = 8'b11111000; // 1962 : 248 - 0xf8
      11'h7AB: dout  = 8'b11111000; // 1963 : 248 - 0xf8
      11'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      11'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      11'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout  = 8'b11111100; // 1968 : 252 - 0xfc -- Sprite 0xf6
      11'h7B1: dout  = 8'b11111100; // 1969 : 252 - 0xfc
      11'h7B2: dout  = 8'b11111100; // 1970 : 252 - 0xfc
      11'h7B3: dout  = 8'b11111100; // 1971 : 252 - 0xfc
      11'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout  = 8'b11111110; // 1976 : 254 - 0xfe -- Sprite 0xf7
      11'h7B9: dout  = 8'b11111110; // 1977 : 254 - 0xfe
      11'h7BA: dout  = 8'b11111110; // 1978 : 254 - 0xfe
      11'h7BB: dout  = 8'b11111110; // 1979 : 254 - 0xfe
      11'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout  = 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0xf8
      11'h7C1: dout  = 8'b11111111; // 1985 : 255 - 0xff
      11'h7C2: dout  = 8'b11111111; // 1986 : 255 - 0xff
      11'h7C3: dout  = 8'b11111111; // 1987 : 255 - 0xff
      11'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      11'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout  = 8'b01111111; // 1996 : 127 - 0x7f
      11'h7CD: dout  = 8'b01000000; // 1997 :  64 - 0x40
      11'h7CE: dout  = 8'b01000000; // 1998 :  64 - 0x40
      11'h7CF: dout  = 8'b01000000; // 1999 :  64 - 0x40
      11'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      11'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout  = 8'b11111111; // 2004 : 255 - 0xff
      11'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      11'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout  = 8'b11111110; // 2012 : 254 - 0xfe
      11'h7DD: dout  = 8'b00000010; // 2013 :   2 - 0x2
      11'h7DE: dout  = 8'b00000010; // 2014 :   2 - 0x2
      11'h7DF: dout  = 8'b00000010; // 2015 :   2 - 0x2
      11'h7E0: dout  = 8'b01000000; // 2016 :  64 - 0x40 -- Sprite 0xfc
      11'h7E1: dout  = 8'b01000000; // 2017 :  64 - 0x40
      11'h7E2: dout  = 8'b01000000; // 2018 :  64 - 0x40
      11'h7E3: dout  = 8'b01111111; // 2019 : 127 - 0x7f
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      11'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout  = 8'b11111111; // 2027 : 255 - 0xff
      11'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00000010; // 2032 :   2 - 0x2 -- Sprite 0xfe
      11'h7F1: dout  = 8'b00000010; // 2033 :   2 - 0x2
      11'h7F2: dout  = 8'b00000010; // 2034 :   2 - 0x2
      11'h7F3: dout  = 8'b11111110; // 2035 : 254 - 0xfe
      11'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
