---   Background Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: smario_traspas_patron.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_MARIO_TRASPAS_BG_PLN0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_MARIO_TRASPAS_BG_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_MARIO_TRASPAS_BG_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 0
    "00111000", --    0 -  0x0  :   56 - 0x38 -- Background 0x0
    "01001100", --    1 -  0x1  :   76 - 0x4c
    "11000110", --    2 -  0x2  :  198 - 0xc6
    "11000110", --    3 -  0x3  :  198 - 0xc6
    "11000110", --    4 -  0x4  :  198 - 0xc6
    "01100100", --    5 -  0x5  :  100 - 0x64
    "00111000", --    6 -  0x6  :   56 - 0x38
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00011000", --    8 -  0x8  :   24 - 0x18 -- Background 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "00011000", --   10 -  0xa  :   24 - 0x18
    "00011000", --   11 -  0xb  :   24 - 0x18
    "00011000", --   12 -  0xc  :   24 - 0x18
    "00011000", --   13 -  0xd  :   24 - 0x18
    "01111110", --   14 -  0xe  :  126 - 0x7e
    "00000000", --   15 -  0xf  :    0 - 0x0
    "01111100", --   16 - 0x10  :  124 - 0x7c -- Background 0x2
    "11000110", --   17 - 0x11  :  198 - 0xc6
    "00001110", --   18 - 0x12  :   14 - 0xe
    "00111100", --   19 - 0x13  :   60 - 0x3c
    "01111000", --   20 - 0x14  :  120 - 0x78
    "11100000", --   21 - 0x15  :  224 - 0xe0
    "11111110", --   22 - 0x16  :  254 - 0xfe
    "00000000", --   23 - 0x17  :    0 - 0x0
    "01111110", --   24 - 0x18  :  126 - 0x7e -- Background 0x3
    "00001100", --   25 - 0x19  :   12 - 0xc
    "00011000", --   26 - 0x1a  :   24 - 0x18
    "00111100", --   27 - 0x1b  :   60 - 0x3c
    "00000110", --   28 - 0x1c  :    6 - 0x6
    "11000110", --   29 - 0x1d  :  198 - 0xc6
    "01111100", --   30 - 0x1e  :  124 - 0x7c
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00011100", --   32 - 0x20  :   28 - 0x1c -- Background 0x4
    "00111100", --   33 - 0x21  :   60 - 0x3c
    "01101100", --   34 - 0x22  :  108 - 0x6c
    "11001100", --   35 - 0x23  :  204 - 0xcc
    "11111110", --   36 - 0x24  :  254 - 0xfe
    "00001100", --   37 - 0x25  :   12 - 0xc
    "00001100", --   38 - 0x26  :   12 - 0xc
    "00000000", --   39 - 0x27  :    0 - 0x0
    "11111100", --   40 - 0x28  :  252 - 0xfc -- Background 0x5
    "11000000", --   41 - 0x29  :  192 - 0xc0
    "11111100", --   42 - 0x2a  :  252 - 0xfc
    "00000110", --   43 - 0x2b  :    6 - 0x6
    "00000110", --   44 - 0x2c  :    6 - 0x6
    "11000110", --   45 - 0x2d  :  198 - 0xc6
    "01111100", --   46 - 0x2e  :  124 - 0x7c
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00111100", --   48 - 0x30  :   60 - 0x3c -- Background 0x6
    "01100000", --   49 - 0x31  :   96 - 0x60
    "11000000", --   50 - 0x32  :  192 - 0xc0
    "11111100", --   51 - 0x33  :  252 - 0xfc
    "11000110", --   52 - 0x34  :  198 - 0xc6
    "11000110", --   53 - 0x35  :  198 - 0xc6
    "01111100", --   54 - 0x36  :  124 - 0x7c
    "00000000", --   55 - 0x37  :    0 - 0x0
    "11111110", --   56 - 0x38  :  254 - 0xfe -- Background 0x7
    "11000110", --   57 - 0x39  :  198 - 0xc6
    "00001100", --   58 - 0x3a  :   12 - 0xc
    "00011000", --   59 - 0x3b  :   24 - 0x18
    "00110000", --   60 - 0x3c  :   48 - 0x30
    "00110000", --   61 - 0x3d  :   48 - 0x30
    "00110000", --   62 - 0x3e  :   48 - 0x30
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "01111100", --   64 - 0x40  :  124 - 0x7c -- Background 0x8
    "11000110", --   65 - 0x41  :  198 - 0xc6
    "11000110", --   66 - 0x42  :  198 - 0xc6
    "01111100", --   67 - 0x43  :  124 - 0x7c
    "11000110", --   68 - 0x44  :  198 - 0xc6
    "11000110", --   69 - 0x45  :  198 - 0xc6
    "01111100", --   70 - 0x46  :  124 - 0x7c
    "00000000", --   71 - 0x47  :    0 - 0x0
    "01111100", --   72 - 0x48  :  124 - 0x7c -- Background 0x9
    "11000110", --   73 - 0x49  :  198 - 0xc6
    "11000110", --   74 - 0x4a  :  198 - 0xc6
    "01111110", --   75 - 0x4b  :  126 - 0x7e
    "00000110", --   76 - 0x4c  :    6 - 0x6
    "00001100", --   77 - 0x4d  :   12 - 0xc
    "01111000", --   78 - 0x4e  :  120 - 0x78
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00111000", --   80 - 0x50  :   56 - 0x38 -- Background 0xa
    "01101100", --   81 - 0x51  :  108 - 0x6c
    "11000110", --   82 - 0x52  :  198 - 0xc6
    "11000110", --   83 - 0x53  :  198 - 0xc6
    "11111110", --   84 - 0x54  :  254 - 0xfe
    "11000110", --   85 - 0x55  :  198 - 0xc6
    "11000110", --   86 - 0x56  :  198 - 0xc6
    "00000000", --   87 - 0x57  :    0 - 0x0
    "11111100", --   88 - 0x58  :  252 - 0xfc -- Background 0xb
    "11000110", --   89 - 0x59  :  198 - 0xc6
    "11000110", --   90 - 0x5a  :  198 - 0xc6
    "11111100", --   91 - 0x5b  :  252 - 0xfc
    "11000110", --   92 - 0x5c  :  198 - 0xc6
    "11000110", --   93 - 0x5d  :  198 - 0xc6
    "11111100", --   94 - 0x5e  :  252 - 0xfc
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00111100", --   96 - 0x60  :   60 - 0x3c -- Background 0xc
    "01100110", --   97 - 0x61  :  102 - 0x66
    "11000000", --   98 - 0x62  :  192 - 0xc0
    "11000000", --   99 - 0x63  :  192 - 0xc0
    "11000000", --  100 - 0x64  :  192 - 0xc0
    "01100110", --  101 - 0x65  :  102 - 0x66
    "00111100", --  102 - 0x66  :   60 - 0x3c
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11111000", --  104 - 0x68  :  248 - 0xf8 -- Background 0xd
    "11001100", --  105 - 0x69  :  204 - 0xcc
    "11000110", --  106 - 0x6a  :  198 - 0xc6
    "11000110", --  107 - 0x6b  :  198 - 0xc6
    "11000110", --  108 - 0x6c  :  198 - 0xc6
    "11001100", --  109 - 0x6d  :  204 - 0xcc
    "11111000", --  110 - 0x6e  :  248 - 0xf8
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11111110", --  112 - 0x70  :  254 - 0xfe -- Background 0xe
    "11000000", --  113 - 0x71  :  192 - 0xc0
    "11000000", --  114 - 0x72  :  192 - 0xc0
    "11111100", --  115 - 0x73  :  252 - 0xfc
    "11000000", --  116 - 0x74  :  192 - 0xc0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "11111110", --  118 - 0x76  :  254 - 0xfe
    "00000000", --  119 - 0x77  :    0 - 0x0
    "11111110", --  120 - 0x78  :  254 - 0xfe -- Background 0xf
    "11000000", --  121 - 0x79  :  192 - 0xc0
    "11000000", --  122 - 0x7a  :  192 - 0xc0
    "11111100", --  123 - 0x7b  :  252 - 0xfc
    "11000000", --  124 - 0x7c  :  192 - 0xc0
    "11000000", --  125 - 0x7d  :  192 - 0xc0
    "11000000", --  126 - 0x7e  :  192 - 0xc0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00111110", --  128 - 0x80  :   62 - 0x3e -- Background 0x10
    "01100000", --  129 - 0x81  :   96 - 0x60
    "11000000", --  130 - 0x82  :  192 - 0xc0
    "11001110", --  131 - 0x83  :  206 - 0xce
    "11000110", --  132 - 0x84  :  198 - 0xc6
    "01100110", --  133 - 0x85  :  102 - 0x66
    "00111110", --  134 - 0x86  :   62 - 0x3e
    "00000000", --  135 - 0x87  :    0 - 0x0
    "11000110", --  136 - 0x88  :  198 - 0xc6 -- Background 0x11
    "11000110", --  137 - 0x89  :  198 - 0xc6
    "11000110", --  138 - 0x8a  :  198 - 0xc6
    "11111110", --  139 - 0x8b  :  254 - 0xfe
    "11000110", --  140 - 0x8c  :  198 - 0xc6
    "11000110", --  141 - 0x8d  :  198 - 0xc6
    "11000110", --  142 - 0x8e  :  198 - 0xc6
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01111110", --  144 - 0x90  :  126 - 0x7e -- Background 0x12
    "00011000", --  145 - 0x91  :   24 - 0x18
    "00011000", --  146 - 0x92  :   24 - 0x18
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00011000", --  148 - 0x94  :   24 - 0x18
    "00011000", --  149 - 0x95  :   24 - 0x18
    "01111110", --  150 - 0x96  :  126 - 0x7e
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00011110", --  152 - 0x98  :   30 - 0x1e -- Background 0x13
    "00000110", --  153 - 0x99  :    6 - 0x6
    "00000110", --  154 - 0x9a  :    6 - 0x6
    "00000110", --  155 - 0x9b  :    6 - 0x6
    "11000110", --  156 - 0x9c  :  198 - 0xc6
    "11000110", --  157 - 0x9d  :  198 - 0xc6
    "01111100", --  158 - 0x9e  :  124 - 0x7c
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "11000110", --  160 - 0xa0  :  198 - 0xc6 -- Background 0x14
    "11001100", --  161 - 0xa1  :  204 - 0xcc
    "11011000", --  162 - 0xa2  :  216 - 0xd8
    "11110000", --  163 - 0xa3  :  240 - 0xf0
    "11111000", --  164 - 0xa4  :  248 - 0xf8
    "11011100", --  165 - 0xa5  :  220 - 0xdc
    "11001110", --  166 - 0xa6  :  206 - 0xce
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "01100000", --  168 - 0xa8  :   96 - 0x60 -- Background 0x15
    "01100000", --  169 - 0xa9  :   96 - 0x60
    "01100000", --  170 - 0xaa  :   96 - 0x60
    "01100000", --  171 - 0xab  :   96 - 0x60
    "01100000", --  172 - 0xac  :   96 - 0x60
    "01100000", --  173 - 0xad  :   96 - 0x60
    "01111110", --  174 - 0xae  :  126 - 0x7e
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11000110", --  176 - 0xb0  :  198 - 0xc6 -- Background 0x16
    "11101110", --  177 - 0xb1  :  238 - 0xee
    "11111110", --  178 - 0xb2  :  254 - 0xfe
    "11111110", --  179 - 0xb3  :  254 - 0xfe
    "11010110", --  180 - 0xb4  :  214 - 0xd6
    "11000110", --  181 - 0xb5  :  198 - 0xc6
    "11000110", --  182 - 0xb6  :  198 - 0xc6
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "11000110", --  184 - 0xb8  :  198 - 0xc6 -- Background 0x17
    "11100110", --  185 - 0xb9  :  230 - 0xe6
    "11110110", --  186 - 0xba  :  246 - 0xf6
    "11111110", --  187 - 0xbb  :  254 - 0xfe
    "11011110", --  188 - 0xbc  :  222 - 0xde
    "11001110", --  189 - 0xbd  :  206 - 0xce
    "11000110", --  190 - 0xbe  :  198 - 0xc6
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "01111100", --  192 - 0xc0  :  124 - 0x7c -- Background 0x18
    "11000110", --  193 - 0xc1  :  198 - 0xc6
    "11000110", --  194 - 0xc2  :  198 - 0xc6
    "11000110", --  195 - 0xc3  :  198 - 0xc6
    "11000110", --  196 - 0xc4  :  198 - 0xc6
    "11000110", --  197 - 0xc5  :  198 - 0xc6
    "01111100", --  198 - 0xc6  :  124 - 0x7c
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "11111100", --  200 - 0xc8  :  252 - 0xfc -- Background 0x19
    "11000110", --  201 - 0xc9  :  198 - 0xc6
    "11000110", --  202 - 0xca  :  198 - 0xc6
    "11000110", --  203 - 0xcb  :  198 - 0xc6
    "11111100", --  204 - 0xcc  :  252 - 0xfc
    "11000000", --  205 - 0xcd  :  192 - 0xc0
    "11000000", --  206 - 0xce  :  192 - 0xc0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "01111100", --  208 - 0xd0  :  124 - 0x7c -- Background 0x1a
    "11000110", --  209 - 0xd1  :  198 - 0xc6
    "11000110", --  210 - 0xd2  :  198 - 0xc6
    "11000110", --  211 - 0xd3  :  198 - 0xc6
    "11011110", --  212 - 0xd4  :  222 - 0xde
    "11001100", --  213 - 0xd5  :  204 - 0xcc
    "01111010", --  214 - 0xd6  :  122 - 0x7a
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "11111100", --  216 - 0xd8  :  252 - 0xfc -- Background 0x1b
    "11000110", --  217 - 0xd9  :  198 - 0xc6
    "11000110", --  218 - 0xda  :  198 - 0xc6
    "11001110", --  219 - 0xdb  :  206 - 0xce
    "11111000", --  220 - 0xdc  :  248 - 0xf8
    "11011100", --  221 - 0xdd  :  220 - 0xdc
    "11001110", --  222 - 0xde  :  206 - 0xce
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "01111000", --  224 - 0xe0  :  120 - 0x78 -- Background 0x1c
    "11001100", --  225 - 0xe1  :  204 - 0xcc
    "11000000", --  226 - 0xe2  :  192 - 0xc0
    "01111100", --  227 - 0xe3  :  124 - 0x7c
    "00000110", --  228 - 0xe4  :    6 - 0x6
    "11000110", --  229 - 0xe5  :  198 - 0xc6
    "01111100", --  230 - 0xe6  :  124 - 0x7c
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "01111110", --  232 - 0xe8  :  126 - 0x7e -- Background 0x1d
    "00011000", --  233 - 0xe9  :   24 - 0x18
    "00011000", --  234 - 0xea  :   24 - 0x18
    "00011000", --  235 - 0xeb  :   24 - 0x18
    "00011000", --  236 - 0xec  :   24 - 0x18
    "00011000", --  237 - 0xed  :   24 - 0x18
    "00011000", --  238 - 0xee  :   24 - 0x18
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11000110", --  240 - 0xf0  :  198 - 0xc6 -- Background 0x1e
    "11000110", --  241 - 0xf1  :  198 - 0xc6
    "11000110", --  242 - 0xf2  :  198 - 0xc6
    "11000110", --  243 - 0xf3  :  198 - 0xc6
    "11000110", --  244 - 0xf4  :  198 - 0xc6
    "11000110", --  245 - 0xf5  :  198 - 0xc6
    "01111100", --  246 - 0xf6  :  124 - 0x7c
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "11000110", --  248 - 0xf8  :  198 - 0xc6 -- Background 0x1f
    "11000110", --  249 - 0xf9  :  198 - 0xc6
    "11000110", --  250 - 0xfa  :  198 - 0xc6
    "11101110", --  251 - 0xfb  :  238 - 0xee
    "01111100", --  252 - 0xfc  :  124 - 0x7c
    "00111000", --  253 - 0xfd  :   56 - 0x38
    "00010000", --  254 - 0xfe  :   16 - 0x10
    "00000000", --  255 - 0xff  :    0 - 0x0
    "11000110", --  256 - 0x100  :  198 - 0xc6 -- Background 0x20
    "11000110", --  257 - 0x101  :  198 - 0xc6
    "11010110", --  258 - 0x102  :  214 - 0xd6
    "11111110", --  259 - 0x103  :  254 - 0xfe
    "11111110", --  260 - 0x104  :  254 - 0xfe
    "11101110", --  261 - 0x105  :  238 - 0xee
    "11000110", --  262 - 0x106  :  198 - 0xc6
    "00000000", --  263 - 0x107  :    0 - 0x0
    "11000110", --  264 - 0x108  :  198 - 0xc6 -- Background 0x21
    "11101110", --  265 - 0x109  :  238 - 0xee
    "01111100", --  266 - 0x10a  :  124 - 0x7c
    "00111000", --  267 - 0x10b  :   56 - 0x38
    "01111100", --  268 - 0x10c  :  124 - 0x7c
    "11101110", --  269 - 0x10d  :  238 - 0xee
    "11000110", --  270 - 0x10e  :  198 - 0xc6
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "01100110", --  272 - 0x110  :  102 - 0x66 -- Background 0x22
    "01100110", --  273 - 0x111  :  102 - 0x66
    "01100110", --  274 - 0x112  :  102 - 0x66
    "00111100", --  275 - 0x113  :   60 - 0x3c
    "00011000", --  276 - 0x114  :   24 - 0x18
    "00011000", --  277 - 0x115  :   24 - 0x18
    "00011000", --  278 - 0x116  :   24 - 0x18
    "00000000", --  279 - 0x117  :    0 - 0x0
    "11111110", --  280 - 0x118  :  254 - 0xfe -- Background 0x23
    "00001110", --  281 - 0x119  :   14 - 0xe
    "00011100", --  282 - 0x11a  :   28 - 0x1c
    "00111000", --  283 - 0x11b  :   56 - 0x38
    "01110000", --  284 - 0x11c  :  112 - 0x70
    "11100000", --  285 - 0x11d  :  224 - 0xe0
    "11111110", --  286 - 0x11e  :  254 - 0xfe
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "11111111", --  296 - 0x128  :  255 - 0xff -- Background 0x25
    "11111111", --  297 - 0x129  :  255 - 0xff
    "11111111", --  298 - 0x12a  :  255 - 0xff
    "11111111", --  299 - 0x12b  :  255 - 0xff
    "11111111", --  300 - 0x12c  :  255 - 0xff
    "11111111", --  301 - 0x12d  :  255 - 0xff
    "11111111", --  302 - 0x12e  :  255 - 0xff
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Background 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "11111111", --  312 - 0x138  :  255 - 0xff -- Background 0x27
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11111111", --  316 - 0x13c  :  255 - 0xff
    "11111111", --  317 - 0x13d  :  255 - 0xff
    "11111111", --  318 - 0x13e  :  255 - 0xff
    "11111111", --  319 - 0x13f  :  255 - 0xff
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "01111110", --  323 - 0x143  :  126 - 0x7e
    "01111110", --  324 - 0x144  :  126 - 0x7e
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Background 0x29
    "00000000", --  329 - 0x149  :    0 - 0x0
    "01000100", --  330 - 0x14a  :   68 - 0x44
    "00101000", --  331 - 0x14b  :   40 - 0x28
    "00010000", --  332 - 0x14c  :   16 - 0x10
    "00101000", --  333 - 0x14d  :   40 - 0x28
    "01000100", --  334 - 0x14e  :   68 - 0x44
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "11111111", --  336 - 0x150  :  255 - 0xff -- Background 0x2a
    "11111111", --  337 - 0x151  :  255 - 0xff
    "11111111", --  338 - 0x152  :  255 - 0xff
    "11111111", --  339 - 0x153  :  255 - 0xff
    "11111111", --  340 - 0x154  :  255 - 0xff
    "11111111", --  341 - 0x155  :  255 - 0xff
    "11111111", --  342 - 0x156  :  255 - 0xff
    "11111111", --  343 - 0x157  :  255 - 0xff
    "00011000", --  344 - 0x158  :   24 - 0x18 -- Background 0x2b
    "00111100", --  345 - 0x159  :   60 - 0x3c
    "00111100", --  346 - 0x15a  :   60 - 0x3c
    "00111100", --  347 - 0x15b  :   60 - 0x3c
    "00011000", --  348 - 0x15c  :   24 - 0x18
    "00011000", --  349 - 0x15d  :   24 - 0x18
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00011000", --  351 - 0x15f  :   24 - 0x18
    "11111111", --  352 - 0x160  :  255 - 0xff -- Background 0x2c
    "01111111", --  353 - 0x161  :  127 - 0x7f
    "01111111", --  354 - 0x162  :  127 - 0x7f
    "01111111", --  355 - 0x163  :  127 - 0x7f
    "01111111", --  356 - 0x164  :  127 - 0x7f
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11100011", --  358 - 0x166  :  227 - 0xe3
    "11000001", --  359 - 0x167  :  193 - 0xc1
    "10000000", --  360 - 0x168  :  128 - 0x80 -- Background 0x2d
    "10000000", --  361 - 0x169  :  128 - 0x80
    "10000000", --  362 - 0x16a  :  128 - 0x80
    "11000001", --  363 - 0x16b  :  193 - 0xc1
    "11100011", --  364 - 0x16c  :  227 - 0xe3
    "11111111", --  365 - 0x16d  :  255 - 0xff
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "00111000", --  368 - 0x170  :   56 - 0x38 -- Background 0x2e
    "01111100", --  369 - 0x171  :  124 - 0x7c
    "01111100", --  370 - 0x172  :  124 - 0x7c
    "01111100", --  371 - 0x173  :  124 - 0x7c
    "01111100", --  372 - 0x174  :  124 - 0x7c
    "01111100", --  373 - 0x175  :  124 - 0x7c
    "00111000", --  374 - 0x176  :   56 - 0x38
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000011", --  376 - 0x178  :    3 - 0x3 -- Background 0x2f
    "00000110", --  377 - 0x179  :    6 - 0x6
    "00001100", --  378 - 0x17a  :   12 - 0xc
    "00001100", --  379 - 0x17b  :   12 - 0xc
    "00001000", --  380 - 0x17c  :    8 - 0x8
    "00001000", --  381 - 0x17d  :    8 - 0x8
    "00000100", --  382 - 0x17e  :    4 - 0x4
    "00000011", --  383 - 0x17f  :    3 - 0x3
    "00000001", --  384 - 0x180  :    1 - 0x1 -- Background 0x30
    "00000010", --  385 - 0x181  :    2 - 0x2
    "00000100", --  386 - 0x182  :    4 - 0x4
    "00001000", --  387 - 0x183  :    8 - 0x8
    "00010000", --  388 - 0x184  :   16 - 0x10
    "00100000", --  389 - 0x185  :   32 - 0x20
    "01000000", --  390 - 0x186  :   64 - 0x40
    "10000000", --  391 - 0x187  :  128 - 0x80
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Background 0x31
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000111", --  397 - 0x18d  :    7 - 0x7
    "00111000", --  398 - 0x18e  :   56 - 0x38
    "11000000", --  399 - 0x18f  :  192 - 0xc0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Background 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "11100000", --  405 - 0x195  :  224 - 0xe0
    "00011100", --  406 - 0x196  :   28 - 0x1c
    "00000011", --  407 - 0x197  :    3 - 0x3
    "10000000", --  408 - 0x198  :  128 - 0x80 -- Background 0x33
    "01000000", --  409 - 0x199  :   64 - 0x40
    "00100000", --  410 - 0x19a  :   32 - 0x20
    "00010000", --  411 - 0x19b  :   16 - 0x10
    "00001000", --  412 - 0x19c  :    8 - 0x8
    "00000100", --  413 - 0x19d  :    4 - 0x4
    "00000010", --  414 - 0x19e  :    2 - 0x2
    "00000001", --  415 - 0x19f  :    1 - 0x1
    "00000100", --  416 - 0x1a0  :    4 - 0x4 -- Background 0x34
    "00001110", --  417 - 0x1a1  :   14 - 0xe
    "00001110", --  418 - 0x1a2  :   14 - 0xe
    "00001110", --  419 - 0x1a3  :   14 - 0xe
    "01101110", --  420 - 0x1a4  :  110 - 0x6e
    "01100100", --  421 - 0x1a5  :  100 - 0x64
    "01100000", --  422 - 0x1a6  :   96 - 0x60
    "01100000", --  423 - 0x1a7  :   96 - 0x60
    "00000111", --  424 - 0x1a8  :    7 - 0x7 -- Background 0x35
    "00001111", --  425 - 0x1a9  :   15 - 0xf
    "00011111", --  426 - 0x1aa  :   31 - 0x1f
    "00011111", --  427 - 0x1ab  :   31 - 0x1f
    "01111111", --  428 - 0x1ac  :  127 - 0x7f
    "11111111", --  429 - 0x1ad  :  255 - 0xff
    "11111111", --  430 - 0x1ae  :  255 - 0xff
    "01111111", --  431 - 0x1af  :  127 - 0x7f
    "00000011", --  432 - 0x1b0  :    3 - 0x3 -- Background 0x36
    "00000111", --  433 - 0x1b1  :    7 - 0x7
    "00011111", --  434 - 0x1b2  :   31 - 0x1f
    "00111111", --  435 - 0x1b3  :   63 - 0x3f
    "00111111", --  436 - 0x1b4  :   63 - 0x3f
    "00111111", --  437 - 0x1b5  :   63 - 0x3f
    "01111001", --  438 - 0x1b6  :  121 - 0x79
    "11110111", --  439 - 0x1b7  :  247 - 0xf7
    "11000000", --  440 - 0x1b8  :  192 - 0xc0 -- Background 0x37
    "11100000", --  441 - 0x1b9  :  224 - 0xe0
    "11110000", --  442 - 0x1ba  :  240 - 0xf0
    "11110100", --  443 - 0x1bb  :  244 - 0xf4
    "11111110", --  444 - 0x1bc  :  254 - 0xfe
    "10111111", --  445 - 0x1bd  :  191 - 0xbf
    "11011111", --  446 - 0x1be  :  223 - 0xdf
    "11111111", --  447 - 0x1bf  :  255 - 0xff
    "10010000", --  448 - 0x1c0  :  144 - 0x90 -- Background 0x38
    "10111000", --  449 - 0x1c1  :  184 - 0xb8
    "11111000", --  450 - 0x1c2  :  248 - 0xf8
    "11111010", --  451 - 0x1c3  :  250 - 0xfa
    "11111111", --  452 - 0x1c4  :  255 - 0xff
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11111111", --  454 - 0x1c6  :  255 - 0xff
    "11111110", --  455 - 0x1c7  :  254 - 0xfe
    "00111011", --  456 - 0x1c8  :   59 - 0x3b -- Background 0x39
    "00011101", --  457 - 0x1c9  :   29 - 0x1d
    "00001110", --  458 - 0x1ca  :   14 - 0xe
    "00001111", --  459 - 0x1cb  :   15 - 0xf
    "00000111", --  460 - 0x1cc  :    7 - 0x7
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "11111111", --  464 - 0x1d0  :  255 - 0xff -- Background 0x3a
    "10111111", --  465 - 0x1d1  :  191 - 0xbf
    "00011100", --  466 - 0x1d2  :   28 - 0x1c
    "11000000", --  467 - 0x1d3  :  192 - 0xc0
    "11110011", --  468 - 0x1d4  :  243 - 0xf3
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "01111110", --  470 - 0x1d6  :  126 - 0x7e
    "00011100", --  471 - 0x1d7  :   28 - 0x1c
    "10111111", --  472 - 0x1d8  :  191 - 0xbf -- Background 0x3b
    "01111111", --  473 - 0x1d9  :  127 - 0x7f
    "00111101", --  474 - 0x1da  :   61 - 0x3d
    "10000011", --  475 - 0x1db  :  131 - 0x83
    "11000111", --  476 - 0x1dc  :  199 - 0xc7
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11111111", --  478 - 0x1de  :  255 - 0xff
    "00111100", --  479 - 0x1df  :   60 - 0x3c
    "11111100", --  480 - 0x1e0  :  252 - 0xfc -- Background 0x3c
    "11111110", --  481 - 0x1e1  :  254 - 0xfe
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111110", --  483 - 0x1e3  :  254 - 0xfe
    "11111110", --  484 - 0x1e4  :  254 - 0xfe
    "11111000", --  485 - 0x1e5  :  248 - 0xf8
    "01100000", --  486 - 0x1e6  :   96 - 0x60
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "11000000", --  488 - 0x1e8  :  192 - 0xc0 -- Background 0x3d
    "00100000", --  489 - 0x1e9  :   32 - 0x20
    "00010000", --  490 - 0x1ea  :   16 - 0x10
    "00010000", --  491 - 0x1eb  :   16 - 0x10
    "00010000", --  492 - 0x1ec  :   16 - 0x10
    "00010000", --  493 - 0x1ed  :   16 - 0x10
    "00100000", --  494 - 0x1ee  :   32 - 0x20
    "11000000", --  495 - 0x1ef  :  192 - 0xc0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "01111111", --  501 - 0x1f5  :  127 - 0x7f
    "11100000", --  502 - 0x1f6  :  224 - 0xe0
    "11000000", --  503 - 0x1f7  :  192 - 0xc0
    "10001000", --  504 - 0x1f8  :  136 - 0x88 -- Background 0x3f
    "10011100", --  505 - 0x1f9  :  156 - 0x9c
    "10001000", --  506 - 0x1fa  :  136 - 0x88
    "10000000", --  507 - 0x1fb  :  128 - 0x80
    "10000000", --  508 - 0x1fc  :  128 - 0x80
    "10000000", --  509 - 0x1fd  :  128 - 0x80
    "10000000", --  510 - 0x1fe  :  128 - 0x80
    "10000000", --  511 - 0x1ff  :  128 - 0x80
    "11111110", --  512 - 0x200  :  254 - 0xfe -- Background 0x40
    "11111110", --  513 - 0x201  :  254 - 0xfe
    "11111110", --  514 - 0x202  :  254 - 0xfe
    "11111110", --  515 - 0x203  :  254 - 0xfe
    "11111110", --  516 - 0x204  :  254 - 0xfe
    "11111110", --  517 - 0x205  :  254 - 0xfe
    "11111110", --  518 - 0x206  :  254 - 0xfe
    "11111110", --  519 - 0x207  :  254 - 0xfe
    "00001000", --  520 - 0x208  :    8 - 0x8 -- Background 0x41
    "00010100", --  521 - 0x209  :   20 - 0x14
    "00100100", --  522 - 0x20a  :   36 - 0x24
    "11000100", --  523 - 0x20b  :  196 - 0xc4
    "00000011", --  524 - 0x20c  :    3 - 0x3
    "01000000", --  525 - 0x20d  :   64 - 0x40
    "10100001", --  526 - 0x20e  :  161 - 0xa1
    "00100110", --  527 - 0x20f  :   38 - 0x26
    "11111111", --  528 - 0x210  :  255 - 0xff -- Background 0x42
    "11111111", --  529 - 0x211  :  255 - 0xff
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11111111", --  531 - 0x213  :  255 - 0xff
    "01111111", --  532 - 0x214  :  127 - 0x7f
    "01111111", --  533 - 0x215  :  127 - 0x7f
    "01111111", --  534 - 0x216  :  127 - 0x7f
    "01111111", --  535 - 0x217  :  127 - 0x7f
    "11111111", --  536 - 0x218  :  255 - 0xff -- Background 0x43
    "11111111", --  537 - 0x219  :  255 - 0xff
    "11111111", --  538 - 0x21a  :  255 - 0xff
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11111111", --  542 - 0x21e  :  255 - 0xff
    "11111111", --  543 - 0x21f  :  255 - 0xff
    "01111111", --  544 - 0x220  :  127 - 0x7f -- Background 0x44
    "10000000", --  545 - 0x221  :  128 - 0x80
    "10000000", --  546 - 0x222  :  128 - 0x80
    "10011000", --  547 - 0x223  :  152 - 0x98
    "10011100", --  548 - 0x224  :  156 - 0x9c
    "10001100", --  549 - 0x225  :  140 - 0x8c
    "10000000", --  550 - 0x226  :  128 - 0x80
    "10000000", --  551 - 0x227  :  128 - 0x80
    "11111111", --  552 - 0x228  :  255 - 0xff -- Background 0x45
    "00000001", --  553 - 0x229  :    1 - 0x1
    "00000001", --  554 - 0x22a  :    1 - 0x1
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "00010000", --  556 - 0x22c  :   16 - 0x10
    "00010000", --  557 - 0x22d  :   16 - 0x10
    "00010000", --  558 - 0x22e  :   16 - 0x10
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "10000000", --  560 - 0x230  :  128 - 0x80 -- Background 0x46
    "10000000", --  561 - 0x231  :  128 - 0x80
    "10000000", --  562 - 0x232  :  128 - 0x80
    "10000000", --  563 - 0x233  :  128 - 0x80
    "10000000", --  564 - 0x234  :  128 - 0x80
    "10000000", --  565 - 0x235  :  128 - 0x80
    "10000000", --  566 - 0x236  :  128 - 0x80
    "10000000", --  567 - 0x237  :  128 - 0x80
    "00000001", --  568 - 0x238  :    1 - 0x1 -- Background 0x47
    "00000001", --  569 - 0x239  :    1 - 0x1
    "00000001", --  570 - 0x23a  :    1 - 0x1
    "11111111", --  571 - 0x23b  :  255 - 0xff
    "00010000", --  572 - 0x23c  :   16 - 0x10
    "00010000", --  573 - 0x23d  :   16 - 0x10
    "00010000", --  574 - 0x23e  :   16 - 0x10
    "11111111", --  575 - 0x23f  :  255 - 0xff
    "11111111", --  576 - 0x240  :  255 - 0xff -- Background 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "11111110", --  584 - 0x248  :  254 - 0xfe -- Background 0x49
    "00000001", --  585 - 0x249  :    1 - 0x1
    "00000001", --  586 - 0x24a  :    1 - 0x1
    "00011001", --  587 - 0x24b  :   25 - 0x19
    "00011101", --  588 - 0x24c  :   29 - 0x1d
    "00001101", --  589 - 0x24d  :   13 - 0xd
    "00000001", --  590 - 0x24e  :    1 - 0x1
    "00000001", --  591 - 0x24f  :    1 - 0x1
    "00000001", --  592 - 0x250  :    1 - 0x1 -- Background 0x4a
    "00000001", --  593 - 0x251  :    1 - 0x1
    "00000001", --  594 - 0x252  :    1 - 0x1
    "00000001", --  595 - 0x253  :    1 - 0x1
    "00000001", --  596 - 0x254  :    1 - 0x1
    "00000001", --  597 - 0x255  :    1 - 0x1
    "00000001", --  598 - 0x256  :    1 - 0x1
    "00000001", --  599 - 0x257  :    1 - 0x1
    "00111111", --  600 - 0x258  :   63 - 0x3f -- Background 0x4b
    "01111111", --  601 - 0x259  :  127 - 0x7f
    "01111111", --  602 - 0x25a  :  127 - 0x7f
    "11111111", --  603 - 0x25b  :  255 - 0xff
    "11111111", --  604 - 0x25c  :  255 - 0xff
    "11111111", --  605 - 0x25d  :  255 - 0xff
    "11111111", --  606 - 0x25e  :  255 - 0xff
    "11111111", --  607 - 0x25f  :  255 - 0xff
    "11111111", --  608 - 0x260  :  255 - 0xff -- Background 0x4c
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "01111110", --  614 - 0x266  :  126 - 0x7e
    "00111100", --  615 - 0x267  :   60 - 0x3c
    "11111111", --  616 - 0x268  :  255 - 0xff -- Background 0x4d
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11111111", --  620 - 0x26c  :  255 - 0xff
    "11111111", --  621 - 0x26d  :  255 - 0xff
    "11111111", --  622 - 0x26e  :  255 - 0xff
    "11111111", --  623 - 0x26f  :  255 - 0xff
    "11111111", --  624 - 0x270  :  255 - 0xff -- Background 0x4e
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11111111", --  626 - 0x272  :  255 - 0xff
    "11111111", --  627 - 0x273  :  255 - 0xff
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111111", --  629 - 0x275  :  255 - 0xff
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "11111111", --  632 - 0x278  :  255 - 0xff -- Background 0x4f
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11111111", --  634 - 0x27a  :  255 - 0xff
    "11111111", --  635 - 0x27b  :  255 - 0xff
    "11111111", --  636 - 0x27c  :  255 - 0xff
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11111110", --  638 - 0x27e  :  254 - 0xfe
    "01111100", --  639 - 0x27f  :  124 - 0x7c
    "11111000", --  640 - 0x280  :  248 - 0xf8 -- Background 0x50
    "11111100", --  641 - 0x281  :  252 - 0xfc
    "11111110", --  642 - 0x282  :  254 - 0xfe
    "11111110", --  643 - 0x283  :  254 - 0xfe
    "11111111", --  644 - 0x284  :  255 - 0xff
    "11111111", --  645 - 0x285  :  255 - 0xff
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111111", --  648 - 0x288  :  255 - 0xff -- Background 0x51
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11111111", --  650 - 0x28a  :  255 - 0xff
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "11111111", --  652 - 0x28c  :  255 - 0xff
    "11111111", --  653 - 0x28d  :  255 - 0xff
    "01111110", --  654 - 0x28e  :  126 - 0x7e
    "00111100", --  655 - 0x28f  :   60 - 0x3c
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x52
    "00001000", --  657 - 0x291  :    8 - 0x8
    "00001000", --  658 - 0x292  :    8 - 0x8
    "00001000", --  659 - 0x293  :    8 - 0x8
    "00010000", --  660 - 0x294  :   16 - 0x10
    "00010000", --  661 - 0x295  :   16 - 0x10
    "00010000", --  662 - 0x296  :   16 - 0x10
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Background 0x53
    "01111111", --  665 - 0x299  :  127 - 0x7f
    "01111111", --  666 - 0x29a  :  127 - 0x7f
    "01111000", --  667 - 0x29b  :  120 - 0x78
    "01110011", --  668 - 0x29c  :  115 - 0x73
    "01110011", --  669 - 0x29d  :  115 - 0x73
    "01110011", --  670 - 0x29e  :  115 - 0x73
    "01111111", --  671 - 0x29f  :  127 - 0x7f
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Background 0x54
    "11111111", --  673 - 0x2a1  :  255 - 0xff
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "00111111", --  675 - 0x2a3  :   63 - 0x3f
    "10011111", --  676 - 0x2a4  :  159 - 0x9f
    "10011111", --  677 - 0x2a5  :  159 - 0x9f
    "10011111", --  678 - 0x2a6  :  159 - 0x9f
    "00011111", --  679 - 0x2a7  :   31 - 0x1f
    "01111110", --  680 - 0x2a8  :  126 - 0x7e -- Background 0x55
    "01111110", --  681 - 0x2a9  :  126 - 0x7e
    "01111111", --  682 - 0x2aa  :  127 - 0x7f
    "01111110", --  683 - 0x2ab  :  126 - 0x7e
    "01111110", --  684 - 0x2ac  :  126 - 0x7e
    "01111111", --  685 - 0x2ad  :  127 - 0x7f
    "01111111", --  686 - 0x2ae  :  127 - 0x7f
    "11111111", --  687 - 0x2af  :  255 - 0xff
    "01111111", --  688 - 0x2b0  :  127 - 0x7f -- Background 0x56
    "01111111", --  689 - 0x2b1  :  127 - 0x7f
    "11111111", --  690 - 0x2b2  :  255 - 0xff
    "01111111", --  691 - 0x2b3  :  127 - 0x7f
    "01111111", --  692 - 0x2b4  :  127 - 0x7f
    "11111111", --  693 - 0x2b5  :  255 - 0xff
    "11111111", --  694 - 0x2b6  :  255 - 0xff
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "01111111", --  696 - 0x2b8  :  127 - 0x7f -- Background 0x57
    "10000000", --  697 - 0x2b9  :  128 - 0x80
    "10100000", --  698 - 0x2ba  :  160 - 0xa0
    "10000000", --  699 - 0x2bb  :  128 - 0x80
    "10000000", --  700 - 0x2bc  :  128 - 0x80
    "10000000", --  701 - 0x2bd  :  128 - 0x80
    "10000000", --  702 - 0x2be  :  128 - 0x80
    "10000000", --  703 - 0x2bf  :  128 - 0x80
    "11111110", --  704 - 0x2c0  :  254 - 0xfe -- Background 0x58
    "00000001", --  705 - 0x2c1  :    1 - 0x1
    "00000101", --  706 - 0x2c2  :    5 - 0x5
    "00000001", --  707 - 0x2c3  :    1 - 0x1
    "00000001", --  708 - 0x2c4  :    1 - 0x1
    "00000001", --  709 - 0x2c5  :    1 - 0x1
    "00000001", --  710 - 0x2c6  :    1 - 0x1
    "00000001", --  711 - 0x2c7  :    1 - 0x1
    "10000000", --  712 - 0x2c8  :  128 - 0x80 -- Background 0x59
    "10000000", --  713 - 0x2c9  :  128 - 0x80
    "10000000", --  714 - 0x2ca  :  128 - 0x80
    "10000000", --  715 - 0x2cb  :  128 - 0x80
    "10000000", --  716 - 0x2cc  :  128 - 0x80
    "10100000", --  717 - 0x2cd  :  160 - 0xa0
    "10000000", --  718 - 0x2ce  :  128 - 0x80
    "01111111", --  719 - 0x2cf  :  127 - 0x7f
    "00000001", --  720 - 0x2d0  :    1 - 0x1 -- Background 0x5a
    "00000001", --  721 - 0x2d1  :    1 - 0x1
    "00000001", --  722 - 0x2d2  :    1 - 0x1
    "00000001", --  723 - 0x2d3  :    1 - 0x1
    "00000001", --  724 - 0x2d4  :    1 - 0x1
    "00000101", --  725 - 0x2d5  :    5 - 0x5
    "00000001", --  726 - 0x2d6  :    1 - 0x1
    "11111110", --  727 - 0x2d7  :  254 - 0xfe
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "11111100", --  732 - 0x2dc  :  252 - 0xfc
    "11111110", --  733 - 0x2dd  :  254 - 0xfe
    "00000111", --  734 - 0x2de  :    7 - 0x7
    "00000011", --  735 - 0x2df  :    3 - 0x3
    "00010001", --  736 - 0x2e0  :   17 - 0x11 -- Background 0x5c
    "00111001", --  737 - 0x2e1  :   57 - 0x39
    "00010001", --  738 - 0x2e2  :   17 - 0x11
    "00000001", --  739 - 0x2e3  :    1 - 0x1
    "00000001", --  740 - 0x2e4  :    1 - 0x1
    "00000001", --  741 - 0x2e5  :    1 - 0x1
    "00000001", --  742 - 0x2e6  :    1 - 0x1
    "00000001", --  743 - 0x2e7  :    1 - 0x1
    "11101111", --  744 - 0x2e8  :  239 - 0xef -- Background 0x5d
    "00101000", --  745 - 0x2e9  :   40 - 0x28
    "00101000", --  746 - 0x2ea  :   40 - 0x28
    "00101000", --  747 - 0x2eb  :   40 - 0x28
    "00101000", --  748 - 0x2ec  :   40 - 0x28
    "00101000", --  749 - 0x2ed  :   40 - 0x28
    "11101111", --  750 - 0x2ee  :  239 - 0xef
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "11111110", --  752 - 0x2f0  :  254 - 0xfe -- Background 0x5e
    "10000010", --  753 - 0x2f1  :  130 - 0x82
    "10000010", --  754 - 0x2f2  :  130 - 0x82
    "10000010", --  755 - 0x2f3  :  130 - 0x82
    "10000010", --  756 - 0x2f4  :  130 - 0x82
    "10000010", --  757 - 0x2f5  :  130 - 0x82
    "11111110", --  758 - 0x2f6  :  254 - 0xfe
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "10000000", --  760 - 0x2f8  :  128 - 0x80 -- Background 0x5f
    "10000000", --  761 - 0x2f9  :  128 - 0x80
    "10000000", --  762 - 0x2fa  :  128 - 0x80
    "10011000", --  763 - 0x2fb  :  152 - 0x98
    "10011100", --  764 - 0x2fc  :  156 - 0x9c
    "10001100", --  765 - 0x2fd  :  140 - 0x8c
    "10000000", --  766 - 0x2fe  :  128 - 0x80
    "01111111", --  767 - 0x2ff  :  127 - 0x7f
    "11111111", --  768 - 0x300  :  255 - 0xff -- Background 0x60
    "11111111", --  769 - 0x301  :  255 - 0xff
    "10000011", --  770 - 0x302  :  131 - 0x83
    "11110011", --  771 - 0x303  :  243 - 0xf3
    "11110011", --  772 - 0x304  :  243 - 0xf3
    "11110011", --  773 - 0x305  :  243 - 0xf3
    "11110011", --  774 - 0x306  :  243 - 0xf3
    "11110011", --  775 - 0x307  :  243 - 0xf3
    "11111111", --  776 - 0x308  :  255 - 0xff -- Background 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11110000", --  778 - 0x30a  :  240 - 0xf0
    "11110110", --  779 - 0x30b  :  246 - 0xf6
    "11110110", --  780 - 0x30c  :  246 - 0xf6
    "11110110", --  781 - 0x30d  :  246 - 0xf6
    "11110110", --  782 - 0x30e  :  246 - 0xf6
    "11110110", --  783 - 0x30f  :  246 - 0xf6
    "11111111", --  784 - 0x310  :  255 - 0xff -- Background 0x62
    "11111111", --  785 - 0x311  :  255 - 0xff
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "11111111", --  792 - 0x318  :  255 - 0xff -- Background 0x63
    "11111111", --  793 - 0x319  :  255 - 0xff
    "00000001", --  794 - 0x31a  :    1 - 0x1
    "01010111", --  795 - 0x31b  :   87 - 0x57
    "00101111", --  796 - 0x31c  :   47 - 0x2f
    "01010111", --  797 - 0x31d  :   87 - 0x57
    "00101111", --  798 - 0x31e  :   47 - 0x2f
    "01010111", --  799 - 0x31f  :   87 - 0x57
    "11110011", --  800 - 0x320  :  243 - 0xf3 -- Background 0x64
    "11110011", --  801 - 0x321  :  243 - 0xf3
    "11110011", --  802 - 0x322  :  243 - 0xf3
    "11110011", --  803 - 0x323  :  243 - 0xf3
    "11110011", --  804 - 0x324  :  243 - 0xf3
    "11110011", --  805 - 0x325  :  243 - 0xf3
    "11111111", --  806 - 0x326  :  255 - 0xff
    "00111111", --  807 - 0x327  :   63 - 0x3f
    "11110110", --  808 - 0x328  :  246 - 0xf6 -- Background 0x65
    "11110110", --  809 - 0x329  :  246 - 0xf6
    "11110110", --  810 - 0x32a  :  246 - 0xf6
    "11110110", --  811 - 0x32b  :  246 - 0xf6
    "11110110", --  812 - 0x32c  :  246 - 0xf6
    "11110110", --  813 - 0x32d  :  246 - 0xf6
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Background 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111111", --  823 - 0x337  :  255 - 0xff
    "00101111", --  824 - 0x338  :   47 - 0x2f -- Background 0x67
    "01010111", --  825 - 0x339  :   87 - 0x57
    "00101111", --  826 - 0x33a  :   47 - 0x2f
    "01010111", --  827 - 0x33b  :   87 - 0x57
    "00101111", --  828 - 0x33c  :   47 - 0x2f
    "01010111", --  829 - 0x33d  :   87 - 0x57
    "11111111", --  830 - 0x33e  :  255 - 0xff
    "11111100", --  831 - 0x33f  :  252 - 0xfc
    "00111100", --  832 - 0x340  :   60 - 0x3c -- Background 0x68
    "00111100", --  833 - 0x341  :   60 - 0x3c
    "00111100", --  834 - 0x342  :   60 - 0x3c
    "00111100", --  835 - 0x343  :   60 - 0x3c
    "00111100", --  836 - 0x344  :   60 - 0x3c
    "00111100", --  837 - 0x345  :   60 - 0x3c
    "00111100", --  838 - 0x346  :   60 - 0x3c
    "00111100", --  839 - 0x347  :   60 - 0x3c
    "11111011", --  840 - 0x348  :  251 - 0xfb -- Background 0x69
    "11111011", --  841 - 0x349  :  251 - 0xfb
    "11111011", --  842 - 0x34a  :  251 - 0xfb
    "11111011", --  843 - 0x34b  :  251 - 0xfb
    "11111011", --  844 - 0x34c  :  251 - 0xfb
    "11111011", --  845 - 0x34d  :  251 - 0xfb
    "11111011", --  846 - 0x34e  :  251 - 0xfb
    "11111011", --  847 - 0x34f  :  251 - 0xfb
    "10111100", --  848 - 0x350  :  188 - 0xbc -- Background 0x6a
    "01011100", --  849 - 0x351  :   92 - 0x5c
    "10111100", --  850 - 0x352  :  188 - 0xbc
    "01011100", --  851 - 0x353  :   92 - 0x5c
    "10111100", --  852 - 0x354  :  188 - 0xbc
    "01011100", --  853 - 0x355  :   92 - 0x5c
    "10111100", --  854 - 0x356  :  188 - 0xbc
    "01011100", --  855 - 0x357  :   92 - 0x5c
    "00011111", --  856 - 0x358  :   31 - 0x1f -- Background 0x6b
    "00100000", --  857 - 0x359  :   32 - 0x20
    "01000000", --  858 - 0x35a  :   64 - 0x40
    "01000000", --  859 - 0x35b  :   64 - 0x40
    "10000000", --  860 - 0x35c  :  128 - 0x80
    "10000000", --  861 - 0x35d  :  128 - 0x80
    "10000000", --  862 - 0x35e  :  128 - 0x80
    "10000001", --  863 - 0x35f  :  129 - 0x81
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x6c
    "10000000", --  865 - 0x361  :  128 - 0x80
    "10000000", --  866 - 0x362  :  128 - 0x80
    "11000000", --  867 - 0x363  :  192 - 0xc0
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111110", --  870 - 0x366  :  254 - 0xfe
    "11111110", --  871 - 0x367  :  254 - 0xfe
    "11111111", --  872 - 0x368  :  255 - 0xff -- Background 0x6d
    "01111111", --  873 - 0x369  :  127 - 0x7f
    "01111111", --  874 - 0x36a  :  127 - 0x7f
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "00000111", --  877 - 0x36d  :    7 - 0x7
    "00000011", --  878 - 0x36e  :    3 - 0x3
    "00000011", --  879 - 0x36f  :    3 - 0x3
    "11111111", --  880 - 0x370  :  255 - 0xff -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "10000001", --  885 - 0x375  :  129 - 0x81
    "11000011", --  886 - 0x376  :  195 - 0xc3
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111000", --  888 - 0x378  :  248 - 0xf8 -- Background 0x6f
    "11111100", --  889 - 0x379  :  252 - 0xfc
    "11111110", --  890 - 0x37a  :  254 - 0xfe
    "11111110", --  891 - 0x37b  :  254 - 0xfe
    "11100011", --  892 - 0x37c  :  227 - 0xe3
    "11000001", --  893 - 0x37d  :  193 - 0xc1
    "10000001", --  894 - 0x37e  :  129 - 0x81
    "10000001", --  895 - 0x37f  :  129 - 0x81
    "10000011", --  896 - 0x380  :  131 - 0x83 -- Background 0x70
    "11111111", --  897 - 0x381  :  255 - 0xff
    "11111111", --  898 - 0x382  :  255 - 0xff
    "11111111", --  899 - 0x383  :  255 - 0xff
    "11111111", --  900 - 0x384  :  255 - 0xff
    "11111111", --  901 - 0x385  :  255 - 0xff
    "01111111", --  902 - 0x386  :  127 - 0x7f
    "00011111", --  903 - 0x387  :   31 - 0x1f
    "11111100", --  904 - 0x388  :  252 - 0xfc -- Background 0x71
    "11111100", --  905 - 0x389  :  252 - 0xfc
    "11111100", --  906 - 0x38a  :  252 - 0xfc
    "11111100", --  907 - 0x38b  :  252 - 0xfc
    "11111110", --  908 - 0x38c  :  254 - 0xfe
    "11111110", --  909 - 0x38d  :  254 - 0xfe
    "11111111", --  910 - 0x38e  :  255 - 0xff
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "00000001", --  912 - 0x390  :    1 - 0x1 -- Background 0x72
    "00000001", --  913 - 0x391  :    1 - 0x1
    "00000001", --  914 - 0x392  :    1 - 0x1
    "00000001", --  915 - 0x393  :    1 - 0x1
    "00000011", --  916 - 0x394  :    3 - 0x3
    "00000011", --  917 - 0x395  :    3 - 0x3
    "00000111", --  918 - 0x396  :    7 - 0x7
    "11111111", --  919 - 0x397  :  255 - 0xff
    "11111111", --  920 - 0x398  :  255 - 0xff -- Background 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111111", --  927 - 0x39f  :  255 - 0xff
    "10000001", --  928 - 0x3a0  :  129 - 0x81 -- Background 0x74
    "11000001", --  929 - 0x3a1  :  193 - 0xc1
    "11100011", --  930 - 0x3a2  :  227 - 0xe3
    "11111111", --  931 - 0x3a3  :  255 - 0xff
    "11111111", --  932 - 0x3a4  :  255 - 0xff
    "11111111", --  933 - 0x3a5  :  255 - 0xff
    "11111111", --  934 - 0x3a6  :  255 - 0xff
    "11111110", --  935 - 0x3a7  :  254 - 0xfe
    "11111111", --  936 - 0x3a8  :  255 - 0xff -- Background 0x75
    "11111111", --  937 - 0x3a9  :  255 - 0xff
    "11111111", --  938 - 0x3aa  :  255 - 0xff
    "11111111", --  939 - 0x3ab  :  255 - 0xff
    "11111111", --  940 - 0x3ac  :  255 - 0xff
    "11111011", --  941 - 0x3ad  :  251 - 0xfb
    "10110101", --  942 - 0x3ae  :  181 - 0xb5
    "11001110", --  943 - 0x3af  :  206 - 0xce
    "11111111", --  944 - 0x3b0  :  255 - 0xff -- Background 0x76
    "11111111", --  945 - 0x3b1  :  255 - 0xff
    "11111111", --  946 - 0x3b2  :  255 - 0xff
    "11111111", --  947 - 0x3b3  :  255 - 0xff
    "11111111", --  948 - 0x3b4  :  255 - 0xff
    "11011111", --  949 - 0x3b5  :  223 - 0xdf
    "10101101", --  950 - 0x3b6  :  173 - 0xad
    "01110011", --  951 - 0x3b7  :  115 - 0x73
    "01110111", --  952 - 0x3b8  :  119 - 0x77 -- Background 0x77
    "01110111", --  953 - 0x3b9  :  119 - 0x77
    "01110111", --  954 - 0x3ba  :  119 - 0x77
    "01110111", --  955 - 0x3bb  :  119 - 0x77
    "01110111", --  956 - 0x3bc  :  119 - 0x77
    "01110111", --  957 - 0x3bd  :  119 - 0x77
    "01110111", --  958 - 0x3be  :  119 - 0x77
    "01110111", --  959 - 0x3bf  :  119 - 0x77
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "01110111", --  968 - 0x3c8  :  119 - 0x77 -- Background 0x79
    "01110111", --  969 - 0x3c9  :  119 - 0x77
    "01110111", --  970 - 0x3ca  :  119 - 0x77
    "01110111", --  971 - 0x3cb  :  119 - 0x77
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000001", --  976 - 0x3d0  :    1 - 0x1 -- Background 0x7a
    "00000001", --  977 - 0x3d1  :    1 - 0x1
    "00000001", --  978 - 0x3d2  :    1 - 0x1
    "00011001", --  979 - 0x3d3  :   25 - 0x19
    "00011101", --  980 - 0x3d4  :   29 - 0x1d
    "00001101", --  981 - 0x3d5  :   13 - 0xd
    "00000001", --  982 - 0x3d6  :    1 - 0x1
    "11111110", --  983 - 0x3d7  :  254 - 0xfe
    "00100000", --  984 - 0x3d8  :   32 - 0x20 -- Background 0x7b
    "01111000", --  985 - 0x3d9  :  120 - 0x78
    "01111111", --  986 - 0x3da  :  127 - 0x7f
    "11111110", --  987 - 0x3db  :  254 - 0xfe
    "11111110", --  988 - 0x3dc  :  254 - 0xfe
    "11111110", --  989 - 0x3dd  :  254 - 0xfe
    "11111110", --  990 - 0x3de  :  254 - 0xfe
    "11111110", --  991 - 0x3df  :  254 - 0xfe
    "00000100", --  992 - 0x3e0  :    4 - 0x4 -- Background 0x7c
    "10011010", --  993 - 0x3e1  :  154 - 0x9a
    "11111010", --  994 - 0x3e2  :  250 - 0xfa
    "11111101", --  995 - 0x3e3  :  253 - 0xfd
    "11111101", --  996 - 0x3e4  :  253 - 0xfd
    "11111101", --  997 - 0x3e5  :  253 - 0xfd
    "11111101", --  998 - 0x3e6  :  253 - 0xfd
    "11111101", --  999 - 0x3e7  :  253 - 0xfd
    "01111110", -- 1000 - 0x3e8  :  126 - 0x7e -- Background 0x7d
    "00111000", -- 1001 - 0x3e9  :   56 - 0x38
    "00100001", -- 1002 - 0x3ea  :   33 - 0x21
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000001", -- 1004 - 0x3ec  :    1 - 0x1
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000001", -- 1006 - 0x3ee  :    1 - 0x1
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "11111010", -- 1008 - 0x3f0  :  250 - 0xfa -- Background 0x7e
    "10001010", -- 1009 - 0x3f1  :  138 - 0x8a
    "10000100", -- 1010 - 0x3f2  :  132 - 0x84
    "10000000", -- 1011 - 0x3f3  :  128 - 0x80
    "10000000", -- 1012 - 0x3f4  :  128 - 0x80
    "10000000", -- 1013 - 0x3f5  :  128 - 0x80
    "10000000", -- 1014 - 0x3f6  :  128 - 0x80
    "10000000", -- 1015 - 0x3f7  :  128 - 0x80
    "00000010", -- 1016 - 0x3f8  :    2 - 0x2 -- Background 0x7f
    "00000100", -- 1017 - 0x3f9  :    4 - 0x4
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00010000", -- 1019 - 0x3fb  :   16 - 0x10
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "01000000", -- 1021 - 0x3fd  :   64 - 0x40
    "10000000", -- 1022 - 0x3fe  :  128 - 0x80
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00001011", -- 1024 - 0x400  :   11 - 0xb -- Background 0x80
    "00001011", -- 1025 - 0x401  :   11 - 0xb
    "00111011", -- 1026 - 0x402  :   59 - 0x3b
    "00001011", -- 1027 - 0x403  :   11 - 0xb
    "11111011", -- 1028 - 0x404  :  251 - 0xfb
    "00001011", -- 1029 - 0x405  :   11 - 0xb
    "00001011", -- 1030 - 0x406  :   11 - 0xb
    "00001010", -- 1031 - 0x407  :   10 - 0xa
    "10010000", -- 1032 - 0x408  :  144 - 0x90 -- Background 0x81
    "00010000", -- 1033 - 0x409  :   16 - 0x10
    "00011111", -- 1034 - 0x40a  :   31 - 0x1f
    "00010000", -- 1035 - 0x40b  :   16 - 0x10
    "00011111", -- 1036 - 0x40c  :   31 - 0x1f
    "00010000", -- 1037 - 0x40d  :   16 - 0x10
    "00010000", -- 1038 - 0x40e  :   16 - 0x10
    "10010000", -- 1039 - 0x40f  :  144 - 0x90
    "00111111", -- 1040 - 0x410  :   63 - 0x3f -- Background 0x82
    "01111000", -- 1041 - 0x411  :  120 - 0x78
    "11100111", -- 1042 - 0x412  :  231 - 0xe7
    "11001111", -- 1043 - 0x413  :  207 - 0xcf
    "01011000", -- 1044 - 0x414  :   88 - 0x58
    "01011000", -- 1045 - 0x415  :   88 - 0x58
    "01010000", -- 1046 - 0x416  :   80 - 0x50
    "10010000", -- 1047 - 0x417  :  144 - 0x90
    "10110000", -- 1048 - 0x418  :  176 - 0xb0 -- Background 0x83
    "11111100", -- 1049 - 0x419  :  252 - 0xfc
    "11100010", -- 1050 - 0x41a  :  226 - 0xe2
    "11000001", -- 1051 - 0x41b  :  193 - 0xc1
    "11000001", -- 1052 - 0x41c  :  193 - 0xc1
    "10000011", -- 1053 - 0x41d  :  131 - 0x83
    "10001111", -- 1054 - 0x41e  :  143 - 0x8f
    "01111110", -- 1055 - 0x41f  :  126 - 0x7e
    "11111110", -- 1056 - 0x420  :  254 - 0xfe -- Background 0x84
    "00000011", -- 1057 - 0x421  :    3 - 0x3
    "00001111", -- 1058 - 0x422  :   15 - 0xf
    "10010001", -- 1059 - 0x423  :  145 - 0x91
    "01110000", -- 1060 - 0x424  :  112 - 0x70
    "01100000", -- 1061 - 0x425  :   96 - 0x60
    "00100000", -- 1062 - 0x426  :   32 - 0x20
    "00110001", -- 1063 - 0x427  :   49 - 0x31
    "00111111", -- 1064 - 0x428  :   63 - 0x3f -- Background 0x85
    "00111111", -- 1065 - 0x429  :   63 - 0x3f
    "00011101", -- 1066 - 0x42a  :   29 - 0x1d
    "00111001", -- 1067 - 0x42b  :   57 - 0x39
    "01111011", -- 1068 - 0x42c  :  123 - 0x7b
    "11110011", -- 1069 - 0x42d  :  243 - 0xf3
    "10000110", -- 1070 - 0x42e  :  134 - 0x86
    "11111110", -- 1071 - 0x42f  :  254 - 0xfe
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Background 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "10000000", -- 1077 - 0x435  :  128 - 0x80
    "10000000", -- 1078 - 0x436  :  128 - 0x80
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "11111110", -- 1080 - 0x438  :  254 - 0xfe -- Background 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "00000011", -- 1085 - 0x43d  :    3 - 0x3
    "00000011", -- 1086 - 0x43e  :    3 - 0x3
    "11111111", -- 1087 - 0x43f  :  255 - 0xff
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "11111111", -- 1090 - 0x442  :  255 - 0xff
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00111100", -- 1096 - 0x448  :   60 - 0x3c -- Background 0x89
    "11111100", -- 1097 - 0x449  :  252 - 0xfc
    "11111100", -- 1098 - 0x44a  :  252 - 0xfc
    "11111100", -- 1099 - 0x44b  :  252 - 0xfc
    "11111100", -- 1100 - 0x44c  :  252 - 0xfc
    "11111100", -- 1101 - 0x44d  :  252 - 0xfc
    "00000100", -- 1102 - 0x44e  :    4 - 0x4
    "00000100", -- 1103 - 0x44f  :    4 - 0x4
    "11111111", -- 1104 - 0x450  :  255 - 0xff -- Background 0x8a
    "11111111", -- 1105 - 0x451  :  255 - 0xff
    "11111111", -- 1106 - 0x452  :  255 - 0xff
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "10000000", -- 1108 - 0x454  :  128 - 0x80
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- Background 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "00000011", -- 1116 - 0x45c  :    3 - 0x3
    "11111111", -- 1117 - 0x45d  :  255 - 0xff
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11111111", -- 1119 - 0x45f  :  255 - 0xff
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Background 0x8c
    "11111111", -- 1121 - 0x461  :  255 - 0xff
    "11111111", -- 1122 - 0x462  :  255 - 0xff
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "11111111", -- 1126 - 0x466  :  255 - 0xff
    "11111111", -- 1127 - 0x467  :  255 - 0xff
    "11111100", -- 1128 - 0x468  :  252 - 0xfc -- Background 0x8d
    "11111100", -- 1129 - 0x469  :  252 - 0xfc
    "11111110", -- 1130 - 0x46a  :  254 - 0xfe
    "11111110", -- 1131 - 0x46b  :  254 - 0xfe
    "11111110", -- 1132 - 0x46c  :  254 - 0xfe
    "00000010", -- 1133 - 0x46d  :    2 - 0x2
    "11111110", -- 1134 - 0x46e  :  254 - 0xfe
    "11111110", -- 1135 - 0x46f  :  254 - 0xfe
    "11111111", -- 1136 - 0x470  :  255 - 0xff -- Background 0x8e
    "10000000", -- 1137 - 0x471  :  128 - 0x80
    "10000000", -- 1138 - 0x472  :  128 - 0x80
    "10000000", -- 1139 - 0x473  :  128 - 0x80
    "10000000", -- 1140 - 0x474  :  128 - 0x80
    "10000000", -- 1141 - 0x475  :  128 - 0x80
    "10000000", -- 1142 - 0x476  :  128 - 0x80
    "10000000", -- 1143 - 0x477  :  128 - 0x80
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- Background 0x8f
    "00000011", -- 1145 - 0x479  :    3 - 0x3
    "00000011", -- 1146 - 0x47a  :    3 - 0x3
    "00000011", -- 1147 - 0x47b  :    3 - 0x3
    "00000011", -- 1148 - 0x47c  :    3 - 0x3
    "00000011", -- 1149 - 0x47d  :    3 - 0x3
    "00000011", -- 1150 - 0x47e  :    3 - 0x3
    "00000011", -- 1151 - 0x47f  :    3 - 0x3
    "00000010", -- 1152 - 0x480  :    2 - 0x2 -- Background 0x90
    "00000010", -- 1153 - 0x481  :    2 - 0x2
    "00000010", -- 1154 - 0x482  :    2 - 0x2
    "00000010", -- 1155 - 0x483  :    2 - 0x2
    "00000010", -- 1156 - 0x484  :    2 - 0x2
    "00000010", -- 1157 - 0x485  :    2 - 0x2
    "00000100", -- 1158 - 0x486  :    4 - 0x4
    "00000100", -- 1159 - 0x487  :    4 - 0x4
    "10000000", -- 1160 - 0x488  :  128 - 0x80 -- Background 0x91
    "10000000", -- 1161 - 0x489  :  128 - 0x80
    "10101010", -- 1162 - 0x48a  :  170 - 0xaa
    "11010101", -- 1163 - 0x48b  :  213 - 0xd5
    "10101010", -- 1164 - 0x48c  :  170 - 0xaa
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "00000011", -- 1168 - 0x490  :    3 - 0x3 -- Background 0x92
    "00000011", -- 1169 - 0x491  :    3 - 0x3
    "10101011", -- 1170 - 0x492  :  171 - 0xab
    "01010111", -- 1171 - 0x493  :   87 - 0x57
    "10101011", -- 1172 - 0x494  :  171 - 0xab
    "11111111", -- 1173 - 0x495  :  255 - 0xff
    "11111111", -- 1174 - 0x496  :  255 - 0xff
    "11111110", -- 1175 - 0x497  :  254 - 0xfe
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- Background 0x93
    "01010101", -- 1177 - 0x499  :   85 - 0x55
    "10101010", -- 1178 - 0x49a  :  170 - 0xaa
    "01010101", -- 1179 - 0x49b  :   85 - 0x55
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000100", -- 1184 - 0x4a0  :    4 - 0x4 -- Background 0x94
    "01010100", -- 1185 - 0x4a1  :   84 - 0x54
    "10101100", -- 1186 - 0x4a2  :  172 - 0xac
    "01011100", -- 1187 - 0x4a3  :   92 - 0x5c
    "11111100", -- 1188 - 0x4a4  :  252 - 0xfc
    "11111100", -- 1189 - 0x4a5  :  252 - 0xfc
    "11111100", -- 1190 - 0x4a6  :  252 - 0xfc
    "00111100", -- 1191 - 0x4a7  :   60 - 0x3c
    "00111111", -- 1192 - 0x4a8  :   63 - 0x3f -- Background 0x95
    "00111111", -- 1193 - 0x4a9  :   63 - 0x3f
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00111111", -- 1195 - 0x4ab  :   63 - 0x3f
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "11111111", -- 1199 - 0x4af  :  255 - 0xff
    "01111110", -- 1200 - 0x4b0  :  126 - 0x7e -- Background 0x96
    "01111100", -- 1201 - 0x4b1  :  124 - 0x7c
    "01111100", -- 1202 - 0x4b2  :  124 - 0x7c
    "01111000", -- 1203 - 0x4b3  :  120 - 0x78
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "00011111", -- 1208 - 0x4b8  :   31 - 0x1f -- Background 0x97
    "00001111", -- 1209 - 0x4b9  :   15 - 0xf
    "00001111", -- 1210 - 0x4ba  :   15 - 0xf
    "00000111", -- 1211 - 0x4bb  :    7 - 0x7
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "11111111", -- 1215 - 0x4bf  :  255 - 0xff
    "11111110", -- 1216 - 0x4c0  :  254 - 0xfe -- Background 0x98
    "11111100", -- 1217 - 0x4c1  :  252 - 0xfc
    "11111100", -- 1218 - 0x4c2  :  252 - 0xfc
    "11111000", -- 1219 - 0x4c3  :  248 - 0xf8
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "11111111", -- 1228 - 0x4cc  :  255 - 0xff
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00011000", -- 1232 - 0x4d0  :   24 - 0x18 -- Background 0x9a
    "00011000", -- 1233 - 0x4d1  :   24 - 0x18
    "00011000", -- 1234 - 0x4d2  :   24 - 0x18
    "00011000", -- 1235 - 0x4d3  :   24 - 0x18
    "00011000", -- 1236 - 0x4d4  :   24 - 0x18
    "00011000", -- 1237 - 0x4d5  :   24 - 0x18
    "00011000", -- 1238 - 0x4d6  :   24 - 0x18
    "00011000", -- 1239 - 0x4d7  :   24 - 0x18
    "00000111", -- 1240 - 0x4d8  :    7 - 0x7 -- Background 0x9b
    "00011111", -- 1241 - 0x4d9  :   31 - 0x1f
    "00111111", -- 1242 - 0x4da  :   63 - 0x3f
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "01111111", -- 1244 - 0x4dc  :  127 - 0x7f
    "01111111", -- 1245 - 0x4dd  :  127 - 0x7f
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11100001", -- 1248 - 0x4e0  :  225 - 0xe1 -- Background 0x9c
    "11111001", -- 1249 - 0x4e1  :  249 - 0xf9
    "11111101", -- 1250 - 0x4e2  :  253 - 0xfd
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111110", -- 1252 - 0x4e4  :  254 - 0xfe
    "11111110", -- 1253 - 0x4e5  :  254 - 0xfe
    "11111111", -- 1254 - 0x4e6  :  255 - 0xff
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "11110000", -- 1256 - 0x4e8  :  240 - 0xf0 -- Background 0x9d
    "00010000", -- 1257 - 0x4e9  :   16 - 0x10
    "00010000", -- 1258 - 0x4ea  :   16 - 0x10
    "00010000", -- 1259 - 0x4eb  :   16 - 0x10
    "00010000", -- 1260 - 0x4ec  :   16 - 0x10
    "00010000", -- 1261 - 0x4ed  :   16 - 0x10
    "00010000", -- 1262 - 0x4ee  :   16 - 0x10
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "00011111", -- 1264 - 0x4f0  :   31 - 0x1f -- Background 0x9e
    "00010000", -- 1265 - 0x4f1  :   16 - 0x10
    "00010000", -- 1266 - 0x4f2  :   16 - 0x10
    "00010000", -- 1267 - 0x4f3  :   16 - 0x10
    "00010000", -- 1268 - 0x4f4  :   16 - 0x10
    "00010000", -- 1269 - 0x4f5  :   16 - 0x10
    "00010000", -- 1270 - 0x4f6  :   16 - 0x10
    "11111111", -- 1271 - 0x4f7  :  255 - 0xff
    "10010010", -- 1272 - 0x4f8  :  146 - 0x92 -- Background 0x9f
    "10010010", -- 1273 - 0x4f9  :  146 - 0x92
    "10010010", -- 1274 - 0x4fa  :  146 - 0x92
    "11111110", -- 1275 - 0x4fb  :  254 - 0xfe
    "11111110", -- 1276 - 0x4fc  :  254 - 0xfe
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00001010", -- 1280 - 0x500  :   10 - 0xa -- Background 0xa0
    "00001010", -- 1281 - 0x501  :   10 - 0xa
    "00111010", -- 1282 - 0x502  :   58 - 0x3a
    "00001010", -- 1283 - 0x503  :   10 - 0xa
    "11111011", -- 1284 - 0x504  :  251 - 0xfb
    "00001011", -- 1285 - 0x505  :   11 - 0xb
    "00001011", -- 1286 - 0x506  :   11 - 0xb
    "00001011", -- 1287 - 0x507  :   11 - 0xb
    "10010000", -- 1288 - 0x508  :  144 - 0x90 -- Background 0xa1
    "10010000", -- 1289 - 0x509  :  144 - 0x90
    "10011111", -- 1290 - 0x50a  :  159 - 0x9f
    "10010000", -- 1291 - 0x50b  :  144 - 0x90
    "10011111", -- 1292 - 0x50c  :  159 - 0x9f
    "10010000", -- 1293 - 0x50d  :  144 - 0x90
    "10010000", -- 1294 - 0x50e  :  144 - 0x90
    "10010000", -- 1295 - 0x50f  :  144 - 0x90
    "00000001", -- 1296 - 0x510  :    1 - 0x1 -- Background 0xa2
    "00000001", -- 1297 - 0x511  :    1 - 0x1
    "00000001", -- 1298 - 0x512  :    1 - 0x1
    "00000001", -- 1299 - 0x513  :    1 - 0x1
    "00000001", -- 1300 - 0x514  :    1 - 0x1
    "00000001", -- 1301 - 0x515  :    1 - 0x1
    "00000001", -- 1302 - 0x516  :    1 - 0x1
    "00000001", -- 1303 - 0x517  :    1 - 0x1
    "10000000", -- 1304 - 0x518  :  128 - 0x80 -- Background 0xa3
    "10000000", -- 1305 - 0x519  :  128 - 0x80
    "10000000", -- 1306 - 0x51a  :  128 - 0x80
    "10000000", -- 1307 - 0x51b  :  128 - 0x80
    "10000000", -- 1308 - 0x51c  :  128 - 0x80
    "10000000", -- 1309 - 0x51d  :  128 - 0x80
    "10000000", -- 1310 - 0x51e  :  128 - 0x80
    "10000000", -- 1311 - 0x51f  :  128 - 0x80
    "00001000", -- 1312 - 0x520  :    8 - 0x8 -- Background 0xa4
    "10001000", -- 1313 - 0x521  :  136 - 0x88
    "10010001", -- 1314 - 0x522  :  145 - 0x91
    "11010001", -- 1315 - 0x523  :  209 - 0xd1
    "01010011", -- 1316 - 0x524  :   83 - 0x53
    "01010011", -- 1317 - 0x525  :   83 - 0x53
    "01110011", -- 1318 - 0x526  :  115 - 0x73
    "00111111", -- 1319 - 0x527  :   63 - 0x3f
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000111", -- 1322 - 0x52a  :    7 - 0x7
    "00001111", -- 1323 - 0x52b  :   15 - 0xf
    "00001100", -- 1324 - 0x52c  :   12 - 0xc
    "00011011", -- 1325 - 0x52d  :   27 - 0x1b
    "00011011", -- 1326 - 0x52e  :   27 - 0x1b
    "00011011", -- 1327 - 0x52f  :   27 - 0x1b
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "11100000", -- 1330 - 0x532  :  224 - 0xe0
    "11110000", -- 1331 - 0x533  :  240 - 0xf0
    "11110000", -- 1332 - 0x534  :  240 - 0xf0
    "11111000", -- 1333 - 0x535  :  248 - 0xf8
    "11111000", -- 1334 - 0x536  :  248 - 0xf8
    "11111000", -- 1335 - 0x537  :  248 - 0xf8
    "00011011", -- 1336 - 0x538  :   27 - 0x1b -- Background 0xa7
    "00011011", -- 1337 - 0x539  :   27 - 0x1b
    "00011011", -- 1338 - 0x53a  :   27 - 0x1b
    "00011011", -- 1339 - 0x53b  :   27 - 0x1b
    "00011011", -- 1340 - 0x53c  :   27 - 0x1b
    "00001111", -- 1341 - 0x53d  :   15 - 0xf
    "00001111", -- 1342 - 0x53e  :   15 - 0xf
    "00000111", -- 1343 - 0x53f  :    7 - 0x7
    "11111000", -- 1344 - 0x540  :  248 - 0xf8 -- Background 0xa8
    "11111000", -- 1345 - 0x541  :  248 - 0xf8
    "11111000", -- 1346 - 0x542  :  248 - 0xf8
    "11111000", -- 1347 - 0x543  :  248 - 0xf8
    "11111000", -- 1348 - 0x544  :  248 - 0xf8
    "11110000", -- 1349 - 0x545  :  240 - 0xf0
    "11110000", -- 1350 - 0x546  :  240 - 0xf0
    "11100000", -- 1351 - 0x547  :  224 - 0xe0
    "11110001", -- 1352 - 0x548  :  241 - 0xf1 -- Background 0xa9
    "00010001", -- 1353 - 0x549  :   17 - 0x11
    "00010001", -- 1354 - 0x54a  :   17 - 0x11
    "00011111", -- 1355 - 0x54b  :   31 - 0x1f
    "00010000", -- 1356 - 0x54c  :   16 - 0x10
    "00010000", -- 1357 - 0x54d  :   16 - 0x10
    "00010000", -- 1358 - 0x54e  :   16 - 0x10
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "00011111", -- 1360 - 0x550  :   31 - 0x1f -- Background 0xaa
    "00010000", -- 1361 - 0x551  :   16 - 0x10
    "00010000", -- 1362 - 0x552  :   16 - 0x10
    "11110000", -- 1363 - 0x553  :  240 - 0xf0
    "00010000", -- 1364 - 0x554  :   16 - 0x10
    "00010000", -- 1365 - 0x555  :   16 - 0x10
    "00010000", -- 1366 - 0x556  :   16 - 0x10
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "01111111", -- 1368 - 0x558  :  127 - 0x7f -- Background 0xab
    "10111111", -- 1369 - 0x559  :  191 - 0xbf
    "11011111", -- 1370 - 0x55a  :  223 - 0xdf
    "11101111", -- 1371 - 0x55b  :  239 - 0xef
    "11110000", -- 1372 - 0x55c  :  240 - 0xf0
    "11110000", -- 1373 - 0x55d  :  240 - 0xf0
    "11110000", -- 1374 - 0x55e  :  240 - 0xf0
    "11110000", -- 1375 - 0x55f  :  240 - 0xf0
    "11110000", -- 1376 - 0x560  :  240 - 0xf0 -- Background 0xac
    "11110000", -- 1377 - 0x561  :  240 - 0xf0
    "11110000", -- 1378 - 0x562  :  240 - 0xf0
    "11110000", -- 1379 - 0x563  :  240 - 0xf0
    "11111111", -- 1380 - 0x564  :  255 - 0xff
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "11111111", -- 1382 - 0x566  :  255 - 0xff
    "11111111", -- 1383 - 0x567  :  255 - 0xff
    "11111111", -- 1384 - 0x568  :  255 - 0xff -- Background 0xad
    "11111111", -- 1385 - 0x569  :  255 - 0xff
    "11111111", -- 1386 - 0x56a  :  255 - 0xff
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "00001111", -- 1388 - 0x56c  :   15 - 0xf
    "00001111", -- 1389 - 0x56d  :   15 - 0xf
    "00001111", -- 1390 - 0x56e  :   15 - 0xf
    "00001111", -- 1391 - 0x56f  :   15 - 0xf
    "00001111", -- 1392 - 0x570  :   15 - 0xf -- Background 0xae
    "00001111", -- 1393 - 0x571  :   15 - 0xf
    "00001111", -- 1394 - 0x572  :   15 - 0xf
    "00001111", -- 1395 - 0x573  :   15 - 0xf
    "11110111", -- 1396 - 0x574  :  247 - 0xf7
    "11111011", -- 1397 - 0x575  :  251 - 0xfb
    "11111101", -- 1398 - 0x576  :  253 - 0xfd
    "11111110", -- 1399 - 0x577  :  254 - 0xfe
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00011000", -- 1406 - 0x57e  :   24 - 0x18
    "00011000", -- 1407 - 0x57f  :   24 - 0x18
    "00011111", -- 1408 - 0x580  :   31 - 0x1f -- Background 0xb0
    "00111111", -- 1409 - 0x581  :   63 - 0x3f
    "01111111", -- 1410 - 0x582  :  127 - 0x7f
    "01111111", -- 1411 - 0x583  :  127 - 0x7f
    "01111111", -- 1412 - 0x584  :  127 - 0x7f
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "11111111", -- 1416 - 0x588  :  255 - 0xff -- Background 0xb1
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11111111", -- 1418 - 0x58a  :  255 - 0xff
    "01111111", -- 1419 - 0x58b  :  127 - 0x7f
    "01111111", -- 1420 - 0x58c  :  127 - 0x7f
    "01111111", -- 1421 - 0x58d  :  127 - 0x7f
    "00111111", -- 1422 - 0x58e  :   63 - 0x3f
    "00011110", -- 1423 - 0x58f  :   30 - 0x1e
    "11111000", -- 1424 - 0x590  :  248 - 0xf8 -- Background 0xb2
    "11111100", -- 1425 - 0x591  :  252 - 0xfc
    "11111110", -- 1426 - 0x592  :  254 - 0xfe
    "11111110", -- 1427 - 0x593  :  254 - 0xfe
    "11111110", -- 1428 - 0x594  :  254 - 0xfe
    "11111111", -- 1429 - 0x595  :  255 - 0xff
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff -- Background 0xb3
    "11111111", -- 1433 - 0x599  :  255 - 0xff
    "11111111", -- 1434 - 0x59a  :  255 - 0xff
    "11111110", -- 1435 - 0x59b  :  254 - 0xfe
    "11111110", -- 1436 - 0x59c  :  254 - 0xfe
    "11111110", -- 1437 - 0x59d  :  254 - 0xfe
    "11111100", -- 1438 - 0x59e  :  252 - 0xfc
    "01111000", -- 1439 - 0x59f  :  120 - 0x78
    "01111111", -- 1440 - 0x5a0  :  127 - 0x7f -- Background 0xb4
    "10000000", -- 1441 - 0x5a1  :  128 - 0x80
    "10000000", -- 1442 - 0x5a2  :  128 - 0x80
    "10000000", -- 1443 - 0x5a3  :  128 - 0x80
    "10000000", -- 1444 - 0x5a4  :  128 - 0x80
    "10000000", -- 1445 - 0x5a5  :  128 - 0x80
    "10000000", -- 1446 - 0x5a6  :  128 - 0x80
    "10000000", -- 1447 - 0x5a7  :  128 - 0x80
    "11011110", -- 1448 - 0x5a8  :  222 - 0xde -- Background 0xb5
    "01100001", -- 1449 - 0x5a9  :   97 - 0x61
    "01100001", -- 1450 - 0x5aa  :   97 - 0x61
    "01100001", -- 1451 - 0x5ab  :   97 - 0x61
    "01110001", -- 1452 - 0x5ac  :  113 - 0x71
    "01011110", -- 1453 - 0x5ad  :   94 - 0x5e
    "01111111", -- 1454 - 0x5ae  :  127 - 0x7f
    "01100001", -- 1455 - 0x5af  :   97 - 0x61
    "10000000", -- 1456 - 0x5b0  :  128 - 0x80 -- Background 0xb6
    "10000000", -- 1457 - 0x5b1  :  128 - 0x80
    "11000000", -- 1458 - 0x5b2  :  192 - 0xc0
    "11110000", -- 1459 - 0x5b3  :  240 - 0xf0
    "10111111", -- 1460 - 0x5b4  :  191 - 0xbf
    "10001111", -- 1461 - 0x5b5  :  143 - 0x8f
    "10000001", -- 1462 - 0x5b6  :  129 - 0x81
    "01111110", -- 1463 - 0x5b7  :  126 - 0x7e
    "01100001", -- 1464 - 0x5b8  :   97 - 0x61 -- Background 0xb7
    "01100001", -- 1465 - 0x5b9  :   97 - 0x61
    "11000001", -- 1466 - 0x5ba  :  193 - 0xc1
    "11000001", -- 1467 - 0x5bb  :  193 - 0xc1
    "10000001", -- 1468 - 0x5bc  :  129 - 0x81
    "10000001", -- 1469 - 0x5bd  :  129 - 0x81
    "10000011", -- 1470 - 0x5be  :  131 - 0x83
    "11111110", -- 1471 - 0x5bf  :  254 - 0xfe
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000011", -- 1474 - 0x5c2  :    3 - 0x3
    "00001111", -- 1475 - 0x5c3  :   15 - 0xf
    "00011111", -- 1476 - 0x5c4  :   31 - 0x1f
    "00111111", -- 1477 - 0x5c5  :   63 - 0x3f
    "01111111", -- 1478 - 0x5c6  :  127 - 0x7f
    "01111111", -- 1479 - 0x5c7  :  127 - 0x7f
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- Background 0xb9
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "11000000", -- 1482 - 0x5ca  :  192 - 0xc0
    "11110000", -- 1483 - 0x5cb  :  240 - 0xf0
    "11111000", -- 1484 - 0x5cc  :  248 - 0xf8
    "11111100", -- 1485 - 0x5cd  :  252 - 0xfc
    "11111110", -- 1486 - 0x5ce  :  254 - 0xfe
    "11111110", -- 1487 - 0x5cf  :  254 - 0xfe
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Background 0xba
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "11111111", -- 1490 - 0x5d2  :  255 - 0xff
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "11111111", -- 1492 - 0x5d4  :  255 - 0xff
    "11111111", -- 1493 - 0x5d5  :  255 - 0xff
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "11111111", -- 1496 - 0x5d8  :  255 - 0xff -- Background 0xbb
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111111", -- 1499 - 0x5db  :  255 - 0xff
    "11111111", -- 1500 - 0x5dc  :  255 - 0xff
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "01111111", -- 1504 - 0x5e0  :  127 - 0x7f -- Background 0xbc
    "01111111", -- 1505 - 0x5e1  :  127 - 0x7f
    "01111111", -- 1506 - 0x5e2  :  127 - 0x7f
    "00111111", -- 1507 - 0x5e3  :   63 - 0x3f
    "00111111", -- 1508 - 0x5e4  :   63 - 0x3f
    "00011111", -- 1509 - 0x5e5  :   31 - 0x1f
    "00001111", -- 1510 - 0x5e6  :   15 - 0xf
    "00000111", -- 1511 - 0x5e7  :    7 - 0x7
    "11111110", -- 1512 - 0x5e8  :  254 - 0xfe -- Background 0xbd
    "11111110", -- 1513 - 0x5e9  :  254 - 0xfe
    "11111110", -- 1514 - 0x5ea  :  254 - 0xfe
    "11111100", -- 1515 - 0x5eb  :  252 - 0xfc
    "11111100", -- 1516 - 0x5ec  :  252 - 0xfc
    "11111000", -- 1517 - 0x5ed  :  248 - 0xf8
    "11110000", -- 1518 - 0x5ee  :  240 - 0xf0
    "11110000", -- 1519 - 0x5ef  :  240 - 0xf0
    "00001111", -- 1520 - 0x5f0  :   15 - 0xf -- Background 0xbe
    "00001111", -- 1521 - 0x5f1  :   15 - 0xf
    "00001111", -- 1522 - 0x5f2  :   15 - 0xf
    "00001111", -- 1523 - 0x5f3  :   15 - 0xf
    "00001111", -- 1524 - 0x5f4  :   15 - 0xf
    "00001111", -- 1525 - 0x5f5  :   15 - 0xf
    "00000111", -- 1526 - 0x5f6  :    7 - 0x7
    "00001111", -- 1527 - 0x5f7  :   15 - 0xf
    "11110000", -- 1528 - 0x5f8  :  240 - 0xf0 -- Background 0xbf
    "11110000", -- 1529 - 0x5f9  :  240 - 0xf0
    "11110000", -- 1530 - 0x5fa  :  240 - 0xf0
    "11110000", -- 1531 - 0x5fb  :  240 - 0xf0
    "11110000", -- 1532 - 0x5fc  :  240 - 0xf0
    "11110000", -- 1533 - 0x5fd  :  240 - 0xf0
    "11100000", -- 1534 - 0x5fe  :  224 - 0xe0
    "11110000", -- 1535 - 0x5ff  :  240 - 0xf0
    "10000001", -- 1536 - 0x600  :  129 - 0x81 -- Background 0xc0
    "11000001", -- 1537 - 0x601  :  193 - 0xc1
    "10100011", -- 1538 - 0x602  :  163 - 0xa3
    "10100011", -- 1539 - 0x603  :  163 - 0xa3
    "10011101", -- 1540 - 0x604  :  157 - 0x9d
    "10000001", -- 1541 - 0x605  :  129 - 0x81
    "10000001", -- 1542 - 0x606  :  129 - 0x81
    "10000001", -- 1543 - 0x607  :  129 - 0x81
    "11100011", -- 1544 - 0x608  :  227 - 0xe3 -- Background 0xc1
    "11110111", -- 1545 - 0x609  :  247 - 0xf7
    "11000001", -- 1546 - 0x60a  :  193 - 0xc1
    "11000001", -- 1547 - 0x60b  :  193 - 0xc1
    "11000001", -- 1548 - 0x60c  :  193 - 0xc1
    "11000001", -- 1549 - 0x60d  :  193 - 0xc1
    "11110111", -- 1550 - 0x60e  :  247 - 0xf7
    "11100011", -- 1551 - 0x60f  :  227 - 0xe3
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000111", -- 1554 - 0x612  :    7 - 0x7
    "00001111", -- 1555 - 0x613  :   15 - 0xf
    "00001100", -- 1556 - 0x614  :   12 - 0xc
    "00011011", -- 1557 - 0x615  :   27 - 0x1b
    "00011011", -- 1558 - 0x616  :   27 - 0x1b
    "00011011", -- 1559 - 0x617  :   27 - 0x1b
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "11100000", -- 1562 - 0x61a  :  224 - 0xe0
    "11110000", -- 1563 - 0x61b  :  240 - 0xf0
    "11110000", -- 1564 - 0x61c  :  240 - 0xf0
    "11111000", -- 1565 - 0x61d  :  248 - 0xf8
    "11111000", -- 1566 - 0x61e  :  248 - 0xf8
    "11111000", -- 1567 - 0x61f  :  248 - 0xf8
    "00011011", -- 1568 - 0x620  :   27 - 0x1b -- Background 0xc4
    "00011011", -- 1569 - 0x621  :   27 - 0x1b
    "00011011", -- 1570 - 0x622  :   27 - 0x1b
    "00011011", -- 1571 - 0x623  :   27 - 0x1b
    "00011011", -- 1572 - 0x624  :   27 - 0x1b
    "00001111", -- 1573 - 0x625  :   15 - 0xf
    "00001111", -- 1574 - 0x626  :   15 - 0xf
    "00000111", -- 1575 - 0x627  :    7 - 0x7
    "11111000", -- 1576 - 0x628  :  248 - 0xf8 -- Background 0xc5
    "11111000", -- 1577 - 0x629  :  248 - 0xf8
    "11111000", -- 1578 - 0x62a  :  248 - 0xf8
    "11111000", -- 1579 - 0x62b  :  248 - 0xf8
    "11111000", -- 1580 - 0x62c  :  248 - 0xf8
    "11110000", -- 1581 - 0x62d  :  240 - 0xf0
    "11110000", -- 1582 - 0x62e  :  240 - 0xf0
    "11100000", -- 1583 - 0x62f  :  224 - 0xe0
    "11100000", -- 1584 - 0x630  :  224 - 0xe0 -- Background 0xc6
    "11111111", -- 1585 - 0x631  :  255 - 0xff
    "11111111", -- 1586 - 0x632  :  255 - 0xff
    "11111111", -- 1587 - 0x633  :  255 - 0xff
    "11111111", -- 1588 - 0x634  :  255 - 0xff
    "11111111", -- 1589 - 0x635  :  255 - 0xff
    "11111111", -- 1590 - 0x636  :  255 - 0xff
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "00000111", -- 1592 - 0x638  :    7 - 0x7 -- Background 0xc7
    "11111111", -- 1593 - 0x639  :  255 - 0xff
    "11111111", -- 1594 - 0x63a  :  255 - 0xff
    "11111111", -- 1595 - 0x63b  :  255 - 0xff
    "11111111", -- 1596 - 0x63c  :  255 - 0xff
    "11111111", -- 1597 - 0x63d  :  255 - 0xff
    "11111111", -- 1598 - 0x63e  :  255 - 0xff
    "11111111", -- 1599 - 0x63f  :  255 - 0xff
    "11111111", -- 1600 - 0x640  :  255 - 0xff -- Background 0xc8
    "11111111", -- 1601 - 0x641  :  255 - 0xff
    "11111111", -- 1602 - 0x642  :  255 - 0xff
    "11111111", -- 1603 - 0x643  :  255 - 0xff
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "11111110", -- 1605 - 0x645  :  254 - 0xfe
    "11111111", -- 1606 - 0x646  :  255 - 0xff
    "11101111", -- 1607 - 0x647  :  239 - 0xef
    "11111111", -- 1608 - 0x648  :  255 - 0xff -- Background 0xc9
    "11011111", -- 1609 - 0x649  :  223 - 0xdf
    "11101111", -- 1610 - 0x64a  :  239 - 0xef
    "10101111", -- 1611 - 0x64b  :  175 - 0xaf
    "10101111", -- 1612 - 0x64c  :  175 - 0xaf
    "01101111", -- 1613 - 0x64d  :  111 - 0x6f
    "11101111", -- 1614 - 0x64e  :  239 - 0xef
    "11100111", -- 1615 - 0x64f  :  231 - 0xe7
    "00011111", -- 1616 - 0x650  :   31 - 0x1f -- Background 0xca
    "00011111", -- 1617 - 0x651  :   31 - 0x1f
    "00111111", -- 1618 - 0x652  :   63 - 0x3f
    "00111111", -- 1619 - 0x653  :   63 - 0x3f
    "01110000", -- 1620 - 0x654  :  112 - 0x70
    "01100011", -- 1621 - 0x655  :   99 - 0x63
    "11100111", -- 1622 - 0x656  :  231 - 0xe7
    "11100101", -- 1623 - 0x657  :  229 - 0xe5
    "11110000", -- 1624 - 0x658  :  240 - 0xf0 -- Background 0xcb
    "11110000", -- 1625 - 0x659  :  240 - 0xf0
    "11111000", -- 1626 - 0x65a  :  248 - 0xf8
    "11111000", -- 1627 - 0x65b  :  248 - 0xf8
    "00001100", -- 1628 - 0x65c  :   12 - 0xc
    "11000100", -- 1629 - 0x65d  :  196 - 0xc4
    "11100100", -- 1630 - 0x65e  :  228 - 0xe4
    "10100110", -- 1631 - 0x65f  :  166 - 0xa6
    "11101001", -- 1632 - 0x660  :  233 - 0xe9 -- Background 0xcc
    "11101001", -- 1633 - 0x661  :  233 - 0xe9
    "11101001", -- 1634 - 0x662  :  233 - 0xe9
    "11101111", -- 1635 - 0x663  :  239 - 0xef
    "11100010", -- 1636 - 0x664  :  226 - 0xe2
    "11100011", -- 1637 - 0x665  :  227 - 0xe3
    "11110000", -- 1638 - 0x666  :  240 - 0xf0
    "11111111", -- 1639 - 0x667  :  255 - 0xff
    "10010110", -- 1640 - 0x668  :  150 - 0x96 -- Background 0xcd
    "10010110", -- 1641 - 0x669  :  150 - 0x96
    "10010110", -- 1642 - 0x66a  :  150 - 0x96
    "11110110", -- 1643 - 0x66b  :  246 - 0xf6
    "01000110", -- 1644 - 0x66c  :   70 - 0x46
    "11000110", -- 1645 - 0x66d  :  198 - 0xc6
    "00001110", -- 1646 - 0x66e  :   14 - 0xe
    "11111110", -- 1647 - 0x66f  :  254 - 0xfe
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Background 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "01111110", -- 1654 - 0x676  :  126 - 0x7e
    "00111100", -- 1655 - 0x677  :   60 - 0x3c
    "00111100", -- 1656 - 0x678  :   60 - 0x3c -- Background 0xcf
    "01000010", -- 1657 - 0x679  :   66 - 0x42
    "10011001", -- 1658 - 0x67a  :  153 - 0x99
    "10100001", -- 1659 - 0x67b  :  161 - 0xa1
    "10100001", -- 1660 - 0x67c  :  161 - 0xa1
    "10011001", -- 1661 - 0x67d  :  153 - 0x99
    "01000010", -- 1662 - 0x67e  :   66 - 0x42
    "00111100", -- 1663 - 0x67f  :   60 - 0x3c
    "00001111", -- 1664 - 0x680  :   15 - 0xf -- Background 0xd0
    "00011111", -- 1665 - 0x681  :   31 - 0x1f
    "00011111", -- 1666 - 0x682  :   31 - 0x1f
    "00111111", -- 1667 - 0x683  :   63 - 0x3f
    "00111111", -- 1668 - 0x684  :   63 - 0x3f
    "01111111", -- 1669 - 0x685  :  127 - 0x7f
    "01111111", -- 1670 - 0x686  :  127 - 0x7f
    "01111111", -- 1671 - 0x687  :  127 - 0x7f
    "11110000", -- 1672 - 0x688  :  240 - 0xf0 -- Background 0xd1
    "11111000", -- 1673 - 0x689  :  248 - 0xf8
    "11111000", -- 1674 - 0x68a  :  248 - 0xf8
    "11111100", -- 1675 - 0x68b  :  252 - 0xfc
    "11111100", -- 1676 - 0x68c  :  252 - 0xfc
    "11111110", -- 1677 - 0x68d  :  254 - 0xfe
    "11111110", -- 1678 - 0x68e  :  254 - 0xfe
    "11111110", -- 1679 - 0x68f  :  254 - 0xfe
    "01111111", -- 1680 - 0x690  :  127 - 0x7f -- Background 0xd2
    "01111111", -- 1681 - 0x691  :  127 - 0x7f
    "00111111", -- 1682 - 0x692  :   63 - 0x3f
    "00111111", -- 1683 - 0x693  :   63 - 0x3f
    "00111111", -- 1684 - 0x694  :   63 - 0x3f
    "00111111", -- 1685 - 0x695  :   63 - 0x3f
    "00011111", -- 1686 - 0x696  :   31 - 0x1f
    "00011111", -- 1687 - 0x697  :   31 - 0x1f
    "11111110", -- 1688 - 0x698  :  254 - 0xfe -- Background 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111100", -- 1692 - 0x69c  :  252 - 0xfc
    "11111100", -- 1693 - 0x69d  :  252 - 0xfc
    "11111110", -- 1694 - 0x69e  :  254 - 0xfe
    "11111110", -- 1695 - 0x69f  :  254 - 0xfe
    "01111111", -- 1696 - 0x6a0  :  127 - 0x7f -- Background 0xd4
    "01111111", -- 1697 - 0x6a1  :  127 - 0x7f
    "01111111", -- 1698 - 0x6a2  :  127 - 0x7f
    "00111111", -- 1699 - 0x6a3  :   63 - 0x3f
    "00111111", -- 1700 - 0x6a4  :   63 - 0x3f
    "00111111", -- 1701 - 0x6a5  :   63 - 0x3f
    "00111111", -- 1702 - 0x6a6  :   63 - 0x3f
    "00011111", -- 1703 - 0x6a7  :   31 - 0x1f
    "11111110", -- 1704 - 0x6a8  :  254 - 0xfe -- Background 0xd5
    "11111110", -- 1705 - 0x6a9  :  254 - 0xfe
    "11111111", -- 1706 - 0x6aa  :  255 - 0xff
    "11111111", -- 1707 - 0x6ab  :  255 - 0xff
    "11111111", -- 1708 - 0x6ac  :  255 - 0xff
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111110", -- 1711 - 0x6af  :  254 - 0xfe
    "00011111", -- 1712 - 0x6b0  :   31 - 0x1f -- Background 0xd6
    "00001111", -- 1713 - 0x6b1  :   15 - 0xf
    "00001111", -- 1714 - 0x6b2  :   15 - 0xf
    "00000111", -- 1715 - 0x6b3  :    7 - 0x7
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "11111110", -- 1720 - 0x6b8  :  254 - 0xfe -- Background 0xd7
    "11111100", -- 1721 - 0x6b9  :  252 - 0xfc
    "11111100", -- 1722 - 0x6ba  :  252 - 0xfc
    "11111000", -- 1723 - 0x6bb  :  248 - 0xf8
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "01111110", -- 1728 - 0x6c0  :  126 - 0x7e -- Background 0xd8
    "01111110", -- 1729 - 0x6c1  :  126 - 0x7e
    "01111110", -- 1730 - 0x6c2  :  126 - 0x7e
    "01111110", -- 1731 - 0x6c3  :  126 - 0x7e
    "01111111", -- 1732 - 0x6c4  :  127 - 0x7f
    "01111111", -- 1733 - 0x6c5  :  127 - 0x7f
    "01111111", -- 1734 - 0x6c6  :  127 - 0x7f
    "01111111", -- 1735 - 0x6c7  :  127 - 0x7f
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- Background 0xd9
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11111111", -- 1740 - 0x6cc  :  255 - 0xff
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111111", -- 1742 - 0x6ce  :  255 - 0xff
    "11111110", -- 1743 - 0x6cf  :  254 - 0xfe
    "11111110", -- 1744 - 0x6d0  :  254 - 0xfe -- Background 0xda
    "11111110", -- 1745 - 0x6d1  :  254 - 0xfe
    "11111110", -- 1746 - 0x6d2  :  254 - 0xfe
    "11111110", -- 1747 - 0x6d3  :  254 - 0xfe
    "11111111", -- 1748 - 0x6d4  :  255 - 0xff
    "11111111", -- 1749 - 0x6d5  :  255 - 0xff
    "11111111", -- 1750 - 0x6d6  :  255 - 0xff
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "01111111", -- 1752 - 0x6d8  :  127 - 0x7f -- Background 0xdb
    "01111111", -- 1753 - 0x6d9  :  127 - 0x7f
    "01111111", -- 1754 - 0x6da  :  127 - 0x7f
    "01111111", -- 1755 - 0x6db  :  127 - 0x7f
    "01111111", -- 1756 - 0x6dc  :  127 - 0x7f
    "01111111", -- 1757 - 0x6dd  :  127 - 0x7f
    "01111111", -- 1758 - 0x6de  :  127 - 0x7f
    "01111111", -- 1759 - 0x6df  :  127 - 0x7f
    "11111111", -- 1760 - 0x6e0  :  255 - 0xff -- Background 0xdc
    "11111111", -- 1761 - 0x6e1  :  255 - 0xff
    "11111111", -- 1762 - 0x6e2  :  255 - 0xff
    "11111111", -- 1763 - 0x6e3  :  255 - 0xff
    "11111100", -- 1764 - 0x6e4  :  252 - 0xfc
    "11111110", -- 1765 - 0x6e5  :  254 - 0xfe
    "11111110", -- 1766 - 0x6e6  :  254 - 0xfe
    "01111110", -- 1767 - 0x6e7  :  126 - 0x7e
    "11111111", -- 1768 - 0x6e8  :  255 - 0xff -- Background 0xdd
    "11111111", -- 1769 - 0x6e9  :  255 - 0xff
    "11111111", -- 1770 - 0x6ea  :  255 - 0xff
    "11111111", -- 1771 - 0x6eb  :  255 - 0xff
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "01111111", -- 1776 - 0x6f0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "01111111", -- 1778 - 0x6f2  :  127 - 0x7f
    "01111111", -- 1779 - 0x6f3  :  127 - 0x7f
    "01111111", -- 1780 - 0x6f4  :  127 - 0x7f
    "01111111", -- 1781 - 0x6f5  :  127 - 0x7f
    "01111111", -- 1782 - 0x6f6  :  127 - 0x7f
    "01111111", -- 1783 - 0x6f7  :  127 - 0x7f
    "11111111", -- 1784 - 0x6f8  :  255 - 0xff -- Background 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11111111", -- 1788 - 0x6fc  :  255 - 0xff
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111110", -- 1791 - 0x6ff  :  254 - 0xfe
    "01111110", -- 1792 - 0x700  :  126 - 0x7e -- Background 0xe0
    "01111110", -- 1793 - 0x701  :  126 - 0x7e
    "01111111", -- 1794 - 0x702  :  127 - 0x7f
    "01111111", -- 1795 - 0x703  :  127 - 0x7f
    "01111111", -- 1796 - 0x704  :  127 - 0x7f
    "01111111", -- 1797 - 0x705  :  127 - 0x7f
    "01111111", -- 1798 - 0x706  :  127 - 0x7f
    "01111111", -- 1799 - 0x707  :  127 - 0x7f
    "00111111", -- 1800 - 0x708  :   63 - 0x3f -- Background 0xe1
    "00111111", -- 1801 - 0x709  :   63 - 0x3f
    "00111111", -- 1802 - 0x70a  :   63 - 0x3f
    "00111111", -- 1803 - 0x70b  :   63 - 0x3f
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "01111110", -- 1808 - 0x710  :  126 - 0x7e -- Background 0xe2
    "01111100", -- 1809 - 0x711  :  124 - 0x7c
    "01111100", -- 1810 - 0x712  :  124 - 0x7c
    "01111000", -- 1811 - 0x713  :  120 - 0x78
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "11111110", -- 1816 - 0x718  :  254 - 0xfe -- Background 0xe3
    "11111110", -- 1817 - 0x719  :  254 - 0xfe
    "11111111", -- 1818 - 0x71a  :  255 - 0xff
    "11111111", -- 1819 - 0x71b  :  255 - 0xff
    "01111111", -- 1820 - 0x71c  :  127 - 0x7f
    "01111111", -- 1821 - 0x71d  :  127 - 0x7f
    "01111111", -- 1822 - 0x71e  :  127 - 0x7f
    "01111111", -- 1823 - 0x71f  :  127 - 0x7f
    "01111111", -- 1824 - 0x720  :  127 - 0x7f -- Background 0xe4
    "01111111", -- 1825 - 0x721  :  127 - 0x7f
    "00111111", -- 1826 - 0x722  :   63 - 0x3f
    "00111111", -- 1827 - 0x723  :   63 - 0x3f
    "00111111", -- 1828 - 0x724  :   63 - 0x3f
    "00111111", -- 1829 - 0x725  :   63 - 0x3f
    "00011111", -- 1830 - 0x726  :   31 - 0x1f
    "00011111", -- 1831 - 0x727  :   31 - 0x1f
    "00111111", -- 1832 - 0x728  :   63 - 0x3f -- Background 0xe5
    "10111111", -- 1833 - 0x729  :  191 - 0xbf
    "11111111", -- 1834 - 0x72a  :  255 - 0xff
    "11111111", -- 1835 - 0x72b  :  255 - 0xff
    "11111100", -- 1836 - 0x72c  :  252 - 0xfc
    "11111100", -- 1837 - 0x72d  :  252 - 0xfc
    "11111110", -- 1838 - 0x72e  :  254 - 0xfe
    "11111110", -- 1839 - 0x72f  :  254 - 0xfe
    "01111111", -- 1840 - 0x730  :  127 - 0x7f -- Background 0xe6
    "01111111", -- 1841 - 0x731  :  127 - 0x7f
    "01111110", -- 1842 - 0x732  :  126 - 0x7e
    "01111110", -- 1843 - 0x733  :  126 - 0x7e
    "01111111", -- 1844 - 0x734  :  127 - 0x7f
    "01111111", -- 1845 - 0x735  :  127 - 0x7f
    "01111111", -- 1846 - 0x736  :  127 - 0x7f
    "01111111", -- 1847 - 0x737  :  127 - 0x7f
    "01111110", -- 1848 - 0x738  :  126 - 0x7e -- Background 0xe7
    "01111110", -- 1849 - 0x739  :  126 - 0x7e
    "01111110", -- 1850 - 0x73a  :  126 - 0x7e
    "01111110", -- 1851 - 0x73b  :  126 - 0x7e
    "01111111", -- 1852 - 0x73c  :  127 - 0x7f
    "01111111", -- 1853 - 0x73d  :  127 - 0x7f
    "01111111", -- 1854 - 0x73e  :  127 - 0x7f
    "01111111", -- 1855 - 0x73f  :  127 - 0x7f
    "10000001", -- 1856 - 0x740  :  129 - 0x81 -- Background 0xe8
    "11000011", -- 1857 - 0x741  :  195 - 0xc3
    "11000011", -- 1858 - 0x742  :  195 - 0xc3
    "11100111", -- 1859 - 0x743  :  231 - 0xe7
    "11100111", -- 1860 - 0x744  :  231 - 0xe7
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "00001111", -- 1864 - 0x748  :   15 - 0xf -- Background 0xe9
    "01000011", -- 1865 - 0x749  :   67 - 0x43
    "01011011", -- 1866 - 0x74a  :   91 - 0x5b
    "01010011", -- 1867 - 0x74b  :   83 - 0x53
    "00110001", -- 1868 - 0x74c  :   49 - 0x31
    "00011001", -- 1869 - 0x74d  :   25 - 0x19
    "00001111", -- 1870 - 0x74e  :   15 - 0xf
    "00000111", -- 1871 - 0x74f  :    7 - 0x7
    "11000001", -- 1872 - 0x750  :  193 - 0xc1 -- Background 0xea
    "11000011", -- 1873 - 0x751  :  195 - 0xc3
    "11000110", -- 1874 - 0x752  :  198 - 0xc6
    "10000100", -- 1875 - 0x753  :  132 - 0x84
    "11111100", -- 1876 - 0x754  :  252 - 0xfc
    "11111100", -- 1877 - 0x755  :  252 - 0xfc
    "00001110", -- 1878 - 0x756  :   14 - 0xe
    "00000010", -- 1879 - 0x757  :    2 - 0x2
    "00010000", -- 1880 - 0x758  :   16 - 0x10 -- Background 0xeb
    "00100000", -- 1881 - 0x759  :   32 - 0x20
    "00100010", -- 1882 - 0x75a  :   34 - 0x22
    "10111010", -- 1883 - 0x75b  :  186 - 0xba
    "11100110", -- 1884 - 0x75c  :  230 - 0xe6
    "11100001", -- 1885 - 0x75d  :  225 - 0xe1
    "11000000", -- 1886 - 0x75e  :  192 - 0xc0
    "11000000", -- 1887 - 0x75f  :  192 - 0xc0
    "00100000", -- 1888 - 0x760  :   32 - 0x20 -- Background 0xec
    "10100110", -- 1889 - 0x761  :  166 - 0xa6
    "01010100", -- 1890 - 0x762  :   84 - 0x54
    "00100110", -- 1891 - 0x763  :   38 - 0x26
    "00100000", -- 1892 - 0x764  :   32 - 0x20
    "11000110", -- 1893 - 0x765  :  198 - 0xc6
    "01010100", -- 1894 - 0x766  :   84 - 0x54
    "00100110", -- 1895 - 0x767  :   38 - 0x26
    "00100000", -- 1896 - 0x768  :   32 - 0x20 -- Background 0xed
    "10000101", -- 1897 - 0x769  :  133 - 0x85
    "00000001", -- 1898 - 0x76a  :    1 - 0x1
    "01000100", -- 1899 - 0x76b  :   68 - 0x44
    "00100000", -- 1900 - 0x76c  :   32 - 0x20
    "10000110", -- 1901 - 0x76d  :  134 - 0x86
    "01010100", -- 1902 - 0x76e  :   84 - 0x54
    "01001000", -- 1903 - 0x76f  :   72 - 0x48
    "00100000", -- 1904 - 0x770  :   32 - 0x20 -- Background 0xee
    "10111010", -- 1905 - 0x771  :  186 - 0xba
    "11001001", -- 1906 - 0x772  :  201 - 0xc9
    "01001010", -- 1907 - 0x773  :   74 - 0x4a
    "00100000", -- 1908 - 0x774  :   32 - 0x20
    "10100110", -- 1909 - 0x775  :  166 - 0xa6
    "00001010", -- 1910 - 0x776  :   10 - 0xa
    "11010000", -- 1911 - 0x777  :  208 - 0xd0
    "11010001", -- 1912 - 0x778  :  209 - 0xd1 -- Background 0xef
    "00100000", -- 1913 - 0x779  :   32 - 0x20
    "11000110", -- 1914 - 0x77a  :  198 - 0xc6
    "00001010", -- 1915 - 0x77b  :   10 - 0xa
    "11010010", -- 1916 - 0x77c  :  210 - 0xd2
    "11010011", -- 1917 - 0x77d  :  211 - 0xd3
    "11011011", -- 1918 - 0x77e  :  219 - 0xdb
    "11011011", -- 1919 - 0x77f  :  219 - 0xdb
    "00001010", -- 1920 - 0x780  :   10 - 0xa -- Background 0xf0
    "11010100", -- 1921 - 0x781  :  212 - 0xd4
    "11010101", -- 1922 - 0x782  :  213 - 0xd5
    "11010100", -- 1923 - 0x783  :  212 - 0xd4
    "11011001", -- 1924 - 0x784  :  217 - 0xd9
    "11011011", -- 1925 - 0x785  :  219 - 0xdb
    "11100010", -- 1926 - 0x786  :  226 - 0xe2
    "11010100", -- 1927 - 0x787  :  212 - 0xd4
    "11010110", -- 1928 - 0x788  :  214 - 0xd6 -- Background 0xf1
    "11010111", -- 1929 - 0x789  :  215 - 0xd7
    "11100001", -- 1930 - 0x78a  :  225 - 0xe1
    "00100110", -- 1931 - 0x78b  :   38 - 0x26
    "11010110", -- 1932 - 0x78c  :  214 - 0xd6
    "11011101", -- 1933 - 0x78d  :  221 - 0xdd
    "11100001", -- 1934 - 0x78e  :  225 - 0xe1
    "11100001", -- 1935 - 0x78f  :  225 - 0xe1
    "11011110", -- 1936 - 0x790  :  222 - 0xde -- Background 0xf2
    "11010001", -- 1937 - 0x791  :  209 - 0xd1
    "11011000", -- 1938 - 0x792  :  216 - 0xd8
    "11010000", -- 1939 - 0x793  :  208 - 0xd0
    "11010001", -- 1940 - 0x794  :  209 - 0xd1
    "00100110", -- 1941 - 0x795  :   38 - 0x26
    "11011110", -- 1942 - 0x796  :  222 - 0xde
    "11010001", -- 1943 - 0x797  :  209 - 0xd1
    "01000110", -- 1944 - 0x798  :   70 - 0x46 -- Background 0xf3
    "00010100", -- 1945 - 0x799  :   20 - 0x14
    "11011011", -- 1946 - 0x79a  :  219 - 0xdb
    "01000010", -- 1947 - 0x79b  :   66 - 0x42
    "01000010", -- 1948 - 0x79c  :   66 - 0x42
    "11011011", -- 1949 - 0x79d  :  219 - 0xdb
    "01000010", -- 1950 - 0x79e  :   66 - 0x42
    "11011011", -- 1951 - 0x79f  :  219 - 0xdb
    "01000010", -- 1952 - 0x7a0  :   66 - 0x42 -- Background 0xf4
    "11011011", -- 1953 - 0x7a1  :  219 - 0xdb
    "01000010", -- 1954 - 0x7a2  :   66 - 0x42
    "11011011", -- 1955 - 0x7a3  :  219 - 0xdb
    "01000010", -- 1956 - 0x7a4  :   66 - 0x42
    "00100110", -- 1957 - 0x7a5  :   38 - 0x26
    "00100001", -- 1958 - 0x7a6  :   33 - 0x21
    "01100110", -- 1959 - 0x7a7  :  102 - 0x66
    "11011011", -- 1960 - 0x7a8  :  219 - 0xdb -- Background 0xf5
    "00100110", -- 1961 - 0x7a9  :   38 - 0x26
    "11011011", -- 1962 - 0x7aa  :  219 - 0xdb
    "11011111", -- 1963 - 0x7ab  :  223 - 0xdf
    "11011011", -- 1964 - 0x7ac  :  219 - 0xdb
    "11011111", -- 1965 - 0x7ad  :  223 - 0xdf
    "11011011", -- 1966 - 0x7ae  :  219 - 0xdb
    "11011011", -- 1967 - 0x7af  :  219 - 0xdb
    "11011011", -- 1968 - 0x7b0  :  219 - 0xdb -- Background 0xf6
    "11011110", -- 1969 - 0x7b1  :  222 - 0xde
    "01000011", -- 1970 - 0x7b2  :   67 - 0x43
    "11011011", -- 1971 - 0x7b3  :  219 - 0xdb
    "11100000", -- 1972 - 0x7b4  :  224 - 0xe0
    "11011011", -- 1973 - 0x7b5  :  219 - 0xdb
    "11011011", -- 1974 - 0x7b6  :  219 - 0xdb
    "11011011", -- 1975 - 0x7b7  :  219 - 0xdb
    "11100011", -- 1976 - 0x7b8  :  227 - 0xe3 -- Background 0xf7
    "00100110", -- 1977 - 0x7b9  :   38 - 0x26
    "00100001", -- 1978 - 0x7ba  :   33 - 0x21
    "10100110", -- 1979 - 0x7bb  :  166 - 0xa6
    "00010100", -- 1980 - 0x7bc  :   20 - 0x14
    "11011011", -- 1981 - 0x7bd  :  219 - 0xdb
    "11011011", -- 1982 - 0x7be  :  219 - 0xdb
    "11011011", -- 1983 - 0x7bf  :  219 - 0xdb
    "11011011", -- 1984 - 0x7c0  :  219 - 0xdb -- Background 0xf8
    "11011001", -- 1985 - 0x7c1  :  217 - 0xd9
    "11011011", -- 1986 - 0x7c2  :  219 - 0xdb
    "11011011", -- 1987 - 0x7c3  :  219 - 0xdb
    "11010100", -- 1988 - 0x7c4  :  212 - 0xd4
    "11011001", -- 1989 - 0x7c5  :  217 - 0xd9
    "11010100", -- 1990 - 0x7c6  :  212 - 0xd4
    "11011001", -- 1991 - 0x7c7  :  217 - 0xd9
    "10010101", -- 1992 - 0x7c8  :  149 - 0x95 -- Background 0xf9
    "10010101", -- 1993 - 0x7c9  :  149 - 0x95
    "10010101", -- 1994 - 0x7ca  :  149 - 0x95
    "10010101", -- 1995 - 0x7cb  :  149 - 0x95
    "10010101", -- 1996 - 0x7cc  :  149 - 0x95
    "10010111", -- 1997 - 0x7cd  :  151 - 0x97
    "10011000", -- 1998 - 0x7ce  :  152 - 0x98
    "01111000", -- 1999 - 0x7cf  :  120 - 0x78
    "10010101", -- 2000 - 0x7d0  :  149 - 0x95 -- Background 0xfa
    "01111010", -- 2001 - 0x7d1  :  122 - 0x7a
    "00100001", -- 2002 - 0x7d2  :   33 - 0x21
    "11101101", -- 2003 - 0x7d3  :  237 - 0xed
    "00001110", -- 2004 - 0x7d4  :   14 - 0xe
    "11001111", -- 2005 - 0x7d5  :  207 - 0xcf
    "00000001", -- 2006 - 0x7d6  :    1 - 0x1
    "00001001", -- 2007 - 0x7d7  :    9 - 0x9
    "00010111", -- 2008 - 0x7d8  :   23 - 0x17 -- Background 0xfb
    "00001101", -- 2009 - 0x7d9  :   13 - 0xd
    "00011000", -- 2010 - 0x7da  :   24 - 0x18
    "00100010", -- 2011 - 0x7db  :   34 - 0x22
    "01001011", -- 2012 - 0x7dc  :   75 - 0x4b
    "00001101", -- 2013 - 0x7dd  :   13 - 0xd
    "00000001", -- 2014 - 0x7de  :    1 - 0x1
    "00100100", -- 2015 - 0x7df  :   36 - 0x24
    "00001010", -- 2016 - 0x7e0  :   10 - 0xa -- Background 0xfc
    "00010110", -- 2017 - 0x7e1  :   22 - 0x16
    "00001110", -- 2018 - 0x7e2  :   14 - 0xe
    "00100010", -- 2019 - 0x7e3  :   34 - 0x22
    "10001011", -- 2020 - 0x7e4  :  139 - 0x8b
    "00001101", -- 2021 - 0x7e5  :   13 - 0xd
    "00000010", -- 2022 - 0x7e6  :    2 - 0x2
    "00100100", -- 2023 - 0x7e7  :   36 - 0x24
    "00001010", -- 2024 - 0x7e8  :   10 - 0xa -- Background 0xfd
    "00010110", -- 2025 - 0x7e9  :   22 - 0x16
    "00001110", -- 2026 - 0x7ea  :   14 - 0xe
    "00100010", -- 2027 - 0x7eb  :   34 - 0x22
    "11101100", -- 2028 - 0x7ec  :  236 - 0xec
    "00000100", -- 2029 - 0x7ed  :    4 - 0x4
    "00011101", -- 2030 - 0x7ee  :   29 - 0x1d
    "00011000", -- 2031 - 0x7ef  :   24 - 0x18
    "01010110", -- 2032 - 0x7f0  :   86 - 0x56 -- Background 0xfe
    "01010101", -- 2033 - 0x7f1  :   85 - 0x55
    "00100011", -- 2034 - 0x7f2  :   35 - 0x23
    "11100010", -- 2035 - 0x7f3  :  226 - 0xe2
    "00000100", -- 2036 - 0x7f4  :    4 - 0x4
    "10011001", -- 2037 - 0x7f5  :  153 - 0x99
    "10101010", -- 2038 - 0x7f6  :  170 - 0xaa
    "10101010", -- 2039 - 0x7f7  :  170 - 0xaa
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Background 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
