---   Sprites Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN_SPR is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN_SPR;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN_SPR is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table both color planes
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x1
    "00111000", --   17 - 0x11  :   56 - 0x38
    "01111100", --   18 - 0x12  :  124 - 0x7c
    "11111110", --   19 - 0x13  :  254 - 0xfe
    "11111110", --   20 - 0x14  :  254 - 0xfe
    "11111110", --   21 - 0x15  :  254 - 0xfe
    "01111100", --   22 - 0x16  :  124 - 0x7c
    "00111000", --   23 - 0x17  :   56 - 0x38
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00111000", --   25 - 0x19  :   56 - 0x38
    "01111100", --   26 - 0x1a  :  124 - 0x7c
    "11111110", --   27 - 0x1b  :  254 - 0xfe
    "11111110", --   28 - 0x1c  :  254 - 0xfe
    "11111110", --   29 - 0x1d  :  254 - 0xfe
    "01111100", --   30 - 0x1e  :  124 - 0x7c
    "00111000", --   31 - 0x1f  :   56 - 0x38
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00011000", --   51 - 0x33  :   24 - 0x18
    "00011000", --   52 - 0x34  :   24 - 0x18
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- plane 1
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00011000", --   59 - 0x3b  :   24 - 0x18
    "00011000", --   60 - 0x3c  :   24 - 0x18
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "11111111", --   72 - 0x48  :  255 - 0xff -- plane 1
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00001111", --   88 - 0x58  :   15 - 0xf -- plane 1
    "00001111", --   89 - 0x59  :   15 - 0xf
    "00001111", --   90 - 0x5a  :   15 - 0xf
    "00001111", --   91 - 0x5b  :   15 - 0xf
    "00001111", --   92 - 0x5c  :   15 - 0xf
    "00001111", --   93 - 0x5d  :   15 - 0xf
    "00001111", --   94 - 0x5e  :   15 - 0xf
    "00001111", --   95 - 0x5f  :   15 - 0xf
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11110000", --  104 - 0x68  :  240 - 0xf0 -- plane 1
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11110000", --  106 - 0x6a  :  240 - 0xf0
    "11110000", --  107 - 0x6b  :  240 - 0xf0
    "11110000", --  108 - 0x6c  :  240 - 0xf0
    "11110000", --  109 - 0x6d  :  240 - 0xf0
    "11110000", --  110 - 0x6e  :  240 - 0xf0
    "11110000", --  111 - 0x6f  :  240 - 0xf0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0x7
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- plane 1
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x8
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- plane 1
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x9
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00011000", --  148 - 0x94  :   24 - 0x18
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- plane 1
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00011000", --  155 - 0x9b  :   24 - 0x18
    "00011000", --  156 - 0x9c  :   24 - 0x18
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0xa
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- plane 1
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0xb
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- plane 1
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- plane 1
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0xd
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- plane 1
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- plane 1
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- plane 1
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  257 - 0x101  :    0 - 0x0
    "11111111", --  258 - 0x102  :  255 - 0xff
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "11111111", --  261 - 0x105  :  255 - 0xff
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- plane 1
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00100100", --  272 - 0x110  :   36 - 0x24 -- Sprite 0x11
    "00100100", --  273 - 0x111  :   36 - 0x24
    "00100100", --  274 - 0x112  :   36 - 0x24
    "00100100", --  275 - 0x113  :   36 - 0x24
    "00100100", --  276 - 0x114  :   36 - 0x24
    "00100100", --  277 - 0x115  :   36 - 0x24
    "00100100", --  278 - 0x116  :   36 - 0x24
    "00100100", --  279 - 0x117  :   36 - 0x24
    "00000000", --  280 - 0x118  :    0 - 0x0 -- plane 1
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00100100", --  288 - 0x120  :   36 - 0x24 -- Sprite 0x12
    "00100100", --  289 - 0x121  :   36 - 0x24
    "11000011", --  290 - 0x122  :  195 - 0xc3
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "11111111", --  293 - 0x125  :  255 - 0xff
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- plane 1
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  305 - 0x131  :    0 - 0x0
    "11111111", --  306 - 0x132  :  255 - 0xff
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "11000011", --  309 - 0x135  :  195 - 0xc3
    "00100100", --  310 - 0x136  :   36 - 0x24
    "00100100", --  311 - 0x137  :   36 - 0x24
    "00000000", --  312 - 0x138  :    0 - 0x0 -- plane 1
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00100100", --  320 - 0x140  :   36 - 0x24 -- Sprite 0x14
    "00100100", --  321 - 0x141  :   36 - 0x24
    "11000100", --  322 - 0x142  :  196 - 0xc4
    "00000100", --  323 - 0x143  :    4 - 0x4
    "00000100", --  324 - 0x144  :    4 - 0x4
    "11000100", --  325 - 0x145  :  196 - 0xc4
    "00100100", --  326 - 0x146  :   36 - 0x24
    "00100100", --  327 - 0x147  :   36 - 0x24
    "00000000", --  328 - 0x148  :    0 - 0x0 -- plane 1
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00100100", --  336 - 0x150  :   36 - 0x24 -- Sprite 0x15
    "00100100", --  337 - 0x151  :   36 - 0x24
    "00100011", --  338 - 0x152  :   35 - 0x23
    "00100000", --  339 - 0x153  :   32 - 0x20
    "00100000", --  340 - 0x154  :   32 - 0x20
    "00100011", --  341 - 0x155  :   35 - 0x23
    "00100100", --  342 - 0x156  :   36 - 0x24
    "00100100", --  343 - 0x157  :   36 - 0x24
    "00000000", --  344 - 0x158  :    0 - 0x0 -- plane 1
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00001111", --  354 - 0x162  :   15 - 0xf
    "00010000", --  355 - 0x163  :   16 - 0x10
    "11110000", --  356 - 0x164  :  240 - 0xf0
    "00001111", --  357 - 0x165  :   15 - 0xf
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- plane 1
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x17
    "00000000", --  369 - 0x171  :    0 - 0x0
    "11110000", --  370 - 0x172  :  240 - 0xf0
    "00001000", --  371 - 0x173  :    8 - 0x8
    "00001111", --  372 - 0x174  :   15 - 0xf
    "11110000", --  373 - 0x175  :  240 - 0xf0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- plane 1
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  385 - 0x181  :    0 - 0x0
    "11110000", --  386 - 0x182  :  240 - 0xf0
    "00001000", --  387 - 0x183  :    8 - 0x8
    "00001000", --  388 - 0x184  :    8 - 0x8
    "11110000", --  389 - 0x185  :  240 - 0xf0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- plane 1
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x19
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00001111", --  402 - 0x192  :   15 - 0xf
    "00010000", --  403 - 0x193  :   16 - 0x10
    "00010000", --  404 - 0x194  :   16 - 0x10
    "00001111", --  405 - 0x195  :   15 - 0xf
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- plane 1
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00100100", --  416 - 0x1a0  :   36 - 0x24 -- Sprite 0x1a
    "00100100", --  417 - 0x1a1  :   36 - 0x24
    "00100100", --  418 - 0x1a2  :   36 - 0x24
    "00100100", --  419 - 0x1a3  :   36 - 0x24
    "00011000", --  420 - 0x1a4  :   24 - 0x18
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- plane 1
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00011000", --  435 - 0x1b3  :   24 - 0x18
    "00100100", --  436 - 0x1b4  :   36 - 0x24
    "00100100", --  437 - 0x1b5  :   36 - 0x24
    "00100100", --  438 - 0x1b6  :   36 - 0x24
    "00100100", --  439 - 0x1b7  :   36 - 0x24
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- plane 1
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00100100", --  448 - 0x1c0  :   36 - 0x24 -- Sprite 0x1c
    "00100100", --  449 - 0x1c1  :   36 - 0x24
    "11000100", --  450 - 0x1c2  :  196 - 0xc4
    "00000100", --  451 - 0x1c3  :    4 - 0x4
    "00001000", --  452 - 0x1c4  :    8 - 0x8
    "11110000", --  453 - 0x1c5  :  240 - 0xf0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- plane 1
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x1d
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "11110000", --  466 - 0x1d2  :  240 - 0xf0
    "00001000", --  467 - 0x1d3  :    8 - 0x8
    "00000100", --  468 - 0x1d4  :    4 - 0x4
    "11000100", --  469 - 0x1d5  :  196 - 0xc4
    "00100100", --  470 - 0x1d6  :   36 - 0x24
    "00100100", --  471 - 0x1d7  :   36 - 0x24
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- plane 1
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00100100", --  480 - 0x1e0  :   36 - 0x24 -- Sprite 0x1e
    "00100100", --  481 - 0x1e1  :   36 - 0x24
    "00100011", --  482 - 0x1e2  :   35 - 0x23
    "00100000", --  483 - 0x1e3  :   32 - 0x20
    "00010000", --  484 - 0x1e4  :   16 - 0x10
    "00001111", --  485 - 0x1e5  :   15 - 0xf
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- plane 1
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00001111", --  498 - 0x1f2  :   15 - 0xf
    "00010000", --  499 - 0x1f3  :   16 - 0x10
    "00100000", --  500 - 0x1f4  :   32 - 0x20
    "00100011", --  501 - 0x1f5  :   35 - 0x23
    "00100100", --  502 - 0x1f6  :   36 - 0x24
    "00100100", --  503 - 0x1f7  :   36 - 0x24
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- plane 1
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  529 - 0x211  :    0 - 0x0
    "11110000", --  530 - 0x212  :  240 - 0xf0
    "00001000", --  531 - 0x213  :    8 - 0x8
    "00001000", --  532 - 0x214  :    8 - 0x8
    "11110000", --  533 - 0x215  :  240 - 0xf0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00001111", --  536 - 0x218  :   15 - 0xf -- plane 1
    "00001111", --  537 - 0x219  :   15 - 0xf
    "00001111", --  538 - 0x21a  :   15 - 0xf
    "00000111", --  539 - 0x21b  :    7 - 0x7
    "00000111", --  540 - 0x21c  :    7 - 0x7
    "00001111", --  541 - 0x21d  :   15 - 0xf
    "00001111", --  542 - 0x21e  :   15 - 0xf
    "00001111", --  543 - 0x21f  :   15 - 0xf
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00001111", --  546 - 0x222  :   15 - 0xf
    "00010000", --  547 - 0x223  :   16 - 0x10
    "00010000", --  548 - 0x224  :   16 - 0x10
    "00001111", --  549 - 0x225  :   15 - 0xf
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "11110000", --  552 - 0x228  :  240 - 0xf0 -- plane 1
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11110000", --  554 - 0x22a  :  240 - 0xf0
    "11100000", --  555 - 0x22b  :  224 - 0xe0
    "11100000", --  556 - 0x22c  :  224 - 0xe0
    "11110000", --  557 - 0x22d  :  240 - 0xf0
    "11110000", --  558 - 0x22e  :  240 - 0xf0
    "11110000", --  559 - 0x22f  :  240 - 0xf0
    "11111111", --  560 - 0x230  :  255 - 0xff -- Sprite 0x23
    "11111111", --  561 - 0x231  :  255 - 0xff
    "11100001", --  562 - 0x232  :  225 - 0xe1
    "11100001", --  563 - 0x233  :  225 - 0xe1
    "11100001", --  564 - 0x234  :  225 - 0xe1
    "11100001", --  565 - 0x235  :  225 - 0xe1
    "11100001", --  566 - 0x236  :  225 - 0xe1
    "11100001", --  567 - 0x237  :  225 - 0xe1
    "11111111", --  568 - 0x238  :  255 - 0xff -- plane 1
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11100001", --  570 - 0x23a  :  225 - 0xe1
    "11100001", --  571 - 0x23b  :  225 - 0xe1
    "11100001", --  572 - 0x23c  :  225 - 0xe1
    "11100001", --  573 - 0x23d  :  225 - 0xe1
    "11100001", --  574 - 0x23e  :  225 - 0xe1
    "11100001", --  575 - 0x23f  :  225 - 0xe1
    "10000111", --  576 - 0x240  :  135 - 0x87 -- Sprite 0x24
    "11000111", --  577 - 0x241  :  199 - 0xc7
    "11000000", --  578 - 0x242  :  192 - 0xc0
    "11000111", --  579 - 0x243  :  199 - 0xc7
    "11001111", --  580 - 0x244  :  207 - 0xcf
    "11001110", --  581 - 0x245  :  206 - 0xce
    "11001111", --  582 - 0x246  :  207 - 0xcf
    "11000111", --  583 - 0x247  :  199 - 0xc7
    "10000111", --  584 - 0x248  :  135 - 0x87 -- plane 1
    "11000111", --  585 - 0x249  :  199 - 0xc7
    "11000000", --  586 - 0x24a  :  192 - 0xc0
    "11000111", --  587 - 0x24b  :  199 - 0xc7
    "11001111", --  588 - 0x24c  :  207 - 0xcf
    "11001110", --  589 - 0x24d  :  206 - 0xce
    "11001111", --  590 - 0x24e  :  207 - 0xcf
    "11000111", --  591 - 0x24f  :  199 - 0xc7
    "11111000", --  592 - 0x250  :  248 - 0xf8 -- Sprite 0x25
    "11111100", --  593 - 0x251  :  252 - 0xfc
    "00011100", --  594 - 0x252  :   28 - 0x1c
    "11111100", --  595 - 0x253  :  252 - 0xfc
    "11111100", --  596 - 0x254  :  252 - 0xfc
    "00011100", --  597 - 0x255  :   28 - 0x1c
    "11111100", --  598 - 0x256  :  252 - 0xfc
    "11111100", --  599 - 0x257  :  252 - 0xfc
    "11111000", --  600 - 0x258  :  248 - 0xf8 -- plane 1
    "11111100", --  601 - 0x259  :  252 - 0xfc
    "00011100", --  602 - 0x25a  :   28 - 0x1c
    "11111100", --  603 - 0x25b  :  252 - 0xfc
    "11111100", --  604 - 0x25c  :  252 - 0xfc
    "00011100", --  605 - 0x25d  :   28 - 0x1c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x26
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11100111", --  610 - 0x262  :  231 - 0xe7
    "11100111", --  611 - 0x263  :  231 - 0xe7
    "11100111", --  612 - 0x264  :  231 - 0xe7
    "11100111", --  613 - 0x265  :  231 - 0xe7
    "11100111", --  614 - 0x266  :  231 - 0xe7
    "11100111", --  615 - 0x267  :  231 - 0xe7
    "11111111", --  616 - 0x268  :  255 - 0xff -- plane 1
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11100111", --  618 - 0x26a  :  231 - 0xe7
    "11100111", --  619 - 0x26b  :  231 - 0xe7
    "11100111", --  620 - 0x26c  :  231 - 0xe7
    "11100111", --  621 - 0x26d  :  231 - 0xe7
    "11100111", --  622 - 0x26e  :  231 - 0xe7
    "11100111", --  623 - 0x26f  :  231 - 0xe7
    "11110000", --  624 - 0x270  :  240 - 0xf0 -- Sprite 0x27
    "11111001", --  625 - 0x271  :  249 - 0xf9
    "00111001", --  626 - 0x272  :   57 - 0x39
    "00111001", --  627 - 0x273  :   57 - 0x39
    "00111001", --  628 - 0x274  :   57 - 0x39
    "00111001", --  629 - 0x275  :   57 - 0x39
    "00111001", --  630 - 0x276  :   57 - 0x39
    "00111000", --  631 - 0x277  :   56 - 0x38
    "11110000", --  632 - 0x278  :  240 - 0xf0 -- plane 1
    "11111001", --  633 - 0x279  :  249 - 0xf9
    "00111001", --  634 - 0x27a  :   57 - 0x39
    "00111001", --  635 - 0x27b  :   57 - 0x39
    "00111001", --  636 - 0x27c  :   57 - 0x39
    "00111001", --  637 - 0x27d  :   57 - 0x39
    "00111001", --  638 - 0x27e  :   57 - 0x39
    "00111000", --  639 - 0x27f  :   56 - 0x38
    "11111111", --  640 - 0x280  :  255 - 0xff -- Sprite 0x28
    "11111111", --  641 - 0x281  :  255 - 0xff
    "11000000", --  642 - 0x282  :  192 - 0xc0
    "11000000", --  643 - 0x283  :  192 - 0xc0
    "11000000", --  644 - 0x284  :  192 - 0xc0
    "11000000", --  645 - 0x285  :  192 - 0xc0
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111111", --  648 - 0x288  :  255 - 0xff -- plane 1
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11000000", --  650 - 0x28a  :  192 - 0xc0
    "11000000", --  651 - 0x28b  :  192 - 0xc0
    "11000000", --  652 - 0x28c  :  192 - 0xc0
    "11000000", --  653 - 0x28d  :  192 - 0xc0
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "00011111", --  656 - 0x290  :   31 - 0x1f -- Sprite 0x29
    "00111111", --  657 - 0x291  :   63 - 0x3f
    "00110000", --  658 - 0x292  :   48 - 0x30
    "00110000", --  659 - 0x293  :   48 - 0x30
    "00110000", --  660 - 0x294  :   48 - 0x30
    "00110000", --  661 - 0x295  :   48 - 0x30
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00011111", --  663 - 0x297  :   31 - 0x1f
    "00011111", --  664 - 0x298  :   31 - 0x1f -- plane 1
    "00111111", --  665 - 0x299  :   63 - 0x3f
    "00110000", --  666 - 0x29a  :   48 - 0x30
    "00110000", --  667 - 0x29b  :   48 - 0x30
    "00110000", --  668 - 0x29c  :   48 - 0x30
    "00110000", --  669 - 0x29d  :   48 - 0x30
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "00011111", --  671 - 0x29f  :   31 - 0x1f
    "11100011", --  672 - 0x2a0  :  227 - 0xe3 -- Sprite 0x2a
    "11110011", --  673 - 0x2a1  :  243 - 0xf3
    "01110000", --  674 - 0x2a2  :  112 - 0x70
    "01110000", --  675 - 0x2a3  :  112 - 0x70
    "01110000", --  676 - 0x2a4  :  112 - 0x70
    "01110000", --  677 - 0x2a5  :  112 - 0x70
    "11110000", --  678 - 0x2a6  :  240 - 0xf0
    "11100000", --  679 - 0x2a7  :  224 - 0xe0
    "11100011", --  680 - 0x2a8  :  227 - 0xe3 -- plane 1
    "11110011", --  681 - 0x2a9  :  243 - 0xf3
    "01110000", --  682 - 0x2aa  :  112 - 0x70
    "01110000", --  683 - 0x2ab  :  112 - 0x70
    "01110000", --  684 - 0x2ac  :  112 - 0x70
    "01110000", --  685 - 0x2ad  :  112 - 0x70
    "11110000", --  686 - 0x2ae  :  240 - 0xf0
    "11100000", --  687 - 0x2af  :  224 - 0xe0
    "11111110", --  688 - 0x2b0  :  254 - 0xfe -- Sprite 0x2b
    "11111110", --  689 - 0x2b1  :  254 - 0xfe
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "01110000", --  691 - 0x2b3  :  112 - 0x70
    "01110000", --  692 - 0x2b4  :  112 - 0x70
    "01110000", --  693 - 0x2b5  :  112 - 0x70
    "01110000", --  694 - 0x2b6  :  112 - 0x70
    "01110000", --  695 - 0x2b7  :  112 - 0x70
    "11111110", --  696 - 0x2b8  :  254 - 0xfe -- plane 1
    "11111110", --  697 - 0x2b9  :  254 - 0xfe
    "01110000", --  698 - 0x2ba  :  112 - 0x70
    "01110000", --  699 - 0x2bb  :  112 - 0x70
    "01110000", --  700 - 0x2bc  :  112 - 0x70
    "01110000", --  701 - 0x2bd  :  112 - 0x70
    "01110000", --  702 - 0x2be  :  112 - 0x70
    "01110000", --  703 - 0x2bf  :  112 - 0x70
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- plane 1
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "11111111", --  728 - 0x2d8  :  255 - 0xff -- plane 1
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00011000", --  739 - 0x2e3  :   24 - 0x18
    "00011000", --  740 - 0x2e4  :   24 - 0x18
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- plane 1
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- plane 1
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00011000", --  763 - 0x2fb  :   24 - 0x18
    "00011000", --  764 - 0x2fc  :   24 - 0x18
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00011100", --  768 - 0x300  :   28 - 0x1c -- Sprite 0x30
    "00100110", --  769 - 0x301  :   38 - 0x26
    "01100011", --  770 - 0x302  :   99 - 0x63
    "01100011", --  771 - 0x303  :   99 - 0x63
    "01100011", --  772 - 0x304  :   99 - 0x63
    "00110010", --  773 - 0x305  :   50 - 0x32
    "00011100", --  774 - 0x306  :   28 - 0x1c
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0 -- plane 1
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00001100", --  784 - 0x310  :   12 - 0xc -- Sprite 0x31
    "00011100", --  785 - 0x311  :   28 - 0x1c
    "00001100", --  786 - 0x312  :   12 - 0xc
    "00001100", --  787 - 0x313  :   12 - 0xc
    "00001100", --  788 - 0x314  :   12 - 0xc
    "00001100", --  789 - 0x315  :   12 - 0xc
    "00111111", --  790 - 0x316  :   63 - 0x3f
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- plane 1
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00111110", --  800 - 0x320  :   62 - 0x3e -- Sprite 0x32
    "01100011", --  801 - 0x321  :   99 - 0x63
    "00000111", --  802 - 0x322  :    7 - 0x7
    "00011110", --  803 - 0x323  :   30 - 0x1e
    "00111100", --  804 - 0x324  :   60 - 0x3c
    "01110000", --  805 - 0x325  :  112 - 0x70
    "01111111", --  806 - 0x326  :  127 - 0x7f
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- plane 1
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00111111", --  816 - 0x330  :   63 - 0x3f -- Sprite 0x33
    "00000110", --  817 - 0x331  :    6 - 0x6
    "00001100", --  818 - 0x332  :   12 - 0xc
    "00011110", --  819 - 0x333  :   30 - 0x1e
    "00000011", --  820 - 0x334  :    3 - 0x3
    "01100011", --  821 - 0x335  :   99 - 0x63
    "00111110", --  822 - 0x336  :   62 - 0x3e
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- plane 1
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00001110", --  832 - 0x340  :   14 - 0xe -- Sprite 0x34
    "00011110", --  833 - 0x341  :   30 - 0x1e
    "00110110", --  834 - 0x342  :   54 - 0x36
    "01100110", --  835 - 0x343  :  102 - 0x66
    "01111111", --  836 - 0x344  :  127 - 0x7f
    "00000110", --  837 - 0x345  :    6 - 0x6
    "00000110", --  838 - 0x346  :    6 - 0x6
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- plane 1
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "01111110", --  848 - 0x350  :  126 - 0x7e -- Sprite 0x35
    "01100000", --  849 - 0x351  :   96 - 0x60
    "01111110", --  850 - 0x352  :  126 - 0x7e
    "00000011", --  851 - 0x353  :    3 - 0x3
    "00000011", --  852 - 0x354  :    3 - 0x3
    "01100011", --  853 - 0x355  :   99 - 0x63
    "00111110", --  854 - 0x356  :   62 - 0x3e
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- plane 1
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00011110", --  864 - 0x360  :   30 - 0x1e -- Sprite 0x36
    "00110000", --  865 - 0x361  :   48 - 0x30
    "01100000", --  866 - 0x362  :   96 - 0x60
    "01111110", --  867 - 0x363  :  126 - 0x7e
    "01100011", --  868 - 0x364  :   99 - 0x63
    "01100011", --  869 - 0x365  :   99 - 0x63
    "00111110", --  870 - 0x366  :   62 - 0x3e
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- plane 1
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "01111111", --  880 - 0x370  :  127 - 0x7f -- Sprite 0x37
    "01100011", --  881 - 0x371  :   99 - 0x63
    "00000110", --  882 - 0x372  :    6 - 0x6
    "00001100", --  883 - 0x373  :   12 - 0xc
    "00011000", --  884 - 0x374  :   24 - 0x18
    "00011000", --  885 - 0x375  :   24 - 0x18
    "00011000", --  886 - 0x376  :   24 - 0x18
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- plane 1
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00111100", --  896 - 0x380  :   60 - 0x3c -- Sprite 0x38
    "01100010", --  897 - 0x381  :   98 - 0x62
    "01110010", --  898 - 0x382  :  114 - 0x72
    "00111100", --  899 - 0x383  :   60 - 0x3c
    "01001111", --  900 - 0x384  :   79 - 0x4f
    "01000011", --  901 - 0x385  :   67 - 0x43
    "00111110", --  902 - 0x386  :   62 - 0x3e
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- plane 1
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00111110", --  912 - 0x390  :   62 - 0x3e -- Sprite 0x39
    "01100011", --  913 - 0x391  :   99 - 0x63
    "01100011", --  914 - 0x392  :   99 - 0x63
    "00111111", --  915 - 0x393  :   63 - 0x3f
    "00000011", --  916 - 0x394  :    3 - 0x3
    "00000110", --  917 - 0x395  :    6 - 0x6
    "00111100", --  918 - 0x396  :   60 - 0x3c
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- plane 1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "01111110", --  931 - 0x3a3  :  126 - 0x7e
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x3b
    "00000010", --  945 - 0x3b1  :    2 - 0x2
    "00000100", --  946 - 0x3b2  :    4 - 0x4
    "00001000", --  947 - 0x3b3  :    8 - 0x8
    "00010000", --  948 - 0x3b4  :   16 - 0x10
    "00100000", --  949 - 0x3b5  :   32 - 0x20
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- plane 1
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000111", --  961 - 0x3c1  :    7 - 0x7
    "00011111", --  962 - 0x3c2  :   31 - 0x1f
    "00111111", --  963 - 0x3c3  :   63 - 0x3f
    "00111111", --  964 - 0x3c4  :   63 - 0x3f
    "00001111", --  965 - 0x3c5  :   15 - 0xf
    "00000011", --  966 - 0x3c6  :    3 - 0x3
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000111", --  969 - 0x3c9  :    7 - 0x7
    "00011111", --  970 - 0x3ca  :   31 - 0x1f
    "00111111", --  971 - 0x3cb  :   63 - 0x3f
    "00111111", --  972 - 0x3cc  :   63 - 0x3f
    "00001111", --  973 - 0x3cd  :   15 - 0xf
    "00000011", --  974 - 0x3ce  :    3 - 0x3
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x3d
    "11000000", --  977 - 0x3d1  :  192 - 0xc0
    "11110000", --  978 - 0x3d2  :  240 - 0xf0
    "11111000", --  979 - 0x3d3  :  248 - 0xf8
    "11111000", --  980 - 0x3d4  :  248 - 0xf8
    "11111100", --  981 - 0x3d5  :  252 - 0xfc
    "11111100", --  982 - 0x3d6  :  252 - 0xfc
    "11111100", --  983 - 0x3d7  :  252 - 0xfc
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- plane 1
    "11000000", --  985 - 0x3d9  :  192 - 0xc0
    "11110000", --  986 - 0x3da  :  240 - 0xf0
    "11111000", --  987 - 0x3db  :  248 - 0xf8
    "11111000", --  988 - 0x3dc  :  248 - 0xf8
    "11111100", --  989 - 0x3dd  :  252 - 0xfc
    "11111100", --  990 - 0x3de  :  252 - 0xfc
    "11111100", --  991 - 0x3df  :  252 - 0xfc
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000011", --  993 - 0x3e1  :    3 - 0x3
    "00001111", --  994 - 0x3e2  :   15 - 0xf
    "00111111", --  995 - 0x3e3  :   63 - 0x3f
    "00111111", --  996 - 0x3e4  :   63 - 0x3f
    "00011111", --  997 - 0x3e5  :   31 - 0x1f
    "00000111", --  998 - 0x3e6  :    7 - 0x7
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- plane 1
    "00000011", -- 1001 - 0x3e9  :    3 - 0x3
    "00001111", -- 1002 - 0x3ea  :   15 - 0xf
    "00111111", -- 1003 - 0x3eb  :   63 - 0x3f
    "00111111", -- 1004 - 0x3ec  :   63 - 0x3f
    "00011111", -- 1005 - 0x3ed  :   31 - 0x1f
    "00000111", -- 1006 - 0x3ee  :    7 - 0x7
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "11111100", -- 1008 - 0x3f0  :  252 - 0xfc -- Sprite 0x3f
    "11111100", -- 1009 - 0x3f1  :  252 - 0xfc
    "11111100", -- 1010 - 0x3f2  :  252 - 0xfc
    "11111000", -- 1011 - 0x3f3  :  248 - 0xf8
    "11111000", -- 1012 - 0x3f4  :  248 - 0xf8
    "11110000", -- 1013 - 0x3f5  :  240 - 0xf0
    "11000000", -- 1014 - 0x3f6  :  192 - 0xc0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "11111100", -- 1016 - 0x3f8  :  252 - 0xfc -- plane 1
    "11111100", -- 1017 - 0x3f9  :  252 - 0xfc
    "11111100", -- 1018 - 0x3fa  :  252 - 0xfc
    "11111000", -- 1019 - 0x3fb  :  248 - 0xf8
    "11111000", -- 1020 - 0x3fc  :  248 - 0xf8
    "11110000", -- 1021 - 0x3fd  :  240 - 0xf0
    "11000000", -- 1022 - 0x3fe  :  192 - 0xc0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x40
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- plane 1
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00011100", -- 1040 - 0x410  :   28 - 0x1c -- Sprite 0x41
    "00110110", -- 1041 - 0x411  :   54 - 0x36
    "01100011", -- 1042 - 0x412  :   99 - 0x63
    "01100011", -- 1043 - 0x413  :   99 - 0x63
    "01111111", -- 1044 - 0x414  :  127 - 0x7f
    "01100011", -- 1045 - 0x415  :   99 - 0x63
    "01100011", -- 1046 - 0x416  :   99 - 0x63
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- plane 1
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "01111110", -- 1056 - 0x420  :  126 - 0x7e -- Sprite 0x42
    "01100011", -- 1057 - 0x421  :   99 - 0x63
    "01100011", -- 1058 - 0x422  :   99 - 0x63
    "01111110", -- 1059 - 0x423  :  126 - 0x7e
    "01100011", -- 1060 - 0x424  :   99 - 0x63
    "01100011", -- 1061 - 0x425  :   99 - 0x63
    "01111110", -- 1062 - 0x426  :  126 - 0x7e
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- plane 1
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00011110", -- 1072 - 0x430  :   30 - 0x1e -- Sprite 0x43
    "00110011", -- 1073 - 0x431  :   51 - 0x33
    "01100000", -- 1074 - 0x432  :   96 - 0x60
    "01100000", -- 1075 - 0x433  :   96 - 0x60
    "01100000", -- 1076 - 0x434  :   96 - 0x60
    "00110011", -- 1077 - 0x435  :   51 - 0x33
    "00011110", -- 1078 - 0x436  :   30 - 0x1e
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- plane 1
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "01111100", -- 1088 - 0x440  :  124 - 0x7c -- Sprite 0x44
    "01100110", -- 1089 - 0x441  :  102 - 0x66
    "01100011", -- 1090 - 0x442  :   99 - 0x63
    "01100011", -- 1091 - 0x443  :   99 - 0x63
    "01100011", -- 1092 - 0x444  :   99 - 0x63
    "01100110", -- 1093 - 0x445  :  102 - 0x66
    "01111100", -- 1094 - 0x446  :  124 - 0x7c
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0 -- plane 1
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "01111111", -- 1104 - 0x450  :  127 - 0x7f -- Sprite 0x45
    "01100000", -- 1105 - 0x451  :   96 - 0x60
    "01100000", -- 1106 - 0x452  :   96 - 0x60
    "01111110", -- 1107 - 0x453  :  126 - 0x7e
    "01100000", -- 1108 - 0x454  :   96 - 0x60
    "01100000", -- 1109 - 0x455  :   96 - 0x60
    "01111111", -- 1110 - 0x456  :  127 - 0x7f
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0 -- plane 1
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "01111111", -- 1120 - 0x460  :  127 - 0x7f -- Sprite 0x46
    "01100000", -- 1121 - 0x461  :   96 - 0x60
    "01100000", -- 1122 - 0x462  :   96 - 0x60
    "01111110", -- 1123 - 0x463  :  126 - 0x7e
    "01100000", -- 1124 - 0x464  :   96 - 0x60
    "01100000", -- 1125 - 0x465  :   96 - 0x60
    "01100000", -- 1126 - 0x466  :   96 - 0x60
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0 -- plane 1
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00011111", -- 1136 - 0x470  :   31 - 0x1f -- Sprite 0x47
    "00110000", -- 1137 - 0x471  :   48 - 0x30
    "01100000", -- 1138 - 0x472  :   96 - 0x60
    "01100111", -- 1139 - 0x473  :  103 - 0x67
    "01100011", -- 1140 - 0x474  :   99 - 0x63
    "00110011", -- 1141 - 0x475  :   51 - 0x33
    "00011111", -- 1142 - 0x476  :   31 - 0x1f
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0 -- plane 1
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "01100011", -- 1152 - 0x480  :   99 - 0x63 -- Sprite 0x48
    "01100011", -- 1153 - 0x481  :   99 - 0x63
    "01100011", -- 1154 - 0x482  :   99 - 0x63
    "01111111", -- 1155 - 0x483  :  127 - 0x7f
    "01100011", -- 1156 - 0x484  :   99 - 0x63
    "01100011", -- 1157 - 0x485  :   99 - 0x63
    "01100011", -- 1158 - 0x486  :   99 - 0x63
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- plane 1
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00111111", -- 1168 - 0x490  :   63 - 0x3f -- Sprite 0x49
    "00001100", -- 1169 - 0x491  :   12 - 0xc
    "00001100", -- 1170 - 0x492  :   12 - 0xc
    "00001100", -- 1171 - 0x493  :   12 - 0xc
    "00001100", -- 1172 - 0x494  :   12 - 0xc
    "00001100", -- 1173 - 0x495  :   12 - 0xc
    "00111111", -- 1174 - 0x496  :   63 - 0x3f
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- plane 1
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000011", -- 1184 - 0x4a0  :    3 - 0x3 -- Sprite 0x4a
    "00000011", -- 1185 - 0x4a1  :    3 - 0x3
    "00000011", -- 1186 - 0x4a2  :    3 - 0x3
    "00000011", -- 1187 - 0x4a3  :    3 - 0x3
    "00000011", -- 1188 - 0x4a4  :    3 - 0x3
    "01100011", -- 1189 - 0x4a5  :   99 - 0x63
    "00111110", -- 1190 - 0x4a6  :   62 - 0x3e
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "01100011", -- 1200 - 0x4b0  :   99 - 0x63 -- Sprite 0x4b
    "01100110", -- 1201 - 0x4b1  :  102 - 0x66
    "01101100", -- 1202 - 0x4b2  :  108 - 0x6c
    "01111000", -- 1203 - 0x4b3  :  120 - 0x78
    "01111100", -- 1204 - 0x4b4  :  124 - 0x7c
    "01100110", -- 1205 - 0x4b5  :  102 - 0x66
    "01100011", -- 1206 - 0x4b6  :   99 - 0x63
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "01100000", -- 1216 - 0x4c0  :   96 - 0x60 -- Sprite 0x4c
    "01100000", -- 1217 - 0x4c1  :   96 - 0x60
    "01100000", -- 1218 - 0x4c2  :   96 - 0x60
    "01100000", -- 1219 - 0x4c3  :   96 - 0x60
    "01100000", -- 1220 - 0x4c4  :   96 - 0x60
    "01100000", -- 1221 - 0x4c5  :   96 - 0x60
    "01111111", -- 1222 - 0x4c6  :  127 - 0x7f
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "01100011", -- 1232 - 0x4d0  :   99 - 0x63 -- Sprite 0x4d
    "01110111", -- 1233 - 0x4d1  :  119 - 0x77
    "01111111", -- 1234 - 0x4d2  :  127 - 0x7f
    "01111111", -- 1235 - 0x4d3  :  127 - 0x7f
    "01101011", -- 1236 - 0x4d4  :  107 - 0x6b
    "01100011", -- 1237 - 0x4d5  :   99 - 0x63
    "01100011", -- 1238 - 0x4d6  :   99 - 0x63
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "01100011", -- 1248 - 0x4e0  :   99 - 0x63 -- Sprite 0x4e
    "01110011", -- 1249 - 0x4e1  :  115 - 0x73
    "01111011", -- 1250 - 0x4e2  :  123 - 0x7b
    "01111111", -- 1251 - 0x4e3  :  127 - 0x7f
    "01101111", -- 1252 - 0x4e4  :  111 - 0x6f
    "01100111", -- 1253 - 0x4e5  :  103 - 0x67
    "01100011", -- 1254 - 0x4e6  :   99 - 0x63
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00111110", -- 1264 - 0x4f0  :   62 - 0x3e -- Sprite 0x4f
    "01100011", -- 1265 - 0x4f1  :   99 - 0x63
    "01100011", -- 1266 - 0x4f2  :   99 - 0x63
    "01100011", -- 1267 - 0x4f3  :   99 - 0x63
    "01100011", -- 1268 - 0x4f4  :   99 - 0x63
    "01100011", -- 1269 - 0x4f5  :   99 - 0x63
    "00111110", -- 1270 - 0x4f6  :   62 - 0x3e
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "01111110", -- 1280 - 0x500  :  126 - 0x7e -- Sprite 0x50
    "01100011", -- 1281 - 0x501  :   99 - 0x63
    "01100011", -- 1282 - 0x502  :   99 - 0x63
    "01100011", -- 1283 - 0x503  :   99 - 0x63
    "01111110", -- 1284 - 0x504  :  126 - 0x7e
    "01100000", -- 1285 - 0x505  :   96 - 0x60
    "01100000", -- 1286 - 0x506  :   96 - 0x60
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- plane 1
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00111110", -- 1296 - 0x510  :   62 - 0x3e -- Sprite 0x51
    "01100011", -- 1297 - 0x511  :   99 - 0x63
    "01100011", -- 1298 - 0x512  :   99 - 0x63
    "01100011", -- 1299 - 0x513  :   99 - 0x63
    "01101111", -- 1300 - 0x514  :  111 - 0x6f
    "01100110", -- 1301 - 0x515  :  102 - 0x66
    "00111101", -- 1302 - 0x516  :   61 - 0x3d
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- plane 1
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "01111110", -- 1312 - 0x520  :  126 - 0x7e -- Sprite 0x52
    "01100011", -- 1313 - 0x521  :   99 - 0x63
    "01100011", -- 1314 - 0x522  :   99 - 0x63
    "01100111", -- 1315 - 0x523  :  103 - 0x67
    "01111100", -- 1316 - 0x524  :  124 - 0x7c
    "01101110", -- 1317 - 0x525  :  110 - 0x6e
    "01100111", -- 1318 - 0x526  :  103 - 0x67
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- plane 1
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00111100", -- 1328 - 0x530  :   60 - 0x3c -- Sprite 0x53
    "01100110", -- 1329 - 0x531  :  102 - 0x66
    "01100000", -- 1330 - 0x532  :   96 - 0x60
    "00111110", -- 1331 - 0x533  :   62 - 0x3e
    "00000011", -- 1332 - 0x534  :    3 - 0x3
    "01100011", -- 1333 - 0x535  :   99 - 0x63
    "00111110", -- 1334 - 0x536  :   62 - 0x3e
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0 -- plane 1
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00111111", -- 1344 - 0x540  :   63 - 0x3f -- Sprite 0x54
    "00001100", -- 1345 - 0x541  :   12 - 0xc
    "00001100", -- 1346 - 0x542  :   12 - 0xc
    "00001100", -- 1347 - 0x543  :   12 - 0xc
    "00001100", -- 1348 - 0x544  :   12 - 0xc
    "00001100", -- 1349 - 0x545  :   12 - 0xc
    "00001100", -- 1350 - 0x546  :   12 - 0xc
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0 -- plane 1
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "01100011", -- 1360 - 0x550  :   99 - 0x63 -- Sprite 0x55
    "01100011", -- 1361 - 0x551  :   99 - 0x63
    "01100011", -- 1362 - 0x552  :   99 - 0x63
    "01100011", -- 1363 - 0x553  :   99 - 0x63
    "01100011", -- 1364 - 0x554  :   99 - 0x63
    "01100011", -- 1365 - 0x555  :   99 - 0x63
    "00111110", -- 1366 - 0x556  :   62 - 0x3e
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- plane 1
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "01100011", -- 1376 - 0x560  :   99 - 0x63 -- Sprite 0x56
    "01100011", -- 1377 - 0x561  :   99 - 0x63
    "01100011", -- 1378 - 0x562  :   99 - 0x63
    "01110111", -- 1379 - 0x563  :  119 - 0x77
    "00111110", -- 1380 - 0x564  :   62 - 0x3e
    "00011100", -- 1381 - 0x565  :   28 - 0x1c
    "00001000", -- 1382 - 0x566  :    8 - 0x8
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- plane 1
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "01100011", -- 1392 - 0x570  :   99 - 0x63 -- Sprite 0x57
    "01100011", -- 1393 - 0x571  :   99 - 0x63
    "01101011", -- 1394 - 0x572  :  107 - 0x6b
    "01111111", -- 1395 - 0x573  :  127 - 0x7f
    "01111111", -- 1396 - 0x574  :  127 - 0x7f
    "01110111", -- 1397 - 0x575  :  119 - 0x77
    "01100011", -- 1398 - 0x576  :   99 - 0x63
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- plane 1
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "01100011", -- 1408 - 0x580  :   99 - 0x63 -- Sprite 0x58
    "01110111", -- 1409 - 0x581  :  119 - 0x77
    "00111110", -- 1410 - 0x582  :   62 - 0x3e
    "00011100", -- 1411 - 0x583  :   28 - 0x1c
    "00111110", -- 1412 - 0x584  :   62 - 0x3e
    "01110111", -- 1413 - 0x585  :  119 - 0x77
    "01100011", -- 1414 - 0x586  :   99 - 0x63
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- plane 1
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00110011", -- 1424 - 0x590  :   51 - 0x33 -- Sprite 0x59
    "00110011", -- 1425 - 0x591  :   51 - 0x33
    "00110011", -- 1426 - 0x592  :   51 - 0x33
    "00011110", -- 1427 - 0x593  :   30 - 0x1e
    "00001100", -- 1428 - 0x594  :   12 - 0xc
    "00001100", -- 1429 - 0x595  :   12 - 0xc
    "00001100", -- 1430 - 0x596  :   12 - 0xc
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0 -- plane 1
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01111111", -- 1440 - 0x5a0  :  127 - 0x7f -- Sprite 0x5a
    "00000111", -- 1441 - 0x5a1  :    7 - 0x7
    "00001110", -- 1442 - 0x5a2  :   14 - 0xe
    "00011100", -- 1443 - 0x5a3  :   28 - 0x1c
    "00111000", -- 1444 - 0x5a4  :   56 - 0x38
    "01110000", -- 1445 - 0x5a5  :  112 - 0x70
    "01111111", -- 1446 - 0x5a6  :  127 - 0x7f
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00110000", -- 1461 - 0x5b5  :   48 - 0x30
    "00110000", -- 1462 - 0x5b6  :   48 - 0x30
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0 -- Sprite 0x5c
    "11110000", -- 1473 - 0x5c1  :  240 - 0xf0
    "11111100", -- 1474 - 0x5c2  :  252 - 0xfc
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111100", -- 1476 - 0x5c4  :  252 - 0xfc
    "11110000", -- 1477 - 0x5c5  :  240 - 0xf0
    "11000000", -- 1478 - 0x5c6  :  192 - 0xc0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00111100", -- 1488 - 0x5d0  :   60 - 0x3c -- Sprite 0x5d
    "01000010", -- 1489 - 0x5d1  :   66 - 0x42
    "10011001", -- 1490 - 0x5d2  :  153 - 0x99
    "10100001", -- 1491 - 0x5d3  :  161 - 0xa1
    "10100001", -- 1492 - 0x5d4  :  161 - 0xa1
    "10011001", -- 1493 - 0x5d5  :  153 - 0x99
    "01000010", -- 1494 - 0x5d6  :   66 - 0x42
    "00111100", -- 1495 - 0x5d7  :   60 - 0x3c
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00010000", -- 1506 - 0x5e2  :   16 - 0x10
    "00010000", -- 1507 - 0x5e3  :   16 - 0x10
    "00010000", -- 1508 - 0x5e4  :   16 - 0x10
    "00010000", -- 1509 - 0x5e5  :   16 - 0x10
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00010000", -- 1514 - 0x5ea  :   16 - 0x10
    "00010000", -- 1515 - 0x5eb  :   16 - 0x10
    "00010000", -- 1516 - 0x5ec  :   16 - 0x10
    "00010000", -- 1517 - 0x5ed  :   16 - 0x10
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00110110", -- 1520 - 0x5f0  :   54 - 0x36 -- Sprite 0x5f
    "00110110", -- 1521 - 0x5f1  :   54 - 0x36
    "00010010", -- 1522 - 0x5f2  :   18 - 0x12
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000001", -- 1541 - 0x605  :    1 - 0x1
    "00011110", -- 1542 - 0x606  :   30 - 0x1e
    "00111011", -- 1543 - 0x607  :   59 - 0x3b
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- plane 1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0x61
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00001100", -- 1554 - 0x612  :   12 - 0xc
    "00111100", -- 1555 - 0x613  :   60 - 0x3c
    "11010000", -- 1556 - 0x614  :  208 - 0xd0
    "00010000", -- 1557 - 0x615  :   16 - 0x10
    "00100000", -- 1558 - 0x616  :   32 - 0x20
    "01000000", -- 1559 - 0x617  :   64 - 0x40
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- plane 1
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00111110", -- 1568 - 0x620  :   62 - 0x3e -- Sprite 0x62
    "00101101", -- 1569 - 0x621  :   45 - 0x2d
    "00110101", -- 1570 - 0x622  :   53 - 0x35
    "00011101", -- 1571 - 0x623  :   29 - 0x1d
    "00000001", -- 1572 - 0x624  :    1 - 0x1
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- plane 1
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "10110000", -- 1584 - 0x630  :  176 - 0xb0 -- Sprite 0x63
    "10111000", -- 1585 - 0x631  :  184 - 0xb8
    "11111000", -- 1586 - 0x632  :  248 - 0xf8
    "01111000", -- 1587 - 0x633  :  120 - 0x78
    "10011000", -- 1588 - 0x634  :  152 - 0x98
    "11110000", -- 1589 - 0x635  :  240 - 0xf0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0 -- plane 1
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000111", -- 1602 - 0x642  :    7 - 0x7
    "00000011", -- 1603 - 0x643  :    3 - 0x3
    "00001101", -- 1604 - 0x644  :   13 - 0xd
    "00011110", -- 1605 - 0x645  :   30 - 0x1e
    "00010111", -- 1606 - 0x646  :   23 - 0x17
    "00011101", -- 1607 - 0x647  :   29 - 0x1d
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- plane 1
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "10000000", -- 1617 - 0x651  :  128 - 0x80
    "01110000", -- 1618 - 0x652  :  112 - 0x70
    "11100000", -- 1619 - 0x653  :  224 - 0xe0
    "11011000", -- 1620 - 0x654  :  216 - 0xd8
    "10111100", -- 1621 - 0x655  :  188 - 0xbc
    "01110100", -- 1622 - 0x656  :  116 - 0x74
    "11011100", -- 1623 - 0x657  :  220 - 0xdc
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- plane 1
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00011111", -- 1632 - 0x660  :   31 - 0x1f -- Sprite 0x66
    "00001011", -- 1633 - 0x661  :   11 - 0xb
    "00001111", -- 1634 - 0x662  :   15 - 0xf
    "00000101", -- 1635 - 0x663  :    5 - 0x5
    "00000011", -- 1636 - 0x664  :    3 - 0x3
    "00000001", -- 1637 - 0x665  :    1 - 0x1
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- plane 1
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11111100", -- 1648 - 0x670  :  252 - 0xfc -- Sprite 0x67
    "01101000", -- 1649 - 0x671  :  104 - 0x68
    "11111000", -- 1650 - 0x672  :  248 - 0xf8
    "10110000", -- 1651 - 0x673  :  176 - 0xb0
    "11100000", -- 1652 - 0x674  :  224 - 0xe0
    "10000000", -- 1653 - 0x675  :  128 - 0x80
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- plane 1
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- plane 1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000001", -- 1675 - 0x68b  :    1 - 0x1
    "00000001", -- 1676 - 0x68c  :    1 - 0x1
    "00001011", -- 1677 - 0x68d  :   11 - 0xb
    "00011100", -- 1678 - 0x68e  :   28 - 0x1c
    "00111111", -- 1679 - 0x68f  :   63 - 0x3f
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0 -- plane 1
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00110000", -- 1690 - 0x69a  :   48 - 0x30
    "01111000", -- 1691 - 0x69b  :  120 - 0x78
    "10000000", -- 1692 - 0x69c  :  128 - 0x80
    "11110000", -- 1693 - 0x69d  :  240 - 0xf0
    "11111000", -- 1694 - 0x69e  :  248 - 0xf8
    "11111100", -- 1695 - 0x69f  :  252 - 0xfc
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00111111", -- 1704 - 0x6a8  :   63 - 0x3f -- plane 1
    "00111111", -- 1705 - 0x6a9  :   63 - 0x3f
    "00111111", -- 1706 - 0x6aa  :   63 - 0x3f
    "00011111", -- 1707 - 0x6ab  :   31 - 0x1f
    "00011111", -- 1708 - 0x6ac  :   31 - 0x1f
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0x6b
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "11111100", -- 1720 - 0x6b8  :  252 - 0xfc -- plane 1
    "11101100", -- 1721 - 0x6b9  :  236 - 0xec
    "11101100", -- 1722 - 0x6ba  :  236 - 0xec
    "11011000", -- 1723 - 0x6bb  :  216 - 0xd8
    "11111000", -- 1724 - 0x6bc  :  248 - 0xf8
    "11100000", -- 1725 - 0x6bd  :  224 - 0xe0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0x6c
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000001", -- 1730 - 0x6c2  :    1 - 0x1
    "00011101", -- 1731 - 0x6c3  :   29 - 0x1d
    "00111110", -- 1732 - 0x6c4  :   62 - 0x3e
    "00111111", -- 1733 - 0x6c5  :   63 - 0x3f
    "00111111", -- 1734 - 0x6c6  :   63 - 0x3f
    "00111111", -- 1735 - 0x6c7  :   63 - 0x3f
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000001", -- 1738 - 0x6ca  :    1 - 0x1
    "00011101", -- 1739 - 0x6cb  :   29 - 0x1d
    "00111110", -- 1740 - 0x6cc  :   62 - 0x3e
    "00111111", -- 1741 - 0x6cd  :   63 - 0x3f
    "00111111", -- 1742 - 0x6ce  :   63 - 0x3f
    "00111111", -- 1743 - 0x6cf  :   63 - 0x3f
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0x6d
    "10000000", -- 1745 - 0x6d1  :  128 - 0x80
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "01110000", -- 1747 - 0x6d3  :  112 - 0x70
    "11111000", -- 1748 - 0x6d4  :  248 - 0xf8
    "11111100", -- 1749 - 0x6d5  :  252 - 0xfc
    "11111100", -- 1750 - 0x6d6  :  252 - 0xfc
    "11111100", -- 1751 - 0x6d7  :  252 - 0xfc
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- plane 1
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "01110000", -- 1755 - 0x6db  :  112 - 0x70
    "11111000", -- 1756 - 0x6dc  :  248 - 0xf8
    "11111100", -- 1757 - 0x6dd  :  252 - 0xfc
    "11111100", -- 1758 - 0x6de  :  252 - 0xfc
    "11111100", -- 1759 - 0x6df  :  252 - 0xfc
    "00111111", -- 1760 - 0x6e0  :   63 - 0x3f -- Sprite 0x6e
    "00111111", -- 1761 - 0x6e1  :   63 - 0x3f
    "00011111", -- 1762 - 0x6e2  :   31 - 0x1f
    "00011111", -- 1763 - 0x6e3  :   31 - 0x1f
    "00001111", -- 1764 - 0x6e4  :   15 - 0xf
    "00000110", -- 1765 - 0x6e5  :    6 - 0x6
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00111111", -- 1768 - 0x6e8  :   63 - 0x3f -- plane 1
    "00111111", -- 1769 - 0x6e9  :   63 - 0x3f
    "00011111", -- 1770 - 0x6ea  :   31 - 0x1f
    "00011111", -- 1771 - 0x6eb  :   31 - 0x1f
    "00001111", -- 1772 - 0x6ec  :   15 - 0xf
    "00000110", -- 1773 - 0x6ed  :    6 - 0x6
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11101100", -- 1776 - 0x6f0  :  236 - 0xec -- Sprite 0x6f
    "11101100", -- 1777 - 0x6f1  :  236 - 0xec
    "11011000", -- 1778 - 0x6f2  :  216 - 0xd8
    "11111000", -- 1779 - 0x6f3  :  248 - 0xf8
    "11110000", -- 1780 - 0x6f4  :  240 - 0xf0
    "11100000", -- 1781 - 0x6f5  :  224 - 0xe0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "11101100", -- 1784 - 0x6f8  :  236 - 0xec -- plane 1
    "11101100", -- 1785 - 0x6f9  :  236 - 0xec
    "11011000", -- 1786 - 0x6fa  :  216 - 0xd8
    "11111000", -- 1787 - 0x6fb  :  248 - 0xf8
    "11110000", -- 1788 - 0x6fc  :  240 - 0xf0
    "11100000", -- 1789 - 0x6fd  :  224 - 0xe0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0x70
    "00000100", -- 1793 - 0x701  :    4 - 0x4
    "00000011", -- 1794 - 0x702  :    3 - 0x3
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000001", -- 1796 - 0x704  :    1 - 0x1
    "00000111", -- 1797 - 0x705  :    7 - 0x7
    "00001111", -- 1798 - 0x706  :   15 - 0xf
    "00001100", -- 1799 - 0x707  :   12 - 0xc
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- plane 1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0x71
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "11100000", -- 1810 - 0x712  :  224 - 0xe0
    "10000000", -- 1811 - 0x713  :  128 - 0x80
    "01000000", -- 1812 - 0x714  :   64 - 0x40
    "11110000", -- 1813 - 0x715  :  240 - 0xf0
    "10011000", -- 1814 - 0x716  :  152 - 0x98
    "11111000", -- 1815 - 0x717  :  248 - 0xf8
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- plane 1
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00011111", -- 1824 - 0x720  :   31 - 0x1f -- Sprite 0x72
    "00010011", -- 1825 - 0x721  :   19 - 0x13
    "00011111", -- 1826 - 0x722  :   31 - 0x1f
    "00001111", -- 1827 - 0x723  :   15 - 0xf
    "00001001", -- 1828 - 0x724  :    9 - 0x9
    "00000111", -- 1829 - 0x725  :    7 - 0x7
    "00000001", -- 1830 - 0x726  :    1 - 0x1
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- plane 1
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "11100100", -- 1840 - 0x730  :  228 - 0xe4 -- Sprite 0x73
    "00111100", -- 1841 - 0x731  :   60 - 0x3c
    "11100100", -- 1842 - 0x732  :  228 - 0xe4
    "00111000", -- 1843 - 0x733  :   56 - 0x38
    "11111000", -- 1844 - 0x734  :  248 - 0xf8
    "11110000", -- 1845 - 0x735  :  240 - 0xf0
    "11000000", -- 1846 - 0x736  :  192 - 0xc0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- plane 1
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0x74
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- plane 1
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00010001", -- 1868 - 0x74c  :   17 - 0x11
    "00010011", -- 1869 - 0x74d  :   19 - 0x13
    "00011111", -- 1870 - 0x74e  :   31 - 0x1f
    "00011111", -- 1871 - 0x74f  :   31 - 0x1f
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0x75
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- plane 1
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "10000000", -- 1883 - 0x75b  :  128 - 0x80
    "11000100", -- 1884 - 0x75c  :  196 - 0xc4
    "11100100", -- 1885 - 0x75d  :  228 - 0xe4
    "11111100", -- 1886 - 0x75e  :  252 - 0xfc
    "11111100", -- 1887 - 0x75f  :  252 - 0xfc
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0x76
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00011111", -- 1896 - 0x768  :   31 - 0x1f -- plane 1
    "00001110", -- 1897 - 0x769  :   14 - 0xe
    "00000110", -- 1898 - 0x76a  :    6 - 0x6
    "00000010", -- 1899 - 0x76b  :    2 - 0x2
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0x77
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "11111100", -- 1912 - 0x778  :  252 - 0xfc -- plane 1
    "10111000", -- 1913 - 0x779  :  184 - 0xb8
    "10110000", -- 1914 - 0x77a  :  176 - 0xb0
    "10100000", -- 1915 - 0x77b  :  160 - 0xa0
    "10000000", -- 1916 - 0x77c  :  128 - 0x80
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- plane 1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000001", -- 1931 - 0x78b  :    1 - 0x1
    "00000011", -- 1932 - 0x78c  :    3 - 0x3
    "00000110", -- 1933 - 0x78d  :    6 - 0x6
    "00000110", -- 1934 - 0x78e  :    6 - 0x6
    "00001111", -- 1935 - 0x78f  :   15 - 0xf
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0x79
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- plane 1
    "00011000", -- 1945 - 0x799  :   24 - 0x18
    "11110100", -- 1946 - 0x79a  :  244 - 0xf4
    "11111000", -- 1947 - 0x79b  :  248 - 0xf8
    "00111000", -- 1948 - 0x79c  :   56 - 0x38
    "01111100", -- 1949 - 0x79d  :  124 - 0x7c
    "11111100", -- 1950 - 0x79e  :  252 - 0xfc
    "11111100", -- 1951 - 0x79f  :  252 - 0xfc
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00001111", -- 1960 - 0x7a8  :   15 - 0xf -- plane 1
    "00011111", -- 1961 - 0x7a9  :   31 - 0x1f
    "00110000", -- 1962 - 0x7aa  :   48 - 0x30
    "00111000", -- 1963 - 0x7ab  :   56 - 0x38
    "00011101", -- 1964 - 0x7ac  :   29 - 0x1d
    "00000011", -- 1965 - 0x7ad  :    3 - 0x3
    "00000011", -- 1966 - 0x7ae  :    3 - 0x3
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0x7b
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "11111100", -- 1976 - 0x7b8  :  252 - 0xfc -- plane 1
    "11111100", -- 1977 - 0x7b9  :  252 - 0xfc
    "01111100", -- 1978 - 0x7ba  :  124 - 0x7c
    "10001110", -- 1979 - 0x7bb  :  142 - 0x8e
    "10000110", -- 1980 - 0x7bc  :  134 - 0x86
    "10011100", -- 1981 - 0x7bd  :  156 - 0x9c
    "01111000", -- 1982 - 0x7be  :  120 - 0x78
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0x7c
    "00000001", -- 1985 - 0x7c1  :    1 - 0x1
    "00000110", -- 1986 - 0x7c2  :    6 - 0x6
    "00000111", -- 1987 - 0x7c3  :    7 - 0x7
    "00000111", -- 1988 - 0x7c4  :    7 - 0x7
    "00000111", -- 1989 - 0x7c5  :    7 - 0x7
    "00000001", -- 1990 - 0x7c6  :    1 - 0x1
    "00000011", -- 1991 - 0x7c7  :    3 - 0x3
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "00000001", -- 1993 - 0x7c9  :    1 - 0x1
    "00000110", -- 1994 - 0x7ca  :    6 - 0x6
    "00000111", -- 1995 - 0x7cb  :    7 - 0x7
    "00000111", -- 1996 - 0x7cc  :    7 - 0x7
    "00000111", -- 1997 - 0x7cd  :    7 - 0x7
    "00000001", -- 1998 - 0x7ce  :    1 - 0x1
    "00000011", -- 1999 - 0x7cf  :    3 - 0x3
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0x7d
    "11000000", -- 2001 - 0x7d1  :  192 - 0xc0
    "00110000", -- 2002 - 0x7d2  :   48 - 0x30
    "11110000", -- 2003 - 0x7d3  :  240 - 0xf0
    "11110000", -- 2004 - 0x7d4  :  240 - 0xf0
    "11110000", -- 2005 - 0x7d5  :  240 - 0xf0
    "01000000", -- 2006 - 0x7d6  :   64 - 0x40
    "01000000", -- 2007 - 0x7d7  :   64 - 0x40
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- plane 1
    "11000000", -- 2009 - 0x7d9  :  192 - 0xc0
    "00110000", -- 2010 - 0x7da  :   48 - 0x30
    "11110000", -- 2011 - 0x7db  :  240 - 0xf0
    "11110000", -- 2012 - 0x7dc  :  240 - 0xf0
    "11110000", -- 2013 - 0x7dd  :  240 - 0xf0
    "01000000", -- 2014 - 0x7de  :   64 - 0x40
    "01000000", -- 2015 - 0x7df  :   64 - 0x40
    "00000001", -- 2016 - 0x7e0  :    1 - 0x1 -- Sprite 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000001", -- 2018 - 0x7e2  :    1 - 0x1
    "00000011", -- 2019 - 0x7e3  :    3 - 0x3
    "00000001", -- 2020 - 0x7e4  :    1 - 0x1
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000001", -- 2024 - 0x7e8  :    1 - 0x1 -- plane 1
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000001", -- 2026 - 0x7ea  :    1 - 0x1
    "00000011", -- 2027 - 0x7eb  :    3 - 0x3
    "00000001", -- 2028 - 0x7ec  :    1 - 0x1
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "01000000", -- 2032 - 0x7f0  :   64 - 0x40 -- Sprite 0x7f
    "01000000", -- 2033 - 0x7f1  :   64 - 0x40
    "01000000", -- 2034 - 0x7f2  :   64 - 0x40
    "01000000", -- 2035 - 0x7f3  :   64 - 0x40
    "01000000", -- 2036 - 0x7f4  :   64 - 0x40
    "10000000", -- 2037 - 0x7f5  :  128 - 0x80
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "01000000", -- 2040 - 0x7f8  :   64 - 0x40 -- plane 1
    "01000000", -- 2041 - 0x7f9  :   64 - 0x40
    "01000000", -- 2042 - 0x7fa  :   64 - 0x40
    "01000000", -- 2043 - 0x7fb  :   64 - 0x40
    "01000000", -- 2044 - 0x7fc  :   64 - 0x40
    "10000000", -- 2045 - 0x7fd  :  128 - 0x80
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "11111111", -- 2048 - 0x800  :  255 - 0xff -- Sprite 0x80
    "11111111", -- 2049 - 0x801  :  255 - 0xff
    "11111111", -- 2050 - 0x802  :  255 - 0xff
    "11111111", -- 2051 - 0x803  :  255 - 0xff
    "11000000", -- 2052 - 0x804  :  192 - 0xc0
    "11000000", -- 2053 - 0x805  :  192 - 0xc0
    "11000000", -- 2054 - 0x806  :  192 - 0xc0
    "11000111", -- 2055 - 0x807  :  199 - 0xc7
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- plane 1
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000000", -- 2059 - 0x80b  :    0 - 0x0
    "00000000", -- 2060 - 0x80c  :    0 - 0x0
    "00011111", -- 2061 - 0x80d  :   31 - 0x1f
    "00010000", -- 2062 - 0x80e  :   16 - 0x10
    "00010111", -- 2063 - 0x80f  :   23 - 0x17
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Sprite 0x81
    "11111111", -- 2065 - 0x811  :  255 - 0xff
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "11111111", -- 2067 - 0x813  :  255 - 0xff
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "11111111", -- 2071 - 0x817  :  255 - 0xff
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- plane 1
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00000000", -- 2075 - 0x81b  :    0 - 0x0
    "00000000", -- 2076 - 0x81c  :    0 - 0x0
    "11111111", -- 2077 - 0x81d  :  255 - 0xff
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "11111111", -- 2079 - 0x81f  :  255 - 0xff
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Sprite 0x82
    "11111111", -- 2081 - 0x821  :  255 - 0xff
    "11111111", -- 2082 - 0x822  :  255 - 0xff
    "11111111", -- 2083 - 0x823  :  255 - 0xff
    "01111111", -- 2084 - 0x824  :  127 - 0x7f
    "00111111", -- 2085 - 0x825  :   63 - 0x3f
    "00011111", -- 2086 - 0x826  :   31 - 0x1f
    "11001111", -- 2087 - 0x827  :  207 - 0xcf
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- plane 1
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "00000000", -- 2092 - 0x82c  :    0 - 0x0
    "10000000", -- 2093 - 0x82d  :  128 - 0x80
    "00000000", -- 2094 - 0x82e  :    0 - 0x0
    "11000000", -- 2095 - 0x82f  :  192 - 0xc0
    "11111111", -- 2096 - 0x830  :  255 - 0xff -- Sprite 0x83
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "11111111", -- 2098 - 0x832  :  255 - 0xff
    "11110111", -- 2099 - 0x833  :  247 - 0xf7
    "11110111", -- 2100 - 0x834  :  247 - 0xf7
    "11100010", -- 2101 - 0x835  :  226 - 0xe2
    "11100000", -- 2102 - 0x836  :  224 - 0xe0
    "11000110", -- 2103 - 0x837  :  198 - 0xc6
    "00000000", -- 2104 - 0x838  :    0 - 0x0 -- plane 1
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00001000", -- 2109 - 0x83d  :    8 - 0x8
    "00001000", -- 2110 - 0x83e  :    8 - 0x8
    "00010110", -- 2111 - 0x83f  :   22 - 0x16
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Sprite 0x84
    "11111111", -- 2113 - 0x841  :  255 - 0xff
    "11111111", -- 2114 - 0x842  :  255 - 0xff
    "11111111", -- 2115 - 0x843  :  255 - 0xff
    "10111111", -- 2116 - 0x844  :  191 - 0xbf
    "10111111", -- 2117 - 0x845  :  191 - 0xbf
    "00011111", -- 2118 - 0x846  :   31 - 0x1f
    "00011111", -- 2119 - 0x847  :   31 - 0x1f
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- plane 1
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "00000000", -- 2124 - 0x84c  :    0 - 0x0
    "00000000", -- 2125 - 0x84d  :    0 - 0x0
    "01000000", -- 2126 - 0x84e  :   64 - 0x40
    "11000000", -- 2127 - 0x84f  :  192 - 0xc0
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Sprite 0x85
    "11111111", -- 2129 - 0x851  :  255 - 0xff
    "11111111", -- 2130 - 0x852  :  255 - 0xff
    "11111111", -- 2131 - 0x853  :  255 - 0xff
    "11111110", -- 2132 - 0x854  :  254 - 0xfe
    "11111000", -- 2133 - 0x855  :  248 - 0xf8
    "11100000", -- 2134 - 0x856  :  224 - 0xe0
    "11000000", -- 2135 - 0x857  :  192 - 0xc0
    "00000000", -- 2136 - 0x858  :    0 - 0x0 -- plane 1
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000001", -- 2141 - 0x85d  :    1 - 0x1
    "00000111", -- 2142 - 0x85e  :    7 - 0x7
    "00001100", -- 2143 - 0x85f  :   12 - 0xc
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11111111", -- 2147 - 0x863  :  255 - 0xff
    "00000111", -- 2148 - 0x864  :    7 - 0x7
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00111111", -- 2150 - 0x866  :   63 - 0x3f
    "11111111", -- 2151 - 0x867  :  255 - 0xff
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- plane 1
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "11000000", -- 2157 - 0x86d  :  192 - 0xc0
    "00111111", -- 2158 - 0x86e  :   63 - 0x3f
    "11111111", -- 2159 - 0x86f  :  255 - 0xff
    "11111111", -- 2160 - 0x870  :  255 - 0xff -- Sprite 0x87
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "11111111", -- 2165 - 0x875  :  255 - 0xff
    "00111111", -- 2166 - 0x876  :   63 - 0x3f
    "11001111", -- 2167 - 0x877  :  207 - 0xcf
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- plane 1
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "11000000", -- 2175 - 0x87f  :  192 - 0xc0
    "11111111", -- 2176 - 0x880  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "11111111", -- 2178 - 0x882  :  255 - 0xff
    "11111111", -- 2179 - 0x883  :  255 - 0xff
    "11111111", -- 2180 - 0x884  :  255 - 0xff
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "11111111", -- 2182 - 0x886  :  255 - 0xff
    "11111111", -- 2183 - 0x887  :  255 - 0xff
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "00000000", -- 2190 - 0x88e  :    0 - 0x0
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "11111111", -- 2192 - 0x890  :  255 - 0xff -- Sprite 0x89
    "11111111", -- 2193 - 0x891  :  255 - 0xff
    "11111111", -- 2194 - 0x892  :  255 - 0xff
    "01110111", -- 2195 - 0x893  :  119 - 0x77
    "00010011", -- 2196 - 0x894  :   19 - 0x13
    "00000001", -- 2197 - 0x895  :    1 - 0x1
    "00010000", -- 2198 - 0x896  :   16 - 0x10
    "00011000", -- 2199 - 0x897  :   24 - 0x18
    "00000000", -- 2200 - 0x898  :    0 - 0x0 -- plane 1
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000000", -- 2203 - 0x89b  :    0 - 0x0
    "00000000", -- 2204 - 0x89c  :    0 - 0x0
    "01000100", -- 2205 - 0x89d  :   68 - 0x44
    "01010110", -- 2206 - 0x89e  :   86 - 0x56
    "01011011", -- 2207 - 0x89f  :   91 - 0x5b
    "11111111", -- 2208 - 0x8a0  :  255 - 0xff -- Sprite 0x8a
    "11111111", -- 2209 - 0x8a1  :  255 - 0xff
    "11111111", -- 2210 - 0x8a2  :  255 - 0xff
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "11111111", -- 2212 - 0x8a4  :  255 - 0xff
    "11111111", -- 2213 - 0x8a5  :  255 - 0xff
    "11111111", -- 2214 - 0x8a6  :  255 - 0xff
    "01111111", -- 2215 - 0x8a7  :  127 - 0x7f
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00000000", -- 2222 - 0x8ae  :    0 - 0x0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "11111111", -- 2224 - 0x8b0  :  255 - 0xff -- Sprite 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11111111", -- 2226 - 0x8b2  :  255 - 0xff
    "11110111", -- 2227 - 0x8b3  :  247 - 0xf7
    "11100101", -- 2228 - 0x8b4  :  229 - 0xe5
    "11000001", -- 2229 - 0x8b5  :  193 - 0xc1
    "10000100", -- 2230 - 0x8b6  :  132 - 0x84
    "00001100", -- 2231 - 0x8b7  :   12 - 0xc
    "00000000", -- 2232 - 0x8b8  :    0 - 0x0 -- plane 1
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00000000", -- 2234 - 0x8ba  :    0 - 0x0
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00000000", -- 2236 - 0x8bc  :    0 - 0x0
    "00010000", -- 2237 - 0x8bd  :   16 - 0x10
    "00110100", -- 2238 - 0x8be  :   52 - 0x34
    "01101101", -- 2239 - 0x8bf  :  109 - 0x6d
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Sprite 0x8c
    "11111111", -- 2241 - 0x8c1  :  255 - 0xff
    "11111111", -- 2242 - 0x8c2  :  255 - 0xff
    "11111111", -- 2243 - 0x8c3  :  255 - 0xff
    "11111111", -- 2244 - 0x8c4  :  255 - 0xff
    "01111111", -- 2245 - 0x8c5  :  127 - 0x7f
    "01111110", -- 2246 - 0x8c6  :  126 - 0x7e
    "01111110", -- 2247 - 0x8c7  :  126 - 0x7e
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "11111111", -- 2256 - 0x8d0  :  255 - 0xff -- Sprite 0x8d
    "11111111", -- 2257 - 0x8d1  :  255 - 0xff
    "10111111", -- 2258 - 0x8d2  :  191 - 0xbf
    "10110111", -- 2259 - 0x8d3  :  183 - 0xb7
    "00010111", -- 2260 - 0x8d4  :   23 - 0x17
    "00000011", -- 2261 - 0x8d5  :    3 - 0x3
    "00100011", -- 2262 - 0x8d6  :   35 - 0x23
    "00100001", -- 2263 - 0x8d7  :   33 - 0x21
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- plane 1
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "00000000", -- 2267 - 0x8db  :    0 - 0x0
    "01000000", -- 2268 - 0x8dc  :   64 - 0x40
    "01001000", -- 2269 - 0x8dd  :   72 - 0x48
    "10101000", -- 2270 - 0x8de  :  168 - 0xa8
    "10101100", -- 2271 - 0x8df  :  172 - 0xac
    "11111111", -- 2272 - 0x8e0  :  255 - 0xff -- Sprite 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11111011", -- 2274 - 0x8e2  :  251 - 0xfb
    "11111001", -- 2275 - 0x8e3  :  249 - 0xf9
    "11111000", -- 2276 - 0x8e4  :  248 - 0xf8
    "11111000", -- 2277 - 0x8e5  :  248 - 0xf8
    "11111000", -- 2278 - 0x8e6  :  248 - 0xf8
    "11111000", -- 2279 - 0x8e7  :  248 - 0xf8
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "00000000", -- 2283 - 0x8eb  :    0 - 0x0
    "00000010", -- 2284 - 0x8ec  :    2 - 0x2
    "00000010", -- 2285 - 0x8ed  :    2 - 0x2
    "00000010", -- 2286 - 0x8ee  :    2 - 0x2
    "00000010", -- 2287 - 0x8ef  :    2 - 0x2
    "11111111", -- 2288 - 0x8f0  :  255 - 0xff -- Sprite 0x8f
    "11111111", -- 2289 - 0x8f1  :  255 - 0xff
    "01111000", -- 2290 - 0x8f2  :  120 - 0x78
    "00111000", -- 2291 - 0x8f3  :   56 - 0x38
    "00011000", -- 2292 - 0x8f4  :   24 - 0x18
    "00001000", -- 2293 - 0x8f5  :    8 - 0x8
    "10000000", -- 2294 - 0x8f6  :  128 - 0x80
    "11000000", -- 2295 - 0x8f7  :  192 - 0xc0
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0 -- plane 1
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00000000", -- 2298 - 0x8fa  :    0 - 0x0
    "00000011", -- 2299 - 0x8fb  :    3 - 0x3
    "01000011", -- 2300 - 0x8fc  :   67 - 0x43
    "01100010", -- 2301 - 0x8fd  :   98 - 0x62
    "10110010", -- 2302 - 0x8fe  :  178 - 0xb2
    "11011010", -- 2303 - 0x8ff  :  218 - 0xda
    "11111111", -- 2304 - 0x900  :  255 - 0xff -- Sprite 0x90
    "11111111", -- 2305 - 0x901  :  255 - 0xff
    "00000001", -- 2306 - 0x902  :    1 - 0x1
    "00000001", -- 2307 - 0x903  :    1 - 0x1
    "00000001", -- 2308 - 0x904  :    1 - 0x1
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "11111111", -- 2310 - 0x906  :  255 - 0xff
    "11111111", -- 2311 - 0x907  :  255 - 0xff
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- plane 1
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "11111100", -- 2315 - 0x90b  :  252 - 0xfc
    "11111100", -- 2316 - 0x90c  :  252 - 0xfc
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "11111111", -- 2318 - 0x90e  :  255 - 0xff
    "11111111", -- 2319 - 0x90f  :  255 - 0xff
    "11111111", -- 2320 - 0x910  :  255 - 0xff -- Sprite 0x91
    "11111111", -- 2321 - 0x911  :  255 - 0xff
    "11111111", -- 2322 - 0x912  :  255 - 0xff
    "11111111", -- 2323 - 0x913  :  255 - 0xff
    "11111111", -- 2324 - 0x914  :  255 - 0xff
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "01111111", -- 2326 - 0x916  :  127 - 0x7f
    "00111111", -- 2327 - 0x917  :   63 - 0x3f
    "00000000", -- 2328 - 0x918  :    0 - 0x0 -- plane 1
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00000000", -- 2331 - 0x91b  :    0 - 0x0
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "11000111", -- 2336 - 0x920  :  199 - 0xc7 -- Sprite 0x92
    "11000111", -- 2337 - 0x921  :  199 - 0xc7
    "11000111", -- 2338 - 0x922  :  199 - 0xc7
    "11000111", -- 2339 - 0x923  :  199 - 0xc7
    "11000111", -- 2340 - 0x924  :  199 - 0xc7
    "11000111", -- 2341 - 0x925  :  199 - 0xc7
    "11000111", -- 2342 - 0x926  :  199 - 0xc7
    "11000111", -- 2343 - 0x927  :  199 - 0xc7
    "00010111", -- 2344 - 0x928  :   23 - 0x17 -- plane 1
    "00010111", -- 2345 - 0x929  :   23 - 0x17
    "00010111", -- 2346 - 0x92a  :   23 - 0x17
    "00010111", -- 2347 - 0x92b  :   23 - 0x17
    "00010111", -- 2348 - 0x92c  :   23 - 0x17
    "00010111", -- 2349 - 0x92d  :   23 - 0x17
    "00010111", -- 2350 - 0x92e  :   23 - 0x17
    "00010111", -- 2351 - 0x92f  :   23 - 0x17
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Sprite 0x93
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "11111111", -- 2354 - 0x932  :  255 - 0xff
    "11111111", -- 2355 - 0x933  :  255 - 0xff
    "11111001", -- 2356 - 0x934  :  249 - 0xf9
    "11111001", -- 2357 - 0x935  :  249 - 0xf9
    "11111111", -- 2358 - 0x936  :  255 - 0xff
    "11111111", -- 2359 - 0x937  :  255 - 0xff
    "11111111", -- 2360 - 0x938  :  255 - 0xff -- plane 1
    "11111111", -- 2361 - 0x939  :  255 - 0xff
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "11111111", -- 2363 - 0x93b  :  255 - 0xff
    "11111001", -- 2364 - 0x93c  :  249 - 0xf9
    "11111001", -- 2365 - 0x93d  :  249 - 0xf9
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "11111111", -- 2367 - 0x93f  :  255 - 0xff
    "11110111", -- 2368 - 0x940  :  247 - 0xf7 -- Sprite 0x94
    "11111011", -- 2369 - 0x941  :  251 - 0xfb
    "11111011", -- 2370 - 0x942  :  251 - 0xfb
    "11111101", -- 2371 - 0x943  :  253 - 0xfd
    "11111100", -- 2372 - 0x944  :  252 - 0xfc
    "11111100", -- 2373 - 0x945  :  252 - 0xfc
    "01111100", -- 2374 - 0x946  :  124 - 0x7c
    "01111100", -- 2375 - 0x947  :  124 - 0x7c
    "11110000", -- 2376 - 0x948  :  240 - 0xf0 -- plane 1
    "11111000", -- 2377 - 0x949  :  248 - 0xf8
    "11111000", -- 2378 - 0x94a  :  248 - 0xf8
    "11111100", -- 2379 - 0x94b  :  252 - 0xfc
    "11111100", -- 2380 - 0x94c  :  252 - 0xfc
    "11111100", -- 2381 - 0x94d  :  252 - 0xfc
    "01111100", -- 2382 - 0x94e  :  124 - 0x7c
    "01111100", -- 2383 - 0x94f  :  124 - 0x7c
    "11000111", -- 2384 - 0x950  :  199 - 0xc7 -- Sprite 0x95
    "10001111", -- 2385 - 0x951  :  143 - 0x8f
    "10001111", -- 2386 - 0x952  :  143 - 0x8f
    "00011111", -- 2387 - 0x953  :   31 - 0x1f
    "00011111", -- 2388 - 0x954  :   31 - 0x1f
    "00111111", -- 2389 - 0x955  :   63 - 0x3f
    "00111111", -- 2390 - 0x956  :   63 - 0x3f
    "01111111", -- 2391 - 0x957  :  127 - 0x7f
    "00010111", -- 2392 - 0x958  :   23 - 0x17 -- plane 1
    "00101111", -- 2393 - 0x959  :   47 - 0x2f
    "00101111", -- 2394 - 0x95a  :   47 - 0x2f
    "01011111", -- 2395 - 0x95b  :   95 - 0x5f
    "01011111", -- 2396 - 0x95c  :   95 - 0x5f
    "10111111", -- 2397 - 0x95d  :  191 - 0xbf
    "10111111", -- 2398 - 0x95e  :  191 - 0xbf
    "01111111", -- 2399 - 0x95f  :  127 - 0x7f
    "00001111", -- 2400 - 0x960  :   15 - 0xf -- Sprite 0x96
    "00001111", -- 2401 - 0x961  :   15 - 0xf
    "10000111", -- 2402 - 0x962  :  135 - 0x87
    "10000111", -- 2403 - 0x963  :  135 - 0x87
    "11000010", -- 2404 - 0x964  :  194 - 0xc2
    "11000010", -- 2405 - 0x965  :  194 - 0xc2
    "11100000", -- 2406 - 0x966  :  224 - 0xe0
    "11100000", -- 2407 - 0x967  :  224 - 0xe0
    "01100000", -- 2408 - 0x968  :   96 - 0x60 -- plane 1
    "01100000", -- 2409 - 0x969  :   96 - 0x60
    "10110000", -- 2410 - 0x96a  :  176 - 0xb0
    "10110000", -- 2411 - 0x96b  :  176 - 0xb0
    "11011000", -- 2412 - 0x96c  :  216 - 0xd8
    "11011000", -- 2413 - 0x96d  :  216 - 0xd8
    "11101100", -- 2414 - 0x96e  :  236 - 0xec
    "11101100", -- 2415 - 0x96f  :  236 - 0xec
    "10000011", -- 2416 - 0x970  :  131 - 0x83 -- Sprite 0x97
    "10001111", -- 2417 - 0x971  :  143 - 0x8f
    "00001111", -- 2418 - 0x972  :   15 - 0xf
    "00011111", -- 2419 - 0x973  :   31 - 0x1f
    "00011111", -- 2420 - 0x974  :   31 - 0x1f
    "00111111", -- 2421 - 0x975  :   63 - 0x3f
    "00111111", -- 2422 - 0x976  :   63 - 0x3f
    "00111111", -- 2423 - 0x977  :   63 - 0x3f
    "00110011", -- 2424 - 0x978  :   51 - 0x33 -- plane 1
    "00101111", -- 2425 - 0x979  :   47 - 0x2f
    "01101111", -- 2426 - 0x97a  :  111 - 0x6f
    "01011111", -- 2427 - 0x97b  :   95 - 0x5f
    "11011111", -- 2428 - 0x97c  :  223 - 0xdf
    "10111111", -- 2429 - 0x97d  :  191 - 0xbf
    "10111111", -- 2430 - 0x97e  :  191 - 0xbf
    "10111111", -- 2431 - 0x97f  :  191 - 0xbf
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Sprite 0x98
    "11111111", -- 2433 - 0x981  :  255 - 0xff
    "11111111", -- 2434 - 0x982  :  255 - 0xff
    "11111110", -- 2435 - 0x983  :  254 - 0xfe
    "11111001", -- 2436 - 0x984  :  249 - 0xf9
    "11100111", -- 2437 - 0x985  :  231 - 0xe7
    "11111100", -- 2438 - 0x986  :  252 - 0xfc
    "11110000", -- 2439 - 0x987  :  240 - 0xf0
    "11111111", -- 2440 - 0x988  :  255 - 0xff -- plane 1
    "11111111", -- 2441 - 0x989  :  255 - 0xff
    "11111111", -- 2442 - 0x98a  :  255 - 0xff
    "11111110", -- 2443 - 0x98b  :  254 - 0xfe
    "11111001", -- 2444 - 0x98c  :  249 - 0xf9
    "11100111", -- 2445 - 0x98d  :  231 - 0xe7
    "11111100", -- 2446 - 0x98e  :  252 - 0xfc
    "11110011", -- 2447 - 0x98f  :  243 - 0xf3
    "11110111", -- 2448 - 0x990  :  247 - 0xf7 -- Sprite 0x99
    "11111011", -- 2449 - 0x991  :  251 - 0xfb
    "11111011", -- 2450 - 0x992  :  251 - 0xfb
    "01110011", -- 2451 - 0x993  :  115 - 0x73
    "11000001", -- 2452 - 0x994  :  193 - 0xc1
    "00000011", -- 2453 - 0x995  :    3 - 0x3
    "00001111", -- 2454 - 0x996  :   15 - 0xf
    "00111111", -- 2455 - 0x997  :   63 - 0x3f
    "11110000", -- 2456 - 0x998  :  240 - 0xf0 -- plane 1
    "11111000", -- 2457 - 0x999  :  248 - 0xf8
    "11111000", -- 2458 - 0x99a  :  248 - 0xf8
    "01110000", -- 2459 - 0x99b  :  112 - 0x70
    "11001100", -- 2460 - 0x99c  :  204 - 0xcc
    "00110000", -- 2461 - 0x99d  :   48 - 0x30
    "11000000", -- 2462 - 0x99e  :  192 - 0xc0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "11111111", -- 2464 - 0x9a0  :  255 - 0xff -- Sprite 0x9a
    "11111111", -- 2465 - 0x9a1  :  255 - 0xff
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "10000000", -- 2467 - 0x9a3  :  128 - 0x80
    "10000000", -- 2468 - 0x9a4  :  128 - 0x80
    "10000000", -- 2469 - 0x9a5  :  128 - 0x80
    "10001111", -- 2470 - 0x9a6  :  143 - 0x8f
    "10001111", -- 2471 - 0x9a7  :  143 - 0x8f
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00111111", -- 2476 - 0x9ac  :   63 - 0x3f
    "00100000", -- 2477 - 0x9ad  :   32 - 0x20
    "00101111", -- 2478 - 0x9ae  :   47 - 0x2f
    "00101111", -- 2479 - 0x9af  :   47 - 0x2f
    "11111111", -- 2480 - 0x9b0  :  255 - 0xff -- Sprite 0x9b
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "11111111", -- 2482 - 0x9b2  :  255 - 0xff
    "00001111", -- 2483 - 0x9b3  :   15 - 0xf
    "00001111", -- 2484 - 0x9b4  :   15 - 0xf
    "00000111", -- 2485 - 0x9b5  :    7 - 0x7
    "11110111", -- 2486 - 0x9b6  :  247 - 0xf7
    "11110001", -- 2487 - 0x9b7  :  241 - 0xf1
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0 -- plane 1
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "11100000", -- 2492 - 0x9bc  :  224 - 0xe0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "11110000", -- 2494 - 0x9be  :  240 - 0xf0
    "11110000", -- 2495 - 0x9bf  :  240 - 0xf0
    "00011100", -- 2496 - 0x9c0  :   28 - 0x1c -- Sprite 0x9c
    "00011110", -- 2497 - 0x9c1  :   30 - 0x1e
    "00011111", -- 2498 - 0x9c2  :   31 - 0x1f
    "00011111", -- 2499 - 0x9c3  :   31 - 0x1f
    "00011111", -- 2500 - 0x9c4  :   31 - 0x1f
    "00011111", -- 2501 - 0x9c5  :   31 - 0x1f
    "00011111", -- 2502 - 0x9c6  :   31 - 0x1f
    "00011111", -- 2503 - 0x9c7  :   31 - 0x1f
    "01011101", -- 2504 - 0x9c8  :   93 - 0x5d -- plane 1
    "01011110", -- 2505 - 0x9c9  :   94 - 0x5e
    "01011111", -- 2506 - 0x9ca  :   95 - 0x5f
    "01011111", -- 2507 - 0x9cb  :   95 - 0x5f
    "01011111", -- 2508 - 0x9cc  :   95 - 0x5f
    "01011111", -- 2509 - 0x9cd  :   95 - 0x5f
    "01011111", -- 2510 - 0x9ce  :   95 - 0x5f
    "01011111", -- 2511 - 0x9cf  :   95 - 0x5f
    "00111110", -- 2512 - 0x9d0  :   62 - 0x3e -- Sprite 0x9d
    "00011100", -- 2513 - 0x9d1  :   28 - 0x1c
    "00001000", -- 2514 - 0x9d2  :    8 - 0x8
    "10000000", -- 2515 - 0x9d3  :  128 - 0x80
    "11000001", -- 2516 - 0x9d4  :  193 - 0xc1
    "11100011", -- 2517 - 0x9d5  :  227 - 0xe3
    "11110111", -- 2518 - 0x9d6  :  247 - 0xf7
    "11111111", -- 2519 - 0x9d7  :  255 - 0xff
    "10000000", -- 2520 - 0x9d8  :  128 - 0x80 -- plane 1
    "11000001", -- 2521 - 0x9d9  :  193 - 0xc1
    "01100011", -- 2522 - 0x9da  :   99 - 0x63
    "10110110", -- 2523 - 0x9db  :  182 - 0xb6
    "11011001", -- 2524 - 0x9dc  :  217 - 0xd9
    "11101011", -- 2525 - 0x9dd  :  235 - 0xeb
    "11110111", -- 2526 - 0x9de  :  247 - 0xf7
    "11111111", -- 2527 - 0x9df  :  255 - 0xff
    "00011100", -- 2528 - 0x9e0  :   28 - 0x1c -- Sprite 0x9e
    "00111100", -- 2529 - 0x9e1  :   60 - 0x3c
    "01111100", -- 2530 - 0x9e2  :  124 - 0x7c
    "11111100", -- 2531 - 0x9e3  :  252 - 0xfc
    "11111100", -- 2532 - 0x9e4  :  252 - 0xfc
    "11111100", -- 2533 - 0x9e5  :  252 - 0xfc
    "11111100", -- 2534 - 0x9e6  :  252 - 0xfc
    "11111100", -- 2535 - 0x9e7  :  252 - 0xfc
    "11011101", -- 2536 - 0x9e8  :  221 - 0xdd -- plane 1
    "10111101", -- 2537 - 0x9e9  :  189 - 0xbd
    "01111101", -- 2538 - 0x9ea  :  125 - 0x7d
    "11111101", -- 2539 - 0x9eb  :  253 - 0xfd
    "11111101", -- 2540 - 0x9ec  :  253 - 0xfd
    "11111101", -- 2541 - 0x9ed  :  253 - 0xfd
    "11111101", -- 2542 - 0x9ee  :  253 - 0xfd
    "11111101", -- 2543 - 0x9ef  :  253 - 0xfd
    "01111100", -- 2544 - 0x9f0  :  124 - 0x7c -- Sprite 0x9f
    "01111100", -- 2545 - 0x9f1  :  124 - 0x7c
    "01111000", -- 2546 - 0x9f2  :  120 - 0x78
    "01111000", -- 2547 - 0x9f3  :  120 - 0x78
    "01110001", -- 2548 - 0x9f4  :  113 - 0x71
    "01110001", -- 2549 - 0x9f5  :  113 - 0x71
    "01100011", -- 2550 - 0x9f6  :   99 - 0x63
    "01100011", -- 2551 - 0x9f7  :   99 - 0x63
    "00000001", -- 2552 - 0x9f8  :    1 - 0x1 -- plane 1
    "00000001", -- 2553 - 0x9f9  :    1 - 0x1
    "00000010", -- 2554 - 0x9fa  :    2 - 0x2
    "00000010", -- 2555 - 0x9fb  :    2 - 0x2
    "00000101", -- 2556 - 0x9fc  :    5 - 0x5
    "00000101", -- 2557 - 0x9fd  :    5 - 0x5
    "00001011", -- 2558 - 0x9fe  :   11 - 0xb
    "00001011", -- 2559 - 0x9ff  :   11 - 0xb
    "01110001", -- 2560 - 0xa00  :  113 - 0x71 -- Sprite 0xa0
    "01110000", -- 2561 - 0xa01  :  112 - 0x70
    "11111000", -- 2562 - 0xa02  :  248 - 0xf8
    "11111000", -- 2563 - 0xa03  :  248 - 0xf8
    "11111100", -- 2564 - 0xa04  :  252 - 0xfc
    "11111100", -- 2565 - 0xa05  :  252 - 0xfc
    "11111110", -- 2566 - 0xa06  :  254 - 0xfe
    "11111110", -- 2567 - 0xa07  :  254 - 0xfe
    "01110100", -- 2568 - 0xa08  :  116 - 0x74 -- plane 1
    "01110110", -- 2569 - 0xa09  :  118 - 0x76
    "11111010", -- 2570 - 0xa0a  :  250 - 0xfa
    "11111011", -- 2571 - 0xa0b  :  251 - 0xfb
    "11111101", -- 2572 - 0xa0c  :  253 - 0xfd
    "11111101", -- 2573 - 0xa0d  :  253 - 0xfd
    "11111110", -- 2574 - 0xa0e  :  254 - 0xfe
    "11111110", -- 2575 - 0xa0f  :  254 - 0xfe
    "11111000", -- 2576 - 0xa10  :  248 - 0xf8 -- Sprite 0xa1
    "11111000", -- 2577 - 0xa11  :  248 - 0xf8
    "11111000", -- 2578 - 0xa12  :  248 - 0xf8
    "01111000", -- 2579 - 0xa13  :  120 - 0x78
    "01111000", -- 2580 - 0xa14  :  120 - 0x78
    "00111000", -- 2581 - 0xa15  :   56 - 0x38
    "00111000", -- 2582 - 0xa16  :   56 - 0x38
    "00011000", -- 2583 - 0xa17  :   24 - 0x18
    "00000010", -- 2584 - 0xa18  :    2 - 0x2 -- plane 1
    "00000010", -- 2585 - 0xa19  :    2 - 0x2
    "00000010", -- 2586 - 0xa1a  :    2 - 0x2
    "00000010", -- 2587 - 0xa1b  :    2 - 0x2
    "00000010", -- 2588 - 0xa1c  :    2 - 0x2
    "10000010", -- 2589 - 0xa1d  :  130 - 0x82
    "10000010", -- 2590 - 0xa1e  :  130 - 0x82
    "11000010", -- 2591 - 0xa1f  :  194 - 0xc2
    "11100000", -- 2592 - 0xa20  :  224 - 0xe0 -- Sprite 0xa2
    "11110000", -- 2593 - 0xa21  :  240 - 0xf0
    "11111000", -- 2594 - 0xa22  :  248 - 0xf8
    "11111000", -- 2595 - 0xa23  :  248 - 0xf8
    "11111100", -- 2596 - 0xa24  :  252 - 0xfc
    "11111100", -- 2597 - 0xa25  :  252 - 0xfc
    "11111110", -- 2598 - 0xa26  :  254 - 0xfe
    "11111111", -- 2599 - 0xa27  :  255 - 0xff
    "11101010", -- 2600 - 0xa28  :  234 - 0xea -- plane 1
    "11110110", -- 2601 - 0xa29  :  246 - 0xf6
    "11111010", -- 2602 - 0xa2a  :  250 - 0xfa
    "11111010", -- 2603 - 0xa2b  :  250 - 0xfa
    "11111100", -- 2604 - 0xa2c  :  252 - 0xfc
    "11111100", -- 2605 - 0xa2d  :  252 - 0xfc
    "11111110", -- 2606 - 0xa2e  :  254 - 0xfe
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "11111111", -- 2608 - 0xa30  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 2609 - 0xa31  :  255 - 0xff
    "11111111", -- 2610 - 0xa32  :  255 - 0xff
    "11111111", -- 2611 - 0xa33  :  255 - 0xff
    "11111111", -- 2612 - 0xa34  :  255 - 0xff
    "11111111", -- 2613 - 0xa35  :  255 - 0xff
    "11111111", -- 2614 - 0xa36  :  255 - 0xff
    "11111111", -- 2615 - 0xa37  :  255 - 0xff
    "11111111", -- 2616 - 0xa38  :  255 - 0xff -- plane 1
    "11111111", -- 2617 - 0xa39  :  255 - 0xff
    "11111111", -- 2618 - 0xa3a  :  255 - 0xff
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "00011111", -- 2624 - 0xa40  :   31 - 0x1f -- Sprite 0xa4
    "00011111", -- 2625 - 0xa41  :   31 - 0x1f
    "00011111", -- 2626 - 0xa42  :   31 - 0x1f
    "00011111", -- 2627 - 0xa43  :   31 - 0x1f
    "00011111", -- 2628 - 0xa44  :   31 - 0x1f
    "00011111", -- 2629 - 0xa45  :   31 - 0x1f
    "00011111", -- 2630 - 0xa46  :   31 - 0x1f
    "00011111", -- 2631 - 0xa47  :   31 - 0x1f
    "01000000", -- 2632 - 0xa48  :   64 - 0x40 -- plane 1
    "01000000", -- 2633 - 0xa49  :   64 - 0x40
    "01000000", -- 2634 - 0xa4a  :   64 - 0x40
    "01000000", -- 2635 - 0xa4b  :   64 - 0x40
    "01000000", -- 2636 - 0xa4c  :   64 - 0x40
    "01000000", -- 2637 - 0xa4d  :   64 - 0x40
    "01000000", -- 2638 - 0xa4e  :   64 - 0x40
    "01000000", -- 2639 - 0xa4f  :   64 - 0x40
    "11111000", -- 2640 - 0xa50  :  248 - 0xf8 -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "11111000", -- 2643 - 0xa53  :  248 - 0xf8
    "11111000", -- 2644 - 0xa54  :  248 - 0xf8
    "11111000", -- 2645 - 0xa55  :  248 - 0xf8
    "11111000", -- 2646 - 0xa56  :  248 - 0xf8
    "11111000", -- 2647 - 0xa57  :  248 - 0xf8
    "11111000", -- 2648 - 0xa58  :  248 - 0xf8 -- plane 1
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111000", -- 2651 - 0xa5b  :  248 - 0xf8
    "11111011", -- 2652 - 0xa5c  :  251 - 0xfb
    "11111010", -- 2653 - 0xa5d  :  250 - 0xfa
    "11111010", -- 2654 - 0xa5e  :  250 - 0xfa
    "11111010", -- 2655 - 0xa5f  :  250 - 0xfa
    "11111100", -- 2656 - 0xa60  :  252 - 0xfc -- Sprite 0xa6
    "11111000", -- 2657 - 0xa61  :  248 - 0xf8
    "11110000", -- 2658 - 0xa62  :  240 - 0xf0
    "00000001", -- 2659 - 0xa63  :    1 - 0x1
    "00000001", -- 2660 - 0xa64  :    1 - 0x1
    "00000011", -- 2661 - 0xa65  :    3 - 0x3
    "11000011", -- 2662 - 0xa66  :  195 - 0xc3
    "10000111", -- 2663 - 0xa67  :  135 - 0x87
    "11111100", -- 2664 - 0xa68  :  252 - 0xfc -- plane 1
    "11111010", -- 2665 - 0xa69  :  250 - 0xfa
    "11110110", -- 2666 - 0xa6a  :  246 - 0xf6
    "00001101", -- 2667 - 0xa6b  :   13 - 0xd
    "11111001", -- 2668 - 0xa6c  :  249 - 0xf9
    "00000011", -- 2669 - 0xa6d  :    3 - 0x3
    "00010011", -- 2670 - 0xa6e  :   19 - 0x13
    "00110111", -- 2671 - 0xa6f  :   55 - 0x37
    "01111111", -- 2672 - 0xa70  :  127 - 0x7f -- Sprite 0xa7
    "11111001", -- 2673 - 0xa71  :  249 - 0xf9
    "11111001", -- 2674 - 0xa72  :  249 - 0xf9
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111110", -- 2676 - 0xa74  :  254 - 0xfe
    "11111100", -- 2677 - 0xa75  :  252 - 0xfc
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "01111111", -- 2680 - 0xa78  :  127 - 0x7f -- plane 1
    "11111001", -- 2681 - 0xa79  :  249 - 0xf9
    "11111001", -- 2682 - 0xa7a  :  249 - 0xf9
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111110", -- 2684 - 0xa7c  :  254 - 0xfe
    "11111100", -- 2685 - 0xa7d  :  252 - 0xfc
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "11110000", -- 2688 - 0xa80  :  240 - 0xf0 -- Sprite 0xa8
    "11110000", -- 2689 - 0xa81  :  240 - 0xf0
    "11111000", -- 2690 - 0xa82  :  248 - 0xf8
    "01111000", -- 2691 - 0xa83  :  120 - 0x78
    "11111100", -- 2692 - 0xa84  :  252 - 0xfc
    "11110100", -- 2693 - 0xa85  :  244 - 0xf4
    "11110110", -- 2694 - 0xa86  :  246 - 0xf6
    "11111010", -- 2695 - 0xa87  :  250 - 0xfa
    "11110110", -- 2696 - 0xa88  :  246 - 0xf6 -- plane 1
    "11110110", -- 2697 - 0xa89  :  246 - 0xf6
    "11111011", -- 2698 - 0xa8a  :  251 - 0xfb
    "01111011", -- 2699 - 0xa8b  :  123 - 0x7b
    "11111101", -- 2700 - 0xa8c  :  253 - 0xfd
    "11110101", -- 2701 - 0xa8d  :  245 - 0xf5
    "11110110", -- 2702 - 0xa8e  :  246 - 0xf6
    "11111010", -- 2703 - 0xa8f  :  250 - 0xfa
    "00111111", -- 2704 - 0xa90  :   63 - 0x3f -- Sprite 0xa9
    "00111111", -- 2705 - 0xa91  :   63 - 0x3f
    "00111111", -- 2706 - 0xa92  :   63 - 0x3f
    "00111111", -- 2707 - 0xa93  :   63 - 0x3f
    "00111111", -- 2708 - 0xa94  :   63 - 0x3f
    "00011111", -- 2709 - 0xa95  :   31 - 0x1f
    "00001111", -- 2710 - 0xa96  :   15 - 0xf
    "00000111", -- 2711 - 0xa97  :    7 - 0x7
    "10111111", -- 2712 - 0xa98  :  191 - 0xbf -- plane 1
    "10111111", -- 2713 - 0xa99  :  191 - 0xbf
    "00111111", -- 2714 - 0xa9a  :   63 - 0x3f
    "00111111", -- 2715 - 0xa9b  :   63 - 0x3f
    "10111111", -- 2716 - 0xa9c  :  191 - 0xbf
    "10011111", -- 2717 - 0xa9d  :  159 - 0x9f
    "11001111", -- 2718 - 0xa9e  :  207 - 0xcf
    "11010111", -- 2719 - 0xa9f  :  215 - 0xd7
    "11100000", -- 2720 - 0xaa0  :  224 - 0xe0 -- Sprite 0xaa
    "11111000", -- 2721 - 0xaa1  :  248 - 0xf8
    "11111111", -- 2722 - 0xaa2  :  255 - 0xff
    "11110011", -- 2723 - 0xaa3  :  243 - 0xf3
    "11111100", -- 2724 - 0xaa4  :  252 - 0xfc
    "11111111", -- 2725 - 0xaa5  :  255 - 0xff
    "11111111", -- 2726 - 0xaa6  :  255 - 0xff
    "11111111", -- 2727 - 0xaa7  :  255 - 0xff
    "11100100", -- 2728 - 0xaa8  :  228 - 0xe4 -- plane 1
    "11111000", -- 2729 - 0xaa9  :  248 - 0xf8
    "11111111", -- 2730 - 0xaaa  :  255 - 0xff
    "11110011", -- 2731 - 0xaab  :  243 - 0xf3
    "11111100", -- 2732 - 0xaac  :  252 - 0xfc
    "11111111", -- 2733 - 0xaad  :  255 - 0xff
    "11111111", -- 2734 - 0xaae  :  255 - 0xff
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "11111111", -- 2736 - 0xab0  :  255 - 0xff -- Sprite 0xab
    "11111111", -- 2737 - 0xab1  :  255 - 0xff
    "00111111", -- 2738 - 0xab2  :   63 - 0x3f
    "11001111", -- 2739 - 0xab3  :  207 - 0xcf
    "11110011", -- 2740 - 0xab4  :  243 - 0xf3
    "00111101", -- 2741 - 0xab5  :   61 - 0x3d
    "11011000", -- 2742 - 0xab6  :  216 - 0xd8
    "10110000", -- 2743 - 0xab7  :  176 - 0xb0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- plane 1
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "11000000", -- 2747 - 0xabb  :  192 - 0xc0
    "11110000", -- 2748 - 0xabc  :  240 - 0xf0
    "00111100", -- 2749 - 0xabd  :   60 - 0x3c
    "11011000", -- 2750 - 0xabe  :  216 - 0xd8
    "10110110", -- 2751 - 0xabf  :  182 - 0xb6
    "10001111", -- 2752 - 0xac0  :  143 - 0x8f -- Sprite 0xac
    "11101111", -- 2753 - 0xac1  :  239 - 0xef
    "11100000", -- 2754 - 0xac2  :  224 - 0xe0
    "11111000", -- 2755 - 0xac3  :  248 - 0xf8
    "11111000", -- 2756 - 0xac4  :  248 - 0xf8
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "11111111", -- 2758 - 0xac6  :  255 - 0xff
    "11111111", -- 2759 - 0xac7  :  255 - 0xff
    "00001111", -- 2760 - 0xac8  :   15 - 0xf -- plane 1
    "00001111", -- 2761 - 0xac9  :   15 - 0xf
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000011", -- 2763 - 0xacb  :    3 - 0x3
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "11110001", -- 2768 - 0xad0  :  241 - 0xf1 -- Sprite 0xad
    "11110001", -- 2769 - 0xad1  :  241 - 0xf1
    "00000001", -- 2770 - 0xad2  :    1 - 0x1
    "00000001", -- 2771 - 0xad3  :    1 - 0x1
    "00000001", -- 2772 - 0xad4  :    1 - 0x1
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "11110100", -- 2776 - 0xad8  :  244 - 0xf4 -- plane 1
    "11110100", -- 2777 - 0xad9  :  244 - 0xf4
    "00000100", -- 2778 - 0xada  :    4 - 0x4
    "11111100", -- 2779 - 0xadb  :  252 - 0xfc
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00011111", -- 2784 - 0xae0  :   31 - 0x1f -- Sprite 0xae
    "00011111", -- 2785 - 0xae1  :   31 - 0x1f
    "00011111", -- 2786 - 0xae2  :   31 - 0x1f
    "00011111", -- 2787 - 0xae3  :   31 - 0x1f
    "00011111", -- 2788 - 0xae4  :   31 - 0x1f
    "00011111", -- 2789 - 0xae5  :   31 - 0x1f
    "00011111", -- 2790 - 0xae6  :   31 - 0x1f
    "00011111", -- 2791 - 0xae7  :   31 - 0x1f
    "01011111", -- 2792 - 0xae8  :   95 - 0x5f -- plane 1
    "01011111", -- 2793 - 0xae9  :   95 - 0x5f
    "01011111", -- 2794 - 0xaea  :   95 - 0x5f
    "01011111", -- 2795 - 0xaeb  :   95 - 0x5f
    "01011111", -- 2796 - 0xaec  :   95 - 0x5f
    "01011111", -- 2797 - 0xaed  :   95 - 0x5f
    "01011111", -- 2798 - 0xaee  :   95 - 0x5f
    "01011111", -- 2799 - 0xaef  :   95 - 0x5f
    "11111100", -- 2800 - 0xaf0  :  252 - 0xfc -- Sprite 0xaf
    "11111100", -- 2801 - 0xaf1  :  252 - 0xfc
    "11111100", -- 2802 - 0xaf2  :  252 - 0xfc
    "11111100", -- 2803 - 0xaf3  :  252 - 0xfc
    "11110100", -- 2804 - 0xaf4  :  244 - 0xf4
    "11110100", -- 2805 - 0xaf5  :  244 - 0xf4
    "11110100", -- 2806 - 0xaf6  :  244 - 0xf4
    "11110100", -- 2807 - 0xaf7  :  244 - 0xf4
    "11111101", -- 2808 - 0xaf8  :  253 - 0xfd -- plane 1
    "11111101", -- 2809 - 0xaf9  :  253 - 0xfd
    "11111101", -- 2810 - 0xafa  :  253 - 0xfd
    "11111101", -- 2811 - 0xafb  :  253 - 0xfd
    "11110101", -- 2812 - 0xafc  :  245 - 0xf5
    "11110101", -- 2813 - 0xafd  :  245 - 0xf5
    "11110101", -- 2814 - 0xafe  :  245 - 0xf5
    "11110101", -- 2815 - 0xaff  :  245 - 0xf5
    "00001100", -- 2816 - 0xb00  :   12 - 0xc -- Sprite 0xb0
    "00011100", -- 2817 - 0xb01  :   28 - 0x1c
    "00001100", -- 2818 - 0xb02  :   12 - 0xc
    "00001100", -- 2819 - 0xb03  :   12 - 0xc
    "00001100", -- 2820 - 0xb04  :   12 - 0xc
    "00001100", -- 2821 - 0xb05  :   12 - 0xc
    "00111111", -- 2822 - 0xb06  :   63 - 0x3f
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00001100", -- 2824 - 0xb08  :   12 - 0xc -- plane 1
    "00011100", -- 2825 - 0xb09  :   28 - 0x1c
    "00001100", -- 2826 - 0xb0a  :   12 - 0xc
    "00001100", -- 2827 - 0xb0b  :   12 - 0xc
    "00001100", -- 2828 - 0xb0c  :   12 - 0xc
    "00001100", -- 2829 - 0xb0d  :   12 - 0xc
    "00111111", -- 2830 - 0xb0e  :   63 - 0x3f
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00111110", -- 2832 - 0xb10  :   62 - 0x3e -- Sprite 0xb1
    "01100011", -- 2833 - 0xb11  :   99 - 0x63
    "00000111", -- 2834 - 0xb12  :    7 - 0x7
    "00011110", -- 2835 - 0xb13  :   30 - 0x1e
    "00111100", -- 2836 - 0xb14  :   60 - 0x3c
    "01110000", -- 2837 - 0xb15  :  112 - 0x70
    "01111111", -- 2838 - 0xb16  :  127 - 0x7f
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00111110", -- 2840 - 0xb18  :   62 - 0x3e -- plane 1
    "01100011", -- 2841 - 0xb19  :   99 - 0x63
    "00000111", -- 2842 - 0xb1a  :    7 - 0x7
    "00011110", -- 2843 - 0xb1b  :   30 - 0x1e
    "00111100", -- 2844 - 0xb1c  :   60 - 0x3c
    "01110000", -- 2845 - 0xb1d  :  112 - 0x70
    "01111111", -- 2846 - 0xb1e  :  127 - 0x7f
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "01111110", -- 2848 - 0xb20  :  126 - 0x7e -- Sprite 0xb2
    "01100011", -- 2849 - 0xb21  :   99 - 0x63
    "01100011", -- 2850 - 0xb22  :   99 - 0x63
    "01100011", -- 2851 - 0xb23  :   99 - 0x63
    "01111110", -- 2852 - 0xb24  :  126 - 0x7e
    "01100000", -- 2853 - 0xb25  :   96 - 0x60
    "01100000", -- 2854 - 0xb26  :   96 - 0x60
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "01111110", -- 2856 - 0xb28  :  126 - 0x7e -- plane 1
    "01100011", -- 2857 - 0xb29  :   99 - 0x63
    "01100011", -- 2858 - 0xb2a  :   99 - 0x63
    "01100011", -- 2859 - 0xb2b  :   99 - 0x63
    "01111110", -- 2860 - 0xb2c  :  126 - 0x7e
    "01100000", -- 2861 - 0xb2d  :   96 - 0x60
    "01100000", -- 2862 - 0xb2e  :   96 - 0x60
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "01100011", -- 2864 - 0xb30  :   99 - 0x63 -- Sprite 0xb3
    "01100011", -- 2865 - 0xb31  :   99 - 0x63
    "01100011", -- 2866 - 0xb32  :   99 - 0x63
    "01100011", -- 2867 - 0xb33  :   99 - 0x63
    "01100011", -- 2868 - 0xb34  :   99 - 0x63
    "01100011", -- 2869 - 0xb35  :   99 - 0x63
    "00111110", -- 2870 - 0xb36  :   62 - 0x3e
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "01100011", -- 2872 - 0xb38  :   99 - 0x63 -- plane 1
    "01100011", -- 2873 - 0xb39  :   99 - 0x63
    "01100011", -- 2874 - 0xb3a  :   99 - 0x63
    "01100011", -- 2875 - 0xb3b  :   99 - 0x63
    "01100011", -- 2876 - 0xb3c  :   99 - 0x63
    "01100011", -- 2877 - 0xb3d  :   99 - 0x63
    "00111110", -- 2878 - 0xb3e  :   62 - 0x3e
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "01100011", -- 2880 - 0xb40  :   99 - 0x63 -- Sprite 0xb4
    "01100011", -- 2881 - 0xb41  :   99 - 0x63
    "01100011", -- 2882 - 0xb42  :   99 - 0x63
    "01111111", -- 2883 - 0xb43  :  127 - 0x7f
    "01100011", -- 2884 - 0xb44  :   99 - 0x63
    "01100011", -- 2885 - 0xb45  :   99 - 0x63
    "01100011", -- 2886 - 0xb46  :   99 - 0x63
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "01100011", -- 2888 - 0xb48  :   99 - 0x63 -- plane 1
    "01100011", -- 2889 - 0xb49  :   99 - 0x63
    "01100011", -- 2890 - 0xb4a  :   99 - 0x63
    "01111111", -- 2891 - 0xb4b  :  127 - 0x7f
    "01100011", -- 2892 - 0xb4c  :   99 - 0x63
    "01100011", -- 2893 - 0xb4d  :   99 - 0x63
    "01100011", -- 2894 - 0xb4e  :   99 - 0x63
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00111111", -- 2896 - 0xb50  :   63 - 0x3f -- Sprite 0xb5
    "00001100", -- 2897 - 0xb51  :   12 - 0xc
    "00001100", -- 2898 - 0xb52  :   12 - 0xc
    "00001100", -- 2899 - 0xb53  :   12 - 0xc
    "00001100", -- 2900 - 0xb54  :   12 - 0xc
    "00001100", -- 2901 - 0xb55  :   12 - 0xc
    "00111111", -- 2902 - 0xb56  :   63 - 0x3f
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00111111", -- 2904 - 0xb58  :   63 - 0x3f -- plane 1
    "00001100", -- 2905 - 0xb59  :   12 - 0xc
    "00001100", -- 2906 - 0xb5a  :   12 - 0xc
    "00001100", -- 2907 - 0xb5b  :   12 - 0xc
    "00001100", -- 2908 - 0xb5c  :   12 - 0xc
    "00001100", -- 2909 - 0xb5d  :   12 - 0xc
    "00111111", -- 2910 - 0xb5e  :   63 - 0x3f
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Sprite 0xb6
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "01111110", -- 2915 - 0xb63  :  126 - 0x7e
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- plane 1
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "01111110", -- 2923 - 0xb6b  :  126 - 0x7e
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00111100", -- 2928 - 0xb70  :   60 - 0x3c -- Sprite 0xb7
    "01100110", -- 2929 - 0xb71  :  102 - 0x66
    "01100000", -- 2930 - 0xb72  :   96 - 0x60
    "00111110", -- 2931 - 0xb73  :   62 - 0x3e
    "00000011", -- 2932 - 0xb74  :    3 - 0x3
    "01100011", -- 2933 - 0xb75  :   99 - 0x63
    "00111110", -- 2934 - 0xb76  :   62 - 0x3e
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00111100", -- 2936 - 0xb78  :   60 - 0x3c -- plane 1
    "01100110", -- 2937 - 0xb79  :  102 - 0x66
    "01100000", -- 2938 - 0xb7a  :   96 - 0x60
    "00111110", -- 2939 - 0xb7b  :   62 - 0x3e
    "00000011", -- 2940 - 0xb7c  :    3 - 0x3
    "01100011", -- 2941 - 0xb7d  :   99 - 0x63
    "00111110", -- 2942 - 0xb7e  :   62 - 0x3e
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00011110", -- 2944 - 0xb80  :   30 - 0x1e -- Sprite 0xb8
    "00110011", -- 2945 - 0xb81  :   51 - 0x33
    "01100000", -- 2946 - 0xb82  :   96 - 0x60
    "01100000", -- 2947 - 0xb83  :   96 - 0x60
    "01100000", -- 2948 - 0xb84  :   96 - 0x60
    "00110011", -- 2949 - 0xb85  :   51 - 0x33
    "00011110", -- 2950 - 0xb86  :   30 - 0x1e
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00011110", -- 2952 - 0xb88  :   30 - 0x1e -- plane 1
    "00110011", -- 2953 - 0xb89  :   51 - 0x33
    "01100000", -- 2954 - 0xb8a  :   96 - 0x60
    "01100000", -- 2955 - 0xb8b  :   96 - 0x60
    "01100000", -- 2956 - 0xb8c  :   96 - 0x60
    "00110011", -- 2957 - 0xb8d  :   51 - 0x33
    "00011110", -- 2958 - 0xb8e  :   30 - 0x1e
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00111110", -- 2960 - 0xb90  :   62 - 0x3e -- Sprite 0xb9
    "01100011", -- 2961 - 0xb91  :   99 - 0x63
    "01100011", -- 2962 - 0xb92  :   99 - 0x63
    "01100011", -- 2963 - 0xb93  :   99 - 0x63
    "01100011", -- 2964 - 0xb94  :   99 - 0x63
    "01100011", -- 2965 - 0xb95  :   99 - 0x63
    "00111110", -- 2966 - 0xb96  :   62 - 0x3e
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00111110", -- 2968 - 0xb98  :   62 - 0x3e -- plane 1
    "01100011", -- 2969 - 0xb99  :   99 - 0x63
    "01100011", -- 2970 - 0xb9a  :   99 - 0x63
    "01100011", -- 2971 - 0xb9b  :   99 - 0x63
    "01100011", -- 2972 - 0xb9c  :   99 - 0x63
    "01100011", -- 2973 - 0xb9d  :   99 - 0x63
    "00111110", -- 2974 - 0xb9e  :   62 - 0x3e
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "01111110", -- 2976 - 0xba0  :  126 - 0x7e -- Sprite 0xba
    "01100011", -- 2977 - 0xba1  :   99 - 0x63
    "01100011", -- 2978 - 0xba2  :   99 - 0x63
    "01100111", -- 2979 - 0xba3  :  103 - 0x67
    "01111100", -- 2980 - 0xba4  :  124 - 0x7c
    "01101110", -- 2981 - 0xba5  :  110 - 0x6e
    "01100111", -- 2982 - 0xba6  :  103 - 0x67
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "01111110", -- 2984 - 0xba8  :  126 - 0x7e -- plane 1
    "01100011", -- 2985 - 0xba9  :   99 - 0x63
    "01100011", -- 2986 - 0xbaa  :   99 - 0x63
    "01100111", -- 2987 - 0xbab  :  103 - 0x67
    "01111100", -- 2988 - 0xbac  :  124 - 0x7c
    "01101110", -- 2989 - 0xbad  :  110 - 0x6e
    "01100111", -- 2990 - 0xbae  :  103 - 0x67
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "01111111", -- 2992 - 0xbb0  :  127 - 0x7f -- Sprite 0xbb
    "01100000", -- 2993 - 0xbb1  :   96 - 0x60
    "01100000", -- 2994 - 0xbb2  :   96 - 0x60
    "01111110", -- 2995 - 0xbb3  :  126 - 0x7e
    "01100000", -- 2996 - 0xbb4  :   96 - 0x60
    "01100000", -- 2997 - 0xbb5  :   96 - 0x60
    "01111111", -- 2998 - 0xbb6  :  127 - 0x7f
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "01111111", -- 3000 - 0xbb8  :  127 - 0x7f -- plane 1
    "01100000", -- 3001 - 0xbb9  :   96 - 0x60
    "01100000", -- 3002 - 0xbba  :   96 - 0x60
    "01111110", -- 3003 - 0xbbb  :  126 - 0x7e
    "01100000", -- 3004 - 0xbbc  :   96 - 0x60
    "01100000", -- 3005 - 0xbbd  :   96 - 0x60
    "01111111", -- 3006 - 0xbbe  :  127 - 0x7f
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Sprite 0xbc
    "00100010", -- 3009 - 0xbc1  :   34 - 0x22
    "01100101", -- 3010 - 0xbc2  :  101 - 0x65
    "00100101", -- 3011 - 0xbc3  :   37 - 0x25
    "00100101", -- 3012 - 0xbc4  :   37 - 0x25
    "01110010", -- 3013 - 0xbc5  :  114 - 0x72
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Sprite 0xbd
    "01110010", -- 3025 - 0xbd1  :  114 - 0x72
    "01000101", -- 3026 - 0xbd2  :   69 - 0x45
    "01100101", -- 3027 - 0xbd3  :  101 - 0x65
    "00010101", -- 3028 - 0xbd4  :   21 - 0x15
    "01100010", -- 3029 - 0xbd5  :   98 - 0x62
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Sprite 0xbe
    "01100111", -- 3041 - 0xbe1  :  103 - 0x67
    "01010010", -- 3042 - 0xbe2  :   82 - 0x52
    "01100010", -- 3043 - 0xbe3  :   98 - 0x62
    "01000010", -- 3044 - 0xbe4  :   66 - 0x42
    "01000010", -- 3045 - 0xbe5  :   66 - 0x42
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- plane 1
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "01100000", -- 3057 - 0xbf1  :   96 - 0x60
    "10000000", -- 3058 - 0xbf2  :  128 - 0x80
    "01000000", -- 3059 - 0xbf3  :   64 - 0x40
    "00100000", -- 3060 - 0xbf4  :   32 - 0x20
    "11000110", -- 3061 - 0xbf5  :  198 - 0xc6
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "01100011", -- 3072 - 0xc00  :   99 - 0x63 -- Sprite 0xc0
    "01100110", -- 3073 - 0xc01  :  102 - 0x66
    "01101100", -- 3074 - 0xc02  :  108 - 0x6c
    "01111000", -- 3075 - 0xc03  :  120 - 0x78
    "01111100", -- 3076 - 0xc04  :  124 - 0x7c
    "01100110", -- 3077 - 0xc05  :  102 - 0x66
    "01100011", -- 3078 - 0xc06  :   99 - 0x63
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "01100011", -- 3080 - 0xc08  :   99 - 0x63 -- plane 1
    "01100110", -- 3081 - 0xc09  :  102 - 0x66
    "01101100", -- 3082 - 0xc0a  :  108 - 0x6c
    "01111000", -- 3083 - 0xc0b  :  120 - 0x78
    "01111100", -- 3084 - 0xc0c  :  124 - 0x7c
    "01100110", -- 3085 - 0xc0d  :  102 - 0x66
    "01100011", -- 3086 - 0xc0e  :   99 - 0x63
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00111111", -- 3088 - 0xc10  :   63 - 0x3f -- Sprite 0xc1
    "00001100", -- 3089 - 0xc11  :   12 - 0xc
    "00001100", -- 3090 - 0xc12  :   12 - 0xc
    "00001100", -- 3091 - 0xc13  :   12 - 0xc
    "00001100", -- 3092 - 0xc14  :   12 - 0xc
    "00001100", -- 3093 - 0xc15  :   12 - 0xc
    "00111111", -- 3094 - 0xc16  :   63 - 0x3f
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00111111", -- 3096 - 0xc18  :   63 - 0x3f -- plane 1
    "00001100", -- 3097 - 0xc19  :   12 - 0xc
    "00001100", -- 3098 - 0xc1a  :   12 - 0xc
    "00001100", -- 3099 - 0xc1b  :   12 - 0xc
    "00001100", -- 3100 - 0xc1c  :   12 - 0xc
    "00001100", -- 3101 - 0xc1d  :   12 - 0xc
    "00111111", -- 3102 - 0xc1e  :   63 - 0x3f
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "01100011", -- 3104 - 0xc20  :   99 - 0x63 -- Sprite 0xc2
    "01110111", -- 3105 - 0xc21  :  119 - 0x77
    "01111111", -- 3106 - 0xc22  :  127 - 0x7f
    "01111111", -- 3107 - 0xc23  :  127 - 0x7f
    "01101011", -- 3108 - 0xc24  :  107 - 0x6b
    "01100011", -- 3109 - 0xc25  :   99 - 0x63
    "01100011", -- 3110 - 0xc26  :   99 - 0x63
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "01100011", -- 3112 - 0xc28  :   99 - 0x63 -- plane 1
    "01110111", -- 3113 - 0xc29  :  119 - 0x77
    "01111111", -- 3114 - 0xc2a  :  127 - 0x7f
    "01111111", -- 3115 - 0xc2b  :  127 - 0x7f
    "01101011", -- 3116 - 0xc2c  :  107 - 0x6b
    "01100011", -- 3117 - 0xc2d  :   99 - 0x63
    "01100011", -- 3118 - 0xc2e  :   99 - 0x63
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00011100", -- 3120 - 0xc30  :   28 - 0x1c -- Sprite 0xc3
    "00110110", -- 3121 - 0xc31  :   54 - 0x36
    "01100011", -- 3122 - 0xc32  :   99 - 0x63
    "01100011", -- 3123 - 0xc33  :   99 - 0x63
    "01111111", -- 3124 - 0xc34  :  127 - 0x7f
    "01100011", -- 3125 - 0xc35  :   99 - 0x63
    "01100011", -- 3126 - 0xc36  :   99 - 0x63
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00011100", -- 3128 - 0xc38  :   28 - 0x1c -- plane 1
    "00110110", -- 3129 - 0xc39  :   54 - 0x36
    "01100011", -- 3130 - 0xc3a  :   99 - 0x63
    "01100011", -- 3131 - 0xc3b  :   99 - 0x63
    "01111111", -- 3132 - 0xc3c  :  127 - 0x7f
    "01100011", -- 3133 - 0xc3d  :   99 - 0x63
    "01100011", -- 3134 - 0xc3e  :   99 - 0x63
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00011111", -- 3136 - 0xc40  :   31 - 0x1f -- Sprite 0xc4
    "00110000", -- 3137 - 0xc41  :   48 - 0x30
    "01100000", -- 3138 - 0xc42  :   96 - 0x60
    "01100111", -- 3139 - 0xc43  :  103 - 0x67
    "01100011", -- 3140 - 0xc44  :   99 - 0x63
    "00110011", -- 3141 - 0xc45  :   51 - 0x33
    "00011111", -- 3142 - 0xc46  :   31 - 0x1f
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00011111", -- 3144 - 0xc48  :   31 - 0x1f -- plane 1
    "00110000", -- 3145 - 0xc49  :   48 - 0x30
    "01100000", -- 3146 - 0xc4a  :   96 - 0x60
    "01100111", -- 3147 - 0xc4b  :  103 - 0x67
    "01100011", -- 3148 - 0xc4c  :   99 - 0x63
    "00110011", -- 3149 - 0xc4d  :   51 - 0x33
    "00011111", -- 3150 - 0xc4e  :   31 - 0x1f
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "01100011", -- 3152 - 0xc50  :   99 - 0x63 -- Sprite 0xc5
    "01100011", -- 3153 - 0xc51  :   99 - 0x63
    "01100011", -- 3154 - 0xc52  :   99 - 0x63
    "01100011", -- 3155 - 0xc53  :   99 - 0x63
    "01100011", -- 3156 - 0xc54  :   99 - 0x63
    "01100011", -- 3157 - 0xc55  :   99 - 0x63
    "00111110", -- 3158 - 0xc56  :   62 - 0x3e
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "01100011", -- 3160 - 0xc58  :   99 - 0x63 -- plane 1
    "01100011", -- 3161 - 0xc59  :   99 - 0x63
    "01100011", -- 3162 - 0xc5a  :   99 - 0x63
    "01100011", -- 3163 - 0xc5b  :   99 - 0x63
    "01100011", -- 3164 - 0xc5c  :   99 - 0x63
    "01100011", -- 3165 - 0xc5d  :   99 - 0x63
    "00111110", -- 3166 - 0xc5e  :   62 - 0x3e
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "01111110", -- 3168 - 0xc60  :  126 - 0x7e -- Sprite 0xc6
    "01100011", -- 3169 - 0xc61  :   99 - 0x63
    "01100011", -- 3170 - 0xc62  :   99 - 0x63
    "01100111", -- 3171 - 0xc63  :  103 - 0x67
    "01111100", -- 3172 - 0xc64  :  124 - 0x7c
    "01101110", -- 3173 - 0xc65  :  110 - 0x6e
    "01100111", -- 3174 - 0xc66  :  103 - 0x67
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "01111110", -- 3176 - 0xc68  :  126 - 0x7e -- plane 1
    "01100011", -- 3177 - 0xc69  :   99 - 0x63
    "01100011", -- 3178 - 0xc6a  :   99 - 0x63
    "01100111", -- 3179 - 0xc6b  :  103 - 0x67
    "01111100", -- 3180 - 0xc6c  :  124 - 0x7c
    "01101110", -- 3181 - 0xc6d  :  110 - 0x6e
    "01100111", -- 3182 - 0xc6e  :  103 - 0x67
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "01111111", -- 3184 - 0xc70  :  127 - 0x7f -- Sprite 0xc7
    "01100000", -- 3185 - 0xc71  :   96 - 0x60
    "01100000", -- 3186 - 0xc72  :   96 - 0x60
    "01111110", -- 3187 - 0xc73  :  126 - 0x7e
    "01100000", -- 3188 - 0xc74  :   96 - 0x60
    "01100000", -- 3189 - 0xc75  :   96 - 0x60
    "01111111", -- 3190 - 0xc76  :  127 - 0x7f
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "01111111", -- 3192 - 0xc78  :  127 - 0x7f -- plane 1
    "01100000", -- 3193 - 0xc79  :   96 - 0x60
    "01100000", -- 3194 - 0xc7a  :   96 - 0x60
    "01111110", -- 3195 - 0xc7b  :  126 - 0x7e
    "01100000", -- 3196 - 0xc7c  :   96 - 0x60
    "01100000", -- 3197 - 0xc7d  :   96 - 0x60
    "01111111", -- 3198 - 0xc7e  :  127 - 0x7f
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00110110", -- 3200 - 0xc80  :   54 - 0x36 -- Sprite 0xc8
    "00110110", -- 3201 - 0xc81  :   54 - 0x36
    "00010010", -- 3202 - 0xc82  :   18 - 0x12
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00110110", -- 3208 - 0xc88  :   54 - 0x36 -- plane 1
    "00110110", -- 3209 - 0xc89  :   54 - 0x36
    "00010010", -- 3210 - 0xc8a  :   18 - 0x12
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00111110", -- 3216 - 0xc90  :   62 - 0x3e -- Sprite 0xc9
    "01100011", -- 3217 - 0xc91  :   99 - 0x63
    "01100011", -- 3218 - 0xc92  :   99 - 0x63
    "01100011", -- 3219 - 0xc93  :   99 - 0x63
    "01100011", -- 3220 - 0xc94  :   99 - 0x63
    "01100011", -- 3221 - 0xc95  :   99 - 0x63
    "00111110", -- 3222 - 0xc96  :   62 - 0x3e
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00111110", -- 3224 - 0xc98  :   62 - 0x3e -- plane 1
    "01100011", -- 3225 - 0xc99  :   99 - 0x63
    "01100011", -- 3226 - 0xc9a  :   99 - 0x63
    "01100011", -- 3227 - 0xc9b  :   99 - 0x63
    "01100011", -- 3228 - 0xc9c  :   99 - 0x63
    "01100011", -- 3229 - 0xc9d  :   99 - 0x63
    "00111110", -- 3230 - 0xc9e  :   62 - 0x3e
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00111100", -- 3232 - 0xca0  :   60 - 0x3c -- Sprite 0xca
    "01100110", -- 3233 - 0xca1  :  102 - 0x66
    "01100000", -- 3234 - 0xca2  :   96 - 0x60
    "00111110", -- 3235 - 0xca3  :   62 - 0x3e
    "00000011", -- 3236 - 0xca4  :    3 - 0x3
    "01100011", -- 3237 - 0xca5  :   99 - 0x63
    "00111110", -- 3238 - 0xca6  :   62 - 0x3e
    "00000000", -- 3239 - 0xca7  :    0 - 0x0
    "00111100", -- 3240 - 0xca8  :   60 - 0x3c -- plane 1
    "01100110", -- 3241 - 0xca9  :  102 - 0x66
    "01100000", -- 3242 - 0xcaa  :   96 - 0x60
    "00111110", -- 3243 - 0xcab  :   62 - 0x3e
    "00000011", -- 3244 - 0xcac  :    3 - 0x3
    "01100011", -- 3245 - 0xcad  :   99 - 0x63
    "00111110", -- 3246 - 0xcae  :   62 - 0x3e
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00000000", -- 3250 - 0xcb2  :    0 - 0x0
    "00000000", -- 3251 - 0xcb3  :    0 - 0x0
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0 -- plane 1
    "00111000", -- 3257 - 0xcb9  :   56 - 0x38
    "01111100", -- 3258 - 0xcba  :  124 - 0x7c
    "11111110", -- 3259 - 0xcbb  :  254 - 0xfe
    "11111110", -- 3260 - 0xcbc  :  254 - 0xfe
    "11111110", -- 3261 - 0xcbd  :  254 - 0xfe
    "01111100", -- 3262 - 0xcbe  :  124 - 0x7c
    "00111000", -- 3263 - 0xcbf  :   56 - 0x38
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000000", -- 3302 - 0xce6  :    0 - 0x0
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- plane 1
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000000", -- 3309 - 0xced  :    0 - 0x0
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "01000111", -- 3328 - 0xd00  :   71 - 0x47 -- Sprite 0xd0
    "01000111", -- 3329 - 0xd01  :   71 - 0x47
    "00001111", -- 3330 - 0xd02  :   15 - 0xf
    "00001111", -- 3331 - 0xd03  :   15 - 0xf
    "00011111", -- 3332 - 0xd04  :   31 - 0x1f
    "00011111", -- 3333 - 0xd05  :   31 - 0x1f
    "00111111", -- 3334 - 0xd06  :   63 - 0x3f
    "00111111", -- 3335 - 0xd07  :   63 - 0x3f
    "00010111", -- 3336 - 0xd08  :   23 - 0x17 -- plane 1
    "00010111", -- 3337 - 0xd09  :   23 - 0x17
    "00101111", -- 3338 - 0xd0a  :   47 - 0x2f
    "00101111", -- 3339 - 0xd0b  :   47 - 0x2f
    "01011111", -- 3340 - 0xd0c  :   95 - 0x5f
    "01011111", -- 3341 - 0xd0d  :   95 - 0x5f
    "00111111", -- 3342 - 0xd0e  :   63 - 0x3f
    "00111111", -- 3343 - 0xd0f  :   63 - 0x3f
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Sprite 0xd1
    "11001111", -- 3345 - 0xd11  :  207 - 0xcf
    "11001111", -- 3346 - 0xd12  :  207 - 0xcf
    "11111011", -- 3347 - 0xd13  :  251 - 0xfb
    "11110111", -- 3348 - 0xd14  :  247 - 0xf7
    "11100111", -- 3349 - 0xd15  :  231 - 0xe7
    "11111111", -- 3350 - 0xd16  :  255 - 0xff
    "11111111", -- 3351 - 0xd17  :  255 - 0xff
    "11111111", -- 3352 - 0xd18  :  255 - 0xff -- plane 1
    "11001111", -- 3353 - 0xd19  :  207 - 0xcf
    "11001111", -- 3354 - 0xd1a  :  207 - 0xcf
    "11111011", -- 3355 - 0xd1b  :  251 - 0xfb
    "11110111", -- 3356 - 0xd1c  :  247 - 0xf7
    "11100111", -- 3357 - 0xd1d  :  231 - 0xe7
    "11111111", -- 3358 - 0xd1e  :  255 - 0xff
    "11111111", -- 3359 - 0xd1f  :  255 - 0xff
    "00011000", -- 3360 - 0xd20  :   24 - 0x18 -- Sprite 0xd2
    "00001000", -- 3361 - 0xd21  :    8 - 0x8
    "10001000", -- 3362 - 0xd22  :  136 - 0x88
    "10000000", -- 3363 - 0xd23  :  128 - 0x80
    "01000000", -- 3364 - 0xd24  :   64 - 0x40
    "01000000", -- 3365 - 0xd25  :   64 - 0x40
    "10100000", -- 3366 - 0xd26  :  160 - 0xa0
    "10100000", -- 3367 - 0xd27  :  160 - 0xa0
    "01000010", -- 3368 - 0xd28  :   66 - 0x42 -- plane 1
    "01100010", -- 3369 - 0xd29  :   98 - 0x62
    "10100010", -- 3370 - 0xd2a  :  162 - 0xa2
    "10110010", -- 3371 - 0xd2b  :  178 - 0xb2
    "01010010", -- 3372 - 0xd2c  :   82 - 0x52
    "01011010", -- 3373 - 0xd2d  :   90 - 0x5a
    "10101010", -- 3374 - 0xd2e  :  170 - 0xaa
    "10101100", -- 3375 - 0xd2f  :  172 - 0xac
    "11111111", -- 3376 - 0xd30  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11111101", -- 3380 - 0xd34  :  253 - 0xfd
    "11111101", -- 3381 - 0xd35  :  253 - 0xfd
    "11111101", -- 3382 - 0xd36  :  253 - 0xfd
    "11111101", -- 3383 - 0xd37  :  253 - 0xfd
    "11111111", -- 3384 - 0xd38  :  255 - 0xff -- plane 1
    "11111111", -- 3385 - 0xd39  :  255 - 0xff
    "11111111", -- 3386 - 0xd3a  :  255 - 0xff
    "11111111", -- 3387 - 0xd3b  :  255 - 0xff
    "11111101", -- 3388 - 0xd3c  :  253 - 0xfd
    "11111101", -- 3389 - 0xd3d  :  253 - 0xfd
    "11111101", -- 3390 - 0xd3e  :  253 - 0xfd
    "11111101", -- 3391 - 0xd3f  :  253 - 0xfd
    "11000111", -- 3392 - 0xd40  :  199 - 0xc7 -- Sprite 0xd4
    "11110111", -- 3393 - 0xd41  :  247 - 0xf7
    "11110000", -- 3394 - 0xd42  :  240 - 0xf0
    "11111000", -- 3395 - 0xd43  :  248 - 0xf8
    "11111000", -- 3396 - 0xd44  :  248 - 0xf8
    "11111111", -- 3397 - 0xd45  :  255 - 0xff
    "11111111", -- 3398 - 0xd46  :  255 - 0xff
    "11111111", -- 3399 - 0xd47  :  255 - 0xff
    "00000111", -- 3400 - 0xd48  :    7 - 0x7 -- plane 1
    "00000111", -- 3401 - 0xd49  :    7 - 0x7
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000011", -- 3403 - 0xd4b  :    3 - 0x3
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "11111000", -- 3408 - 0xd50  :  248 - 0xf8 -- Sprite 0xd5
    "11111000", -- 3409 - 0xd51  :  248 - 0xf8
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "11111111", -- 3413 - 0xd55  :  255 - 0xff
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "11111010", -- 3416 - 0xd58  :  250 - 0xfa -- plane 1
    "11111010", -- 3417 - 0xd59  :  250 - 0xfa
    "00000010", -- 3418 - 0xd5a  :    2 - 0x2
    "11111110", -- 3419 - 0xd5b  :  254 - 0xfe
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00000000", -- 3422 - 0xd5e  :    0 - 0x0
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "10001111", -- 3424 - 0xd60  :  143 - 0x8f -- Sprite 0xd6
    "11101111", -- 3425 - 0xd61  :  239 - 0xef
    "11000000", -- 3426 - 0xd62  :  192 - 0xc0
    "11110000", -- 3427 - 0xd63  :  240 - 0xf0
    "11100000", -- 3428 - 0xd64  :  224 - 0xe0
    "11111111", -- 3429 - 0xd65  :  255 - 0xff
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "00001111", -- 3432 - 0xd68  :   15 - 0xf -- plane 1
    "00001111", -- 3433 - 0xd69  :   15 - 0xf
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "00000111", -- 3435 - 0xd6b  :    7 - 0x7
    "00000000", -- 3436 - 0xd6c  :    0 - 0x0
    "00000000", -- 3437 - 0xd6d  :    0 - 0x0
    "00000000", -- 3438 - 0xd6e  :    0 - 0x0
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "11111111", -- 3440 - 0xd70  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "00000000", -- 3442 - 0xd72  :    0 - 0x0
    "00000000", -- 3443 - 0xd73  :    0 - 0x0
    "00000000", -- 3444 - 0xd74  :    0 - 0x0
    "11111111", -- 3445 - 0xd75  :  255 - 0xff
    "11111111", -- 3446 - 0xd76  :  255 - 0xff
    "11111111", -- 3447 - 0xd77  :  255 - 0xff
    "11111111", -- 3448 - 0xd78  :  255 - 0xff -- plane 1
    "11111111", -- 3449 - 0xd79  :  255 - 0xff
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "11111111", -- 3451 - 0xd7b  :  255 - 0xff
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "11000011", -- 3456 - 0xd80  :  195 - 0xc3 -- Sprite 0xd8
    "11111111", -- 3457 - 0xd81  :  255 - 0xff
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000000", -- 3460 - 0xd84  :    0 - 0x0
    "11111111", -- 3461 - 0xd85  :  255 - 0xff
    "11111111", -- 3462 - 0xd86  :  255 - 0xff
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11000011", -- 3464 - 0xd88  :  195 - 0xc3 -- plane 1
    "11111111", -- 3465 - 0xd89  :  255 - 0xff
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "11111111", -- 3467 - 0xd8b  :  255 - 0xff
    "00000000", -- 3468 - 0xd8c  :    0 - 0x0
    "00000000", -- 3469 - 0xd8d  :    0 - 0x0
    "00000000", -- 3470 - 0xd8e  :    0 - 0x0
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00000011", -- 3472 - 0xd90  :    3 - 0x3 -- Sprite 0xd9
    "10000001", -- 3473 - 0xd91  :  129 - 0x81
    "00000000", -- 3474 - 0xd92  :    0 - 0x0
    "00000000", -- 3475 - 0xd93  :    0 - 0x0
    "00000011", -- 3476 - 0xd94  :    3 - 0x3
    "11111111", -- 3477 - 0xd95  :  255 - 0xff
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111111", -- 3479 - 0xd97  :  255 - 0xff
    "01101011", -- 3480 - 0xd98  :  107 - 0x6b -- plane 1
    "10110101", -- 3481 - 0xd99  :  181 - 0xb5
    "00110110", -- 3482 - 0xd9a  :   54 - 0x36
    "11111000", -- 3483 - 0xd9b  :  248 - 0xf8
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000000", -- 3486 - 0xd9e  :    0 - 0x0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "11111111", -- 3488 - 0xda0  :  255 - 0xff -- Sprite 0xda
    "11111111", -- 3489 - 0xda1  :  255 - 0xff
    "01111110", -- 3490 - 0xda2  :  126 - 0x7e
    "00000000", -- 3491 - 0xda3  :    0 - 0x0
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "11100000", -- 3493 - 0xda5  :  224 - 0xe0
    "11111111", -- 3494 - 0xda6  :  255 - 0xff
    "11111111", -- 3495 - 0xda7  :  255 - 0xff
    "11111111", -- 3496 - 0xda8  :  255 - 0xff -- plane 1
    "11111111", -- 3497 - 0xda9  :  255 - 0xff
    "01111110", -- 3498 - 0xdaa  :  126 - 0x7e
    "10000001", -- 3499 - 0xdab  :  129 - 0x81
    "00011111", -- 3500 - 0xdac  :   31 - 0x1f
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "01100001", -- 3504 - 0xdb0  :   97 - 0x61 -- Sprite 0xdb
    "11000011", -- 3505 - 0xdb1  :  195 - 0xc3
    "00000111", -- 3506 - 0xdb2  :    7 - 0x7
    "00001111", -- 3507 - 0xdb3  :   15 - 0xf
    "00011111", -- 3508 - 0xdb4  :   31 - 0x1f
    "01111111", -- 3509 - 0xdb5  :  127 - 0x7f
    "11111111", -- 3510 - 0xdb6  :  255 - 0xff
    "11111111", -- 3511 - 0xdb7  :  255 - 0xff
    "01101100", -- 3512 - 0xdb8  :  108 - 0x6c -- plane 1
    "11011000", -- 3513 - 0xdb9  :  216 - 0xd8
    "00110000", -- 3514 - 0xdba  :   48 - 0x30
    "11100000", -- 3515 - 0xdbb  :  224 - 0xe0
    "10000000", -- 3516 - 0xdbc  :  128 - 0x80
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000000", -- 3518 - 0xdbe  :    0 - 0x0
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00011111", -- 3520 - 0xdc0  :   31 - 0x1f -- Sprite 0xdc
    "11011111", -- 3521 - 0xdc1  :  223 - 0xdf
    "11000000", -- 3522 - 0xdc2  :  192 - 0xc0
    "11110000", -- 3523 - 0xdc3  :  240 - 0xf0
    "11110000", -- 3524 - 0xdc4  :  240 - 0xf0
    "11111111", -- 3525 - 0xdc5  :  255 - 0xff
    "11111111", -- 3526 - 0xdc6  :  255 - 0xff
    "11111111", -- 3527 - 0xdc7  :  255 - 0xff
    "00011111", -- 3528 - 0xdc8  :   31 - 0x1f -- plane 1
    "00011111", -- 3529 - 0xdc9  :   31 - 0x1f
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000111", -- 3531 - 0xdcb  :    7 - 0x7
    "00000000", -- 3532 - 0xdcc  :    0 - 0x0
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "00000000", -- 3534 - 0xdce  :    0 - 0x0
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "10000100", -- 3536 - 0xdd0  :  132 - 0x84 -- Sprite 0xdd
    "11111100", -- 3537 - 0xdd1  :  252 - 0xfc
    "00000000", -- 3538 - 0xdd2  :    0 - 0x0
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "11111111", -- 3541 - 0xdd5  :  255 - 0xff
    "11111111", -- 3542 - 0xdd6  :  255 - 0xff
    "11111111", -- 3543 - 0xdd7  :  255 - 0xff
    "10000101", -- 3544 - 0xdd8  :  133 - 0x85 -- plane 1
    "11111101", -- 3545 - 0xdd9  :  253 - 0xfd
    "00000001", -- 3546 - 0xdda  :    1 - 0x1
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "01111111", -- 3552 - 0xde0  :  127 - 0x7f -- Sprite 0xde
    "01111111", -- 3553 - 0xde1  :  127 - 0x7f
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "11111111", -- 3557 - 0xde5  :  255 - 0xff
    "11111111", -- 3558 - 0xde6  :  255 - 0xff
    "11111111", -- 3559 - 0xde7  :  255 - 0xff
    "01111111", -- 3560 - 0xde8  :  127 - 0x7f -- plane 1
    "01111111", -- 3561 - 0xde9  :  127 - 0x7f
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "01011111", -- 3563 - 0xdeb  :   95 - 0x5f
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "11111100", -- 3568 - 0xdf0  :  252 - 0xfc -- Sprite 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111111", -- 3575 - 0xdf7  :  255 - 0xff
    "11111100", -- 3576 - 0xdf8  :  252 - 0xfc -- plane 1
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00110000", -- 3584 - 0xe00  :   48 - 0x30 -- Sprite 0xe0
    "11110000", -- 3585 - 0xe01  :  240 - 0xf0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "11111111", -- 3589 - 0xe05  :  255 - 0xff
    "11111111", -- 3590 - 0xe06  :  255 - 0xff
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "00110100", -- 3592 - 0xe08  :   52 - 0x34 -- plane 1
    "11110110", -- 3593 - 0xe09  :  246 - 0xf6
    "00000010", -- 3594 - 0xe0a  :    2 - 0x2
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "11111111", -- 3600 - 0xe10  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "11111111", -- 3605 - 0xe15  :  255 - 0xff
    "11111111", -- 3606 - 0xe16  :  255 - 0xff
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "11111111", -- 3608 - 0xe18  :  255 - 0xff -- plane 1
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "01111111", -- 3611 - 0xe1b  :  127 - 0x7f
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "11100001", -- 3616 - 0xe20  :  225 - 0xe1 -- Sprite 0xe2
    "11111111", -- 3617 - 0xe21  :  255 - 0xff
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "11111111", -- 3621 - 0xe25  :  255 - 0xff
    "11111111", -- 3622 - 0xe26  :  255 - 0xff
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11100001", -- 3624 - 0xe28  :  225 - 0xe1 -- plane 1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00011111", -- 3632 - 0xe30  :   31 - 0x1f -- Sprite 0xe3
    "00011111", -- 3633 - 0xe31  :   31 - 0x1f
    "00011111", -- 3634 - 0xe32  :   31 - 0x1f
    "00011111", -- 3635 - 0xe33  :   31 - 0x1f
    "00011111", -- 3636 - 0xe34  :   31 - 0x1f
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "01000000", -- 3640 - 0xe38  :   64 - 0x40 -- plane 1
    "01000000", -- 3641 - 0xe39  :   64 - 0x40
    "01000000", -- 3642 - 0xe3a  :   64 - 0x40
    "11000000", -- 3643 - 0xe3b  :  192 - 0xc0
    "00000000", -- 3644 - 0xe3c  :    0 - 0x0
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Sprite 0xe4
    "00011111", -- 3649 - 0xe41  :   31 - 0x1f
    "00111111", -- 3650 - 0xe42  :   63 - 0x3f
    "01111000", -- 3651 - 0xe43  :  120 - 0x78
    "01110111", -- 3652 - 0xe44  :  119 - 0x77
    "01101111", -- 3653 - 0xe45  :  111 - 0x6f
    "01101111", -- 3654 - 0xe46  :  111 - 0x6f
    "01101111", -- 3655 - 0xe47  :  111 - 0x6f
    "00000000", -- 3656 - 0xe48  :    0 - 0x0 -- plane 1
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000111", -- 3660 - 0xe4c  :    7 - 0x7
    "00001111", -- 3661 - 0xe4d  :   15 - 0xf
    "00001111", -- 3662 - 0xe4e  :   15 - 0xf
    "00001111", -- 3663 - 0xe4f  :   15 - 0xf
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Sprite 0xe5
    "11111000", -- 3665 - 0xe51  :  248 - 0xf8
    "11111100", -- 3666 - 0xe52  :  252 - 0xfc
    "00011110", -- 3667 - 0xe53  :   30 - 0x1e
    "11101110", -- 3668 - 0xe54  :  238 - 0xee
    "11110110", -- 3669 - 0xe55  :  246 - 0xf6
    "11110110", -- 3670 - 0xe56  :  246 - 0xf6
    "11110110", -- 3671 - 0xe57  :  246 - 0xf6
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- plane 1
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "11100000", -- 3676 - 0xe5c  :  224 - 0xe0
    "11110000", -- 3677 - 0xe5d  :  240 - 0xf0
    "11110000", -- 3678 - 0xe5e  :  240 - 0xf0
    "11110000", -- 3679 - 0xe5f  :  240 - 0xf0
    "11110110", -- 3680 - 0xe60  :  246 - 0xf6 -- Sprite 0xe6
    "11110110", -- 3681 - 0xe61  :  246 - 0xf6
    "11110110", -- 3682 - 0xe62  :  246 - 0xf6
    "11101110", -- 3683 - 0xe63  :  238 - 0xee
    "00011110", -- 3684 - 0xe64  :   30 - 0x1e
    "11111100", -- 3685 - 0xe65  :  252 - 0xfc
    "11111000", -- 3686 - 0xe66  :  248 - 0xf8
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "11110000", -- 3688 - 0xe68  :  240 - 0xf0 -- plane 1
    "11110000", -- 3689 - 0xe69  :  240 - 0xf0
    "11110000", -- 3690 - 0xe6a  :  240 - 0xf0
    "11100000", -- 3691 - 0xe6b  :  224 - 0xe0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "01101111", -- 3696 - 0xe70  :  111 - 0x6f -- Sprite 0xe7
    "01101111", -- 3697 - 0xe71  :  111 - 0x6f
    "01101111", -- 3698 - 0xe72  :  111 - 0x6f
    "01110111", -- 3699 - 0xe73  :  119 - 0x77
    "01111000", -- 3700 - 0xe74  :  120 - 0x78
    "00111111", -- 3701 - 0xe75  :   63 - 0x3f
    "00011111", -- 3702 - 0xe76  :   31 - 0x1f
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00001111", -- 3704 - 0xe78  :   15 - 0xf -- plane 1
    "00001111", -- 3705 - 0xe79  :   15 - 0xf
    "00001111", -- 3706 - 0xe7a  :   15 - 0xf
    "00000111", -- 3707 - 0xe7b  :    7 - 0x7
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Sprite 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- plane 1
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11110110", -- 3728 - 0xe90  :  246 - 0xf6 -- Sprite 0xe9
    "11110110", -- 3729 - 0xe91  :  246 - 0xf6
    "11110110", -- 3730 - 0xe92  :  246 - 0xf6
    "11110110", -- 3731 - 0xe93  :  246 - 0xf6
    "11110110", -- 3732 - 0xe94  :  246 - 0xf6
    "11110110", -- 3733 - 0xe95  :  246 - 0xf6
    "11110110", -- 3734 - 0xe96  :  246 - 0xf6
    "11110110", -- 3735 - 0xe97  :  246 - 0xf6
    "11110000", -- 3736 - 0xe98  :  240 - 0xf0 -- plane 1
    "11110000", -- 3737 - 0xe99  :  240 - 0xf0
    "11110000", -- 3738 - 0xe9a  :  240 - 0xf0
    "11110000", -- 3739 - 0xe9b  :  240 - 0xf0
    "11110000", -- 3740 - 0xe9c  :  240 - 0xf0
    "11110000", -- 3741 - 0xe9d  :  240 - 0xf0
    "11110000", -- 3742 - 0xe9e  :  240 - 0xf0
    "11110000", -- 3743 - 0xe9f  :  240 - 0xf0
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "11111111", -- 3752 - 0xea8  :  255 - 0xff -- plane 1
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "01101111", -- 3760 - 0xeb0  :  111 - 0x6f -- Sprite 0xeb
    "01101111", -- 3761 - 0xeb1  :  111 - 0x6f
    "01101111", -- 3762 - 0xeb2  :  111 - 0x6f
    "01101111", -- 3763 - 0xeb3  :  111 - 0x6f
    "01101111", -- 3764 - 0xeb4  :  111 - 0x6f
    "01101111", -- 3765 - 0xeb5  :  111 - 0x6f
    "01101111", -- 3766 - 0xeb6  :  111 - 0x6f
    "01101111", -- 3767 - 0xeb7  :  111 - 0x6f
    "00001111", -- 3768 - 0xeb8  :   15 - 0xf -- plane 1
    "00001111", -- 3769 - 0xeb9  :   15 - 0xf
    "00001111", -- 3770 - 0xeba  :   15 - 0xf
    "00001111", -- 3771 - 0xebb  :   15 - 0xf
    "00001111", -- 3772 - 0xebc  :   15 - 0xf
    "00001111", -- 3773 - 0xebd  :   15 - 0xf
    "00001111", -- 3774 - 0xebe  :   15 - 0xf
    "00001111", -- 3775 - 0xebf  :   15 - 0xf
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0 -- plane 1
    "00000000", -- 3801 - 0xed9  :    0 - 0x0
    "00000000", -- 3802 - 0xeda  :    0 - 0x0
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- plane 1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "00000000", -- 3828 - 0xef4  :    0 - 0x0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "00000000", -- 3830 - 0xef6  :    0 - 0x0
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "00000000", -- 3832 - 0xef8  :    0 - 0x0 -- plane 1
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "11111111", -- 3840 - 0xf00  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 3841 - 0xf01  :  255 - 0xff
    "11111111", -- 3842 - 0xf02  :  255 - 0xff
    "11111111", -- 3843 - 0xf03  :  255 - 0xff
    "11111111", -- 3844 - 0xf04  :  255 - 0xff
    "11111111", -- 3845 - 0xf05  :  255 - 0xff
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11111111", -- 3848 - 0xf08  :  255 - 0xff -- plane 1
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "11111111", -- 3850 - 0xf0a  :  255 - 0xff
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "11111111", -- 3860 - 0xf14  :  255 - 0xff
    "11111111", -- 3861 - 0xf15  :  255 - 0xff
    "11111111", -- 3862 - 0xf16  :  255 - 0xff
    "11111111", -- 3863 - 0xf17  :  255 - 0xff
    "11111111", -- 3864 - 0xf18  :  255 - 0xff -- plane 1
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11111111", -- 3867 - 0xf1b  :  255 - 0xff
    "11111111", -- 3868 - 0xf1c  :  255 - 0xff
    "11111111", -- 3869 - 0xf1d  :  255 - 0xff
    "11111111", -- 3870 - 0xf1e  :  255 - 0xff
    "11111111", -- 3871 - 0xf1f  :  255 - 0xff
    "11111111", -- 3872 - 0xf20  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 3873 - 0xf21  :  255 - 0xff
    "11111111", -- 3874 - 0xf22  :  255 - 0xff
    "11111111", -- 3875 - 0xf23  :  255 - 0xff
    "11111111", -- 3876 - 0xf24  :  255 - 0xff
    "11111111", -- 3877 - 0xf25  :  255 - 0xff
    "11111111", -- 3878 - 0xf26  :  255 - 0xff
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff -- plane 1
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11111111", -- 3883 - 0xf2b  :  255 - 0xff
    "11111111", -- 3884 - 0xf2c  :  255 - 0xff
    "11111111", -- 3885 - 0xf2d  :  255 - 0xff
    "11111111", -- 3886 - 0xf2e  :  255 - 0xff
    "11111111", -- 3887 - 0xf2f  :  255 - 0xff
    "11111111", -- 3888 - 0xf30  :  255 - 0xff -- Sprite 0xf3
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "11111111", -- 3891 - 0xf33  :  255 - 0xff
    "11111111", -- 3892 - 0xf34  :  255 - 0xff
    "11111111", -- 3893 - 0xf35  :  255 - 0xff
    "11111111", -- 3894 - 0xf36  :  255 - 0xff
    "11111111", -- 3895 - 0xf37  :  255 - 0xff
    "11111111", -- 3896 - 0xf38  :  255 - 0xff -- plane 1
    "11111111", -- 3897 - 0xf39  :  255 - 0xff
    "11111111", -- 3898 - 0xf3a  :  255 - 0xff
    "11111111", -- 3899 - 0xf3b  :  255 - 0xff
    "11111111", -- 3900 - 0xf3c  :  255 - 0xff
    "11111111", -- 3901 - 0xf3d  :  255 - 0xff
    "11111111", -- 3902 - 0xf3e  :  255 - 0xff
    "11111111", -- 3903 - 0xf3f  :  255 - 0xff
    "11111111", -- 3904 - 0xf40  :  255 - 0xff -- Sprite 0xf4
    "11111111", -- 3905 - 0xf41  :  255 - 0xff
    "11111111", -- 3906 - 0xf42  :  255 - 0xff
    "11111111", -- 3907 - 0xf43  :  255 - 0xff
    "11111111", -- 3908 - 0xf44  :  255 - 0xff
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "11111111", -- 3912 - 0xf48  :  255 - 0xff -- plane 1
    "11111111", -- 3913 - 0xf49  :  255 - 0xff
    "11111111", -- 3914 - 0xf4a  :  255 - 0xff
    "11111111", -- 3915 - 0xf4b  :  255 - 0xff
    "11111111", -- 3916 - 0xf4c  :  255 - 0xff
    "11111111", -- 3917 - 0xf4d  :  255 - 0xff
    "11111111", -- 3918 - 0xf4e  :  255 - 0xff
    "11111111", -- 3919 - 0xf4f  :  255 - 0xff
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Sprite 0xf5
    "11111111", -- 3921 - 0xf51  :  255 - 0xff
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "11111111", -- 3923 - 0xf53  :  255 - 0xff
    "11111111", -- 3924 - 0xf54  :  255 - 0xff
    "11111111", -- 3925 - 0xf55  :  255 - 0xff
    "11111111", -- 3926 - 0xf56  :  255 - 0xff
    "11111111", -- 3927 - 0xf57  :  255 - 0xff
    "11111111", -- 3928 - 0xf58  :  255 - 0xff -- plane 1
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "11111111", -- 3931 - 0xf5b  :  255 - 0xff
    "11111111", -- 3932 - 0xf5c  :  255 - 0xff
    "11111111", -- 3933 - 0xf5d  :  255 - 0xff
    "11111111", -- 3934 - 0xf5e  :  255 - 0xff
    "11111111", -- 3935 - 0xf5f  :  255 - 0xff
    "11111111", -- 3936 - 0xf60  :  255 - 0xff -- Sprite 0xf6
    "11111111", -- 3937 - 0xf61  :  255 - 0xff
    "11111111", -- 3938 - 0xf62  :  255 - 0xff
    "11111111", -- 3939 - 0xf63  :  255 - 0xff
    "11111111", -- 3940 - 0xf64  :  255 - 0xff
    "11111111", -- 3941 - 0xf65  :  255 - 0xff
    "11111111", -- 3942 - 0xf66  :  255 - 0xff
    "11111111", -- 3943 - 0xf67  :  255 - 0xff
    "11111111", -- 3944 - 0xf68  :  255 - 0xff -- plane 1
    "11111111", -- 3945 - 0xf69  :  255 - 0xff
    "11111111", -- 3946 - 0xf6a  :  255 - 0xff
    "11111111", -- 3947 - 0xf6b  :  255 - 0xff
    "11111111", -- 3948 - 0xf6c  :  255 - 0xff
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "11111111", -- 3952 - 0xf70  :  255 - 0xff -- Sprite 0xf7
    "11111111", -- 3953 - 0xf71  :  255 - 0xff
    "11111111", -- 3954 - 0xf72  :  255 - 0xff
    "11111111", -- 3955 - 0xf73  :  255 - 0xff
    "11111111", -- 3956 - 0xf74  :  255 - 0xff
    "11111111", -- 3957 - 0xf75  :  255 - 0xff
    "11111111", -- 3958 - 0xf76  :  255 - 0xff
    "11111111", -- 3959 - 0xf77  :  255 - 0xff
    "11111111", -- 3960 - 0xf78  :  255 - 0xff -- plane 1
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "11111111", -- 3968 - 0xf80  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "11111111", -- 3970 - 0xf82  :  255 - 0xff
    "11111111", -- 3971 - 0xf83  :  255 - 0xff
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "11111111", -- 3974 - 0xf86  :  255 - 0xff
    "11111111", -- 3975 - 0xf87  :  255 - 0xff
    "11111111", -- 3976 - 0xf88  :  255 - 0xff -- plane 1
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111111", -- 3982 - 0xf8e  :  255 - 0xff
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "11111111", -- 3992 - 0xf98  :  255 - 0xff -- plane 1
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111111", -- 3999 - 0xf9f  :  255 - 0xff
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "11111111", -- 4007 - 0xfa7  :  255 - 0xff
    "11111111", -- 4008 - 0xfa8  :  255 - 0xff -- plane 1
    "11111111", -- 4009 - 0xfa9  :  255 - 0xff
    "11111111", -- 4010 - 0xfaa  :  255 - 0xff
    "11111111", -- 4011 - 0xfab  :  255 - 0xff
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "11111111", -- 4015 - 0xfaf  :  255 - 0xff
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "11111111", -- 4024 - 0xfb8  :  255 - 0xff -- plane 1
    "11111111", -- 4025 - 0xfb9  :  255 - 0xff
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "11111111", -- 4031 - 0xfbf  :  255 - 0xff
    "11111111", -- 4032 - 0xfc0  :  255 - 0xff -- Sprite 0xfc
    "11111111", -- 4033 - 0xfc1  :  255 - 0xff
    "11111111", -- 4034 - 0xfc2  :  255 - 0xff
    "11111111", -- 4035 - 0xfc3  :  255 - 0xff
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "11111111", -- 4040 - 0xfc8  :  255 - 0xff -- plane 1
    "11111111", -- 4041 - 0xfc9  :  255 - 0xff
    "11111111", -- 4042 - 0xfca  :  255 - 0xff
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "11111111", -- 4048 - 0xfd0  :  255 - 0xff -- Sprite 0xfd
    "11111111", -- 4049 - 0xfd1  :  255 - 0xff
    "11111111", -- 4050 - 0xfd2  :  255 - 0xff
    "11111111", -- 4051 - 0xfd3  :  255 - 0xff
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff -- plane 1
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "11111111", -- 4064 - 0xfe0  :  255 - 0xff -- Sprite 0xfe
    "11111111", -- 4065 - 0xfe1  :  255 - 0xff
    "11111111", -- 4066 - 0xfe2  :  255 - 0xff
    "11111111", -- 4067 - 0xfe3  :  255 - 0xff
    "11111111", -- 4068 - 0xfe4  :  255 - 0xff
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff -- plane 1
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11111111", -- 4075 - 0xfeb  :  255 - 0xff
    "11111111", -- 4076 - 0xfec  :  255 - 0xff
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff -- plane 1
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
