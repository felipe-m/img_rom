---   Sprites Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: lawnmower_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_LAWN_SPR_PLN0 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_LAWN_SPR_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_LAWN_SPR_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table COLOR PLANE 0
    "11111111", --    0 -  0x0  :  255 - 0xff -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11111111", --    2 -  0x2  :  255 - 0xff
    "11111111", --    3 -  0x3  :  255 - 0xff
    "11111111", --    4 -  0x4  :  255 - 0xff
    "11111111", --    5 -  0x5  :  255 - 0xff
    "11111111", --    6 -  0x6  :  255 - 0xff
    "11111111", --    7 -  0x7  :  255 - 0xff
    "11111111", --    8 -  0x8  :  255 - 0xff -- Sprite 0x1
    "11111111", --    9 -  0x9  :  255 - 0xff
    "11111111", --   10 -  0xa  :  255 - 0xff
    "11111111", --   11 -  0xb  :  255 - 0xff
    "11111111", --   12 -  0xc  :  255 - 0xff
    "11111111", --   13 -  0xd  :  255 - 0xff
    "11111100", --   14 -  0xe  :  252 - 0xfc
    "11111100", --   15 -  0xf  :  252 - 0xfc
    "11111111", --   16 - 0x10  :  255 - 0xff -- Sprite 0x2
    "11111111", --   17 - 0x11  :  255 - 0xff
    "11111111", --   18 - 0x12  :  255 - 0xff
    "11111111", --   19 - 0x13  :  255 - 0xff
    "11111111", --   20 - 0x14  :  255 - 0xff
    "11111111", --   21 - 0x15  :  255 - 0xff
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "11111111", --   24 - 0x18  :  255 - 0xff -- Sprite 0x3
    "11111111", --   25 - 0x19  :  255 - 0xff
    "11111111", --   26 - 0x1a  :  255 - 0xff
    "11111111", --   27 - 0x1b  :  255 - 0xff
    "11111111", --   28 - 0x1c  :  255 - 0xff
    "11111111", --   29 - 0x1d  :  255 - 0xff
    "00011111", --   30 - 0x1e  :   31 - 0x1f
    "01000111", --   31 - 0x1f  :   71 - 0x47
    "11111111", --   32 - 0x20  :  255 - 0xff -- Sprite 0x4
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "11111111", --   36 - 0x24  :  255 - 0xff
    "11111111", --   37 - 0x25  :  255 - 0xff
    "11100000", --   38 - 0x26  :  224 - 0xe0
    "10000000", --   39 - 0x27  :  128 - 0x80
    "11111111", --   40 - 0x28  :  255 - 0xff -- Sprite 0x5
    "11111111", --   41 - 0x29  :  255 - 0xff
    "11111111", --   42 - 0x2a  :  255 - 0xff
    "11111111", --   43 - 0x2b  :  255 - 0xff
    "11111111", --   44 - 0x2c  :  255 - 0xff
    "11110111", --   45 - 0x2d  :  247 - 0xf7
    "00000001", --   46 - 0x2e  :    1 - 0x1
    "00000100", --   47 - 0x2f  :    4 - 0x4
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0x6
    "11111111", --   49 - 0x31  :  255 - 0xff
    "11111111", --   50 - 0x32  :  255 - 0xff
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111111", --   52 - 0x34  :  255 - 0xff
    "11011111", --   53 - 0x35  :  223 - 0xdf
    "00011100", --   54 - 0x36  :   28 - 0x1c
    "01000100", --   55 - 0x37  :   68 - 0x44
    "11111111", --   56 - 0x38  :  255 - 0xff -- Sprite 0x7
    "11111111", --   57 - 0x39  :  255 - 0xff
    "11111111", --   58 - 0x3a  :  255 - 0xff
    "11111111", --   59 - 0x3b  :  255 - 0xff
    "11111111", --   60 - 0x3c  :  255 - 0xff
    "10111111", --   61 - 0x3d  :  191 - 0xbf
    "00111100", --   62 - 0x3e  :   60 - 0x3c
    "01001100", --   63 - 0x3f  :   76 - 0x4c
    "11111100", --   64 - 0x40  :  252 - 0xfc -- Sprite 0x8
    "11111100", --   65 - 0x41  :  252 - 0xfc
    "11111100", --   66 - 0x42  :  252 - 0xfc
    "11111100", --   67 - 0x43  :  252 - 0xfc
    "11111100", --   68 - 0x44  :  252 - 0xfc
    "11111100", --   69 - 0x45  :  252 - 0xfc
    "11111100", --   70 - 0x46  :  252 - 0xfc
    "11111100", --   71 - 0x47  :  252 - 0xfc
    "00010000", --   72 - 0x48  :   16 - 0x10 -- Sprite 0x9
    "00111000", --   73 - 0x49  :   56 - 0x38
    "01111100", --   74 - 0x4a  :  124 - 0x7c
    "11111000", --   75 - 0x4b  :  248 - 0xf8
    "01110000", --   76 - 0x4c  :  112 - 0x70
    "00100010", --   77 - 0x4d  :   34 - 0x22
    "00000101", --   78 - 0x4e  :    5 - 0x5
    "00000010", --   79 - 0x4f  :    2 - 0x2
    "01000111", --   80 - 0x50  :   71 - 0x47 -- Sprite 0xa
    "01000111", --   81 - 0x51  :   71 - 0x47
    "01000111", --   82 - 0x52  :   71 - 0x47
    "01000111", --   83 - 0x53  :   71 - 0x47
    "01000111", --   84 - 0x54  :   71 - 0x47
    "01000111", --   85 - 0x55  :   71 - 0x47
    "01000111", --   86 - 0x56  :   71 - 0x47
    "01000111", --   87 - 0x57  :   71 - 0x47
    "11111111", --   88 - 0x58  :  255 - 0xff -- Sprite 0xb
    "11111110", --   89 - 0x59  :  254 - 0xfe
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111100", --   91 - 0x5b  :  252 - 0xfc
    "11111100", --   92 - 0x5c  :  252 - 0xfc
    "11111100", --   93 - 0x5d  :  252 - 0xfc
    "11111100", --   94 - 0x5e  :  252 - 0xfc
    "11111100", --   95 - 0x5f  :  252 - 0xfc
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0xc
    "00001000", --   97 - 0x61  :    8 - 0x8
    "00011100", --   98 - 0x62  :   28 - 0x1c
    "00111000", --   99 - 0x63  :   56 - 0x38
    "01110000", --  100 - 0x64  :  112 - 0x70
    "00100010", --  101 - 0x65  :   34 - 0x22
    "00000101", --  102 - 0x66  :    5 - 0x5
    "00000010", --  103 - 0x67  :    2 - 0x2
    "00000010", --  104 - 0x68  :    2 - 0x2 -- Sprite 0xd
    "00110001", --  105 - 0x69  :   49 - 0x31
    "01111000", --  106 - 0x6a  :  120 - 0x78
    "11111000", --  107 - 0x6b  :  248 - 0xf8
    "01110000", --  108 - 0x6c  :  112 - 0x70
    "00100010", --  109 - 0x6d  :   34 - 0x22
    "00000101", --  110 - 0x6e  :    5 - 0x5
    "00000010", --  111 - 0x6f  :    2 - 0x2
    "01111100", --  112 - 0x70  :  124 - 0x7c -- Sprite 0xe
    "00111100", --  113 - 0x71  :   60 - 0x3c
    "10011100", --  114 - 0x72  :  156 - 0x9c
    "10001100", --  115 - 0x73  :  140 - 0x8c
    "01001100", --  116 - 0x74  :   76 - 0x4c
    "01000100", --  117 - 0x75  :   68 - 0x44
    "01000100", --  118 - 0x76  :   68 - 0x44
    "01000100", --  119 - 0x77  :   68 - 0x44
    "01000100", --  120 - 0x78  :   68 - 0x44 -- Sprite 0xf
    "01000100", --  121 - 0x79  :   68 - 0x44
    "01000100", --  122 - 0x7a  :   68 - 0x44
    "01000100", --  123 - 0x7b  :   68 - 0x44
    "01000100", --  124 - 0x7c  :   68 - 0x44
    "01000100", --  125 - 0x7d  :   68 - 0x44
    "01000100", --  126 - 0x7e  :   68 - 0x44
    "01000100", --  127 - 0x7f  :   68 - 0x44
    "01001100", --  128 - 0x80  :   76 - 0x4c -- Sprite 0x10
    "00100100", --  129 - 0x81  :   36 - 0x24
    "00100100", --  130 - 0x82  :   36 - 0x24
    "10010100", --  131 - 0x83  :  148 - 0x94
    "00010000", --  132 - 0x84  :   16 - 0x10
    "00001000", --  133 - 0x85  :    8 - 0x8
    "00001000", --  134 - 0x86  :    8 - 0x8
    "00000100", --  135 - 0x87  :    4 - 0x4
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x11
    "00111100", --  137 - 0x89  :   60 - 0x3c
    "01000000", --  138 - 0x8a  :   64 - 0x40
    "01000100", --  139 - 0x8b  :   68 - 0x44
    "01000100", --  140 - 0x8c  :   68 - 0x44
    "01000100", --  141 - 0x8d  :   68 - 0x44
    "01000100", --  142 - 0x8e  :   68 - 0x44
    "01000100", --  143 - 0x8f  :   68 - 0x44
    "00000100", --  144 - 0x90  :    4 - 0x4 -- Sprite 0x12
    "00010010", --  145 - 0x91  :   18 - 0x12
    "00110010", --  146 - 0x92  :   50 - 0x32
    "01111000", --  147 - 0x93  :  120 - 0x78
    "11111000", --  148 - 0x94  :  248 - 0xf8
    "01110000", --  149 - 0x95  :  112 - 0x70
    "00100100", --  150 - 0x96  :   36 - 0x24
    "00000000", --  151 - 0x97  :    0 - 0x0
    "01000100", --  152 - 0x98  :   68 - 0x44 -- Sprite 0x13
    "01000100", --  153 - 0x99  :   68 - 0x44
    "01000100", --  154 - 0x9a  :   68 - 0x44
    "01000100", --  155 - 0x9b  :   68 - 0x44
    "01000100", --  156 - 0x9c  :   68 - 0x44
    "01000100", --  157 - 0x9d  :   68 - 0x44
    "01000100", --  158 - 0x9e  :   68 - 0x44
    "01011100", --  159 - 0x9f  :   92 - 0x5c
    "00010000", --  160 - 0xa0  :   16 - 0x10 -- Sprite 0x14
    "00111000", --  161 - 0xa1  :   56 - 0x38
    "00111100", --  162 - 0xa2  :   60 - 0x3c
    "00111000", --  163 - 0xa3  :   56 - 0x38
    "00010000", --  164 - 0xa4  :   16 - 0x10
    "00000010", --  165 - 0xa5  :    2 - 0x2
    "01000101", --  166 - 0xa6  :   69 - 0x45
    "01000010", --  167 - 0xa7  :   66 - 0x42
    "01000100", --  168 - 0xa8  :   68 - 0x44 -- Sprite 0x15
    "01000100", --  169 - 0xa9  :   68 - 0x44
    "01000100", --  170 - 0xaa  :   68 - 0x44
    "01000100", --  171 - 0xab  :   68 - 0x44
    "01000100", --  172 - 0xac  :   68 - 0x44
    "01011100", --  173 - 0xad  :   92 - 0x5c
    "01000000", --  174 - 0xae  :   64 - 0x40
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "01000000", --  176 - 0xb0  :   64 - 0x40 -- Sprite 0x16
    "01000000", --  177 - 0xb1  :   64 - 0x40
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00011000", --  180 - 0xb4  :   24 - 0x18
    "00111000", --  181 - 0xb5  :   56 - 0x38
    "00010000", --  182 - 0xb6  :   16 - 0x10
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "01000000", --  184 - 0xb8  :   64 - 0x40 -- Sprite 0x17
    "01000000", --  185 - 0xb9  :   64 - 0x40
    "01000000", --  186 - 0xba  :   64 - 0x40
    "01000000", --  187 - 0xbb  :   64 - 0x40
    "01010000", --  188 - 0xbc  :   80 - 0x50
    "01010000", --  189 - 0xbd  :   80 - 0x50
    "01001000", --  190 - 0xbe  :   72 - 0x48
    "01001000", --  191 - 0xbf  :   72 - 0x48
    "01000111", --  192 - 0xc0  :   71 - 0x47 -- Sprite 0x18
    "01000111", --  193 - 0xc1  :   71 - 0x47
    "01000111", --  194 - 0xc2  :   71 - 0x47
    "01000111", --  195 - 0xc3  :   71 - 0x47
    "01000111", --  196 - 0xc4  :   71 - 0x47
    "01011111", --  197 - 0xc5  :   95 - 0x5f
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "11111100", --  200 - 0xc8  :  252 - 0xfc -- Sprite 0x19
    "11111100", --  201 - 0xc9  :  252 - 0xfc
    "11111100", --  202 - 0xca  :  252 - 0xfc
    "11111100", --  203 - 0xcb  :  252 - 0xfc
    "11111100", --  204 - 0xcc  :  252 - 0xfc
    "11011100", --  205 - 0xcd  :  220 - 0xdc
    "00011100", --  206 - 0xce  :   28 - 0x1c
    "01000100", --  207 - 0xcf  :   68 - 0x44
    "00010000", --  208 - 0xd0  :   16 - 0x10 -- Sprite 0x1a
    "00111000", --  209 - 0xd1  :   56 - 0x38
    "01111100", --  210 - 0xd2  :  124 - 0x7c
    "11100000", --  211 - 0xd3  :  224 - 0xe0
    "01000000", --  212 - 0xd4  :   64 - 0x40
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00010000", --  214 - 0xd6  :   16 - 0x10
    "00100000", --  215 - 0xd7  :   32 - 0x20
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "01111100", --  217 - 0xd9  :  124 - 0x7c
    "01000000", --  218 - 0xda  :   64 - 0x40
    "01000100", --  219 - 0xdb  :   68 - 0x44
    "01000100", --  220 - 0xdc  :   68 - 0x44
    "01000100", --  221 - 0xdd  :   68 - 0x44
    "01000100", --  222 - 0xde  :   68 - 0x44
    "01000100", --  223 - 0xdf  :   68 - 0x44
    "00010000", --  224 - 0xe0  :   16 - 0x10 -- Sprite 0x1c
    "00111000", --  225 - 0xe1  :   56 - 0x38
    "01110001", --  226 - 0xe2  :  113 - 0x71
    "11100010", --  227 - 0xe3  :  226 - 0xe2
    "01000100", --  228 - 0xe4  :   68 - 0x44
    "00001000", --  229 - 0xe5  :    8 - 0x8
    "00010000", --  230 - 0xe6  :   16 - 0x10
    "00100000", --  231 - 0xe7  :   32 - 0x20
    "01000000", --  232 - 0xe8  :   64 - 0x40 -- Sprite 0x1d
    "10000100", --  233 - 0xe9  :  132 - 0x84
    "00000010", --  234 - 0xea  :    2 - 0x2
    "00000111", --  235 - 0xeb  :    7 - 0x7
    "00001111", --  236 - 0xec  :   15 - 0xf
    "00011111", --  237 - 0xed  :   31 - 0x1f
    "00111111", --  238 - 0xee  :   63 - 0x3f
    "01111111", --  239 - 0xef  :  127 - 0x7f
    "00010000", --  240 - 0xf0  :   16 - 0x10 -- Sprite 0x1e
    "00011000", --  241 - 0xf1  :   24 - 0x18
    "00001100", --  242 - 0xf2  :   12 - 0xc
    "00000110", --  243 - 0xf3  :    6 - 0x6
    "10000000", --  244 - 0xf4  :  128 - 0x80
    "11000000", --  245 - 0xf5  :  192 - 0xc0
    "11100000", --  246 - 0xf6  :  224 - 0xe0
    "11110000", --  247 - 0xf7  :  240 - 0xf0
    "11111100", --  248 - 0xf8  :  252 - 0xfc -- Sprite 0x1f
    "11111101", --  249 - 0xf9  :  253 - 0xfd
    "11111100", --  250 - 0xfa  :  252 - 0xfc
    "11111110", --  251 - 0xfb  :  254 - 0xfe
    "11111110", --  252 - 0xfc  :  254 - 0xfe
    "11111111", --  253 - 0xfd  :  255 - 0xff
    "11111111", --  254 - 0xfe  :  255 - 0xff
    "11111111", --  255 - 0xff  :  255 - 0xff
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "11111111", --  257 - 0x101  :  255 - 0xff
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11111111", --  262 - 0x106  :  255 - 0xff
    "11111111", --  263 - 0x107  :  255 - 0xff
    "01000100", --  264 - 0x108  :   68 - 0x44 -- Sprite 0x21
    "11000101", --  265 - 0x109  :  197 - 0xc5
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000110", --  267 - 0x10b  :    6 - 0x6
    "00000110", --  268 - 0x10c  :    6 - 0x6
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "01000000", --  272 - 0x110  :   64 - 0x40 -- Sprite 0x22
    "10000001", --  273 - 0x111  :  129 - 0x81
    "00000011", --  274 - 0x112  :    3 - 0x3
    "00000111", --  275 - 0x113  :    7 - 0x7
    "00001111", --  276 - 0x114  :   15 - 0xf
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11111111", --  278 - 0x116  :  255 - 0xff
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111000", --  280 - 0x118  :  248 - 0xf8 -- Sprite 0x23
    "11111100", --  281 - 0x119  :  252 - 0xfc
    "11111110", --  282 - 0x11a  :  254 - 0xfe
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111111", --  284 - 0x11c  :  255 - 0xff
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11111111", --  286 - 0x11e  :  255 - 0xff
    "11111111", --  287 - 0x11f  :  255 - 0xff
    "01000111", --  288 - 0x120  :   71 - 0x47 -- Sprite 0x24
    "11000111", --  289 - 0x121  :  199 - 0xc7
    "00000111", --  290 - 0x122  :    7 - 0x7
    "00000111", --  291 - 0x123  :    7 - 0x7
    "00000111", --  292 - 0x124  :    7 - 0x7
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11111111", --  294 - 0x126  :  255 - 0xff
    "11111111", --  295 - 0x127  :  255 - 0xff
    "11111111", --  296 - 0x128  :  255 - 0xff -- Sprite 0x25
    "11111111", --  297 - 0x129  :  255 - 0xff
    "11111111", --  298 - 0x12a  :  255 - 0xff
    "11111111", --  299 - 0x12b  :  255 - 0xff
    "11111111", --  300 - 0x12c  :  255 - 0xff
    "11111111", --  301 - 0x12d  :  255 - 0xff
    "00011111", --  302 - 0x12e  :   31 - 0x1f
    "00001111", --  303 - 0x12f  :   15 - 0xf
    "11111111", --  304 - 0x130  :  255 - 0xff -- Sprite 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11111100", --  310 - 0x136  :  252 - 0xfc
    "11111000", --  311 - 0x137  :  248 - 0xf8
    "00100111", --  312 - 0x138  :   39 - 0x27 -- Sprite 0x27
    "00010011", --  313 - 0x139  :   19 - 0x13
    "00001001", --  314 - 0x13a  :    9 - 0x9
    "11000100", --  315 - 0x13b  :  196 - 0xc4
    "01100010", --  316 - 0x13c  :   98 - 0x62
    "00100001", --  317 - 0x13d  :   33 - 0x21
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "11111111", --  320 - 0x140  :  255 - 0xff -- Sprite 0x28
    "11111111", --  321 - 0x141  :  255 - 0xff
    "11111111", --  322 - 0x142  :  255 - 0xff
    "11111111", --  323 - 0x143  :  255 - 0xff
    "01111111", --  324 - 0x144  :  127 - 0x7f
    "00111110", --  325 - 0x145  :   62 - 0x3e
    "10011100", --  326 - 0x146  :  156 - 0x9c
    "01001000", --  327 - 0x147  :   72 - 0x48
    "11110000", --  328 - 0x148  :  240 - 0xf0 -- Sprite 0x29
    "11100000", --  329 - 0x149  :  224 - 0xe0
    "11000000", --  330 - 0x14a  :  192 - 0xc0
    "10000000", --  331 - 0x14b  :  128 - 0x80
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000010", --  333 - 0x14d  :    2 - 0x2
    "00000101", --  334 - 0x14e  :    5 - 0x5
    "00000010", --  335 - 0x14f  :    2 - 0x2
    "01000111", --  336 - 0x150  :   71 - 0x47 -- Sprite 0x2a
    "01000110", --  337 - 0x151  :   70 - 0x46
    "01000110", --  338 - 0x152  :   70 - 0x46
    "01000100", --  339 - 0x153  :   68 - 0x44
    "01000100", --  340 - 0x154  :   68 - 0x44
    "01000100", --  341 - 0x155  :   68 - 0x44
    "01000100", --  342 - 0x156  :   68 - 0x44
    "01000100", --  343 - 0x157  :   68 - 0x44
    "01111111", --  344 - 0x158  :  127 - 0x7f -- Sprite 0x2b
    "00111111", --  345 - 0x159  :   63 - 0x3f
    "10011111", --  346 - 0x15a  :  159 - 0x9f
    "10001111", --  347 - 0x15b  :  143 - 0x8f
    "01001111", --  348 - 0x15c  :   79 - 0x4f
    "01000111", --  349 - 0x15d  :   71 - 0x47
    "01000111", --  350 - 0x15e  :   71 - 0x47
    "01000111", --  351 - 0x15f  :   71 - 0x47
    "00100000", --  352 - 0x160  :   32 - 0x20 -- Sprite 0x2c
    "00010000", --  353 - 0x161  :   16 - 0x10
    "00000000", --  354 - 0x162  :    0 - 0x0
    "11000000", --  355 - 0x163  :  192 - 0xc0
    "01100000", --  356 - 0x164  :   96 - 0x60
    "00100010", --  357 - 0x165  :   34 - 0x22
    "00000101", --  358 - 0x166  :    5 - 0x5
    "00000010", --  359 - 0x167  :    2 - 0x2
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Sprite 0x2d
    "01111111", --  361 - 0x169  :  127 - 0x7f
    "01000000", --  362 - 0x16a  :   64 - 0x40
    "01000000", --  363 - 0x16b  :   64 - 0x40
    "01000000", --  364 - 0x16c  :   64 - 0x40
    "01000111", --  365 - 0x16d  :   71 - 0x47
    "01000111", --  366 - 0x16e  :   71 - 0x47
    "01000111", --  367 - 0x16f  :   71 - 0x47
    "01000100", --  368 - 0x170  :   68 - 0x44 -- Sprite 0x2e
    "11000100", --  369 - 0x171  :  196 - 0xc4
    "00000100", --  370 - 0x172  :    4 - 0x4
    "00000100", --  371 - 0x173  :    4 - 0x4
    "00000100", --  372 - 0x174  :    4 - 0x4
    "11111100", --  373 - 0x175  :  252 - 0xfc
    "11111100", --  374 - 0x176  :  252 - 0xfc
    "11111100", --  375 - 0x177  :  252 - 0xfc
    "00000001", --  376 - 0x178  :    1 - 0x1 -- Sprite 0x2f
    "01111100", --  377 - 0x179  :  124 - 0x7c
    "01000000", --  378 - 0x17a  :   64 - 0x40
    "01000100", --  379 - 0x17b  :   68 - 0x44
    "01000100", --  380 - 0x17c  :   68 - 0x44
    "01000100", --  381 - 0x17d  :   68 - 0x44
    "01000100", --  382 - 0x17e  :   68 - 0x44
    "01000100", --  383 - 0x17f  :   68 - 0x44
    "00010000", --  384 - 0x180  :   16 - 0x10 -- Sprite 0x30
    "00111000", --  385 - 0x181  :   56 - 0x38
    "00111100", --  386 - 0x182  :   60 - 0x3c
    "00011000", --  387 - 0x183  :   24 - 0x18
    "00000000", --  388 - 0x184  :    0 - 0x0
    "01000010", --  389 - 0x185  :   66 - 0x42
    "01000100", --  390 - 0x186  :   68 - 0x44
    "01001000", --  391 - 0x187  :   72 - 0x48
    "01000111", --  392 - 0x188  :   71 - 0x47 -- Sprite 0x31
    "01011111", --  393 - 0x189  :   95 - 0x5f
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "01110000", --  396 - 0x18c  :  112 - 0x70
    "00100010", --  397 - 0x18d  :   34 - 0x22
    "00000101", --  398 - 0x18e  :    5 - 0x5
    "00000010", --  399 - 0x18f  :    2 - 0x2
    "11111111", --  400 - 0x190  :  255 - 0xff -- Sprite 0x32
    "11111111", --  401 - 0x191  :  255 - 0xff
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "01110000", --  404 - 0x194  :  112 - 0x70
    "00100010", --  405 - 0x195  :   34 - 0x22
    "00000101", --  406 - 0x196  :    5 - 0x5
    "00000010", --  407 - 0x197  :    2 - 0x2
    "11111111", --  408 - 0x198  :  255 - 0xff -- Sprite 0x33
    "11011111", --  409 - 0x199  :  223 - 0xdf
    "00011111", --  410 - 0x19a  :   31 - 0x1f
    "01000111", --  411 - 0x19b  :   71 - 0x47
    "01000111", --  412 - 0x19c  :   71 - 0x47
    "01000111", --  413 - 0x19d  :   71 - 0x47
    "01000111", --  414 - 0x19e  :   71 - 0x47
    "01000111", --  415 - 0x19f  :   71 - 0x47
    "01000100", --  416 - 0x1a0  :   68 - 0x44 -- Sprite 0x34
    "01000100", --  417 - 0x1a1  :   68 - 0x44
    "01000100", --  418 - 0x1a2  :   68 - 0x44
    "01000100", --  419 - 0x1a3  :   68 - 0x44
    "01000100", --  420 - 0x1a4  :   68 - 0x44
    "01000100", --  421 - 0x1a5  :   68 - 0x44
    "01000100", --  422 - 0x1a6  :   68 - 0x44
    "01000100", --  423 - 0x1a7  :   68 - 0x44
    "00010000", --  424 - 0x1a8  :   16 - 0x10 -- Sprite 0x35
    "00111000", --  425 - 0x1a9  :   56 - 0x38
    "01111100", --  426 - 0x1aa  :  124 - 0x7c
    "11111000", --  427 - 0x1ab  :  248 - 0xf8
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "01111111", --  429 - 0x1ad  :  127 - 0x7f
    "01000000", --  430 - 0x1ae  :   64 - 0x40
    "01000000", --  431 - 0x1af  :   64 - 0x40
    "00010000", --  432 - 0x1b0  :   16 - 0x10 -- Sprite 0x36
    "00111000", --  433 - 0x1b1  :   56 - 0x38
    "01111100", --  434 - 0x1b2  :  124 - 0x7c
    "11111000", --  435 - 0x1b3  :  248 - 0xf8
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "11111111", --  437 - 0x1b5  :  255 - 0xff
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "01000111", --  440 - 0x1b8  :   71 - 0x47 -- Sprite 0x37
    "01000111", --  441 - 0x1b9  :   71 - 0x47
    "01000111", --  442 - 0x1ba  :   71 - 0x47
    "01000111", --  443 - 0x1bb  :   71 - 0x47
    "01000111", --  444 - 0x1bc  :   71 - 0x47
    "11000111", --  445 - 0x1bd  :  199 - 0xc7
    "00000111", --  446 - 0x1be  :    7 - 0x7
    "00000111", --  447 - 0x1bf  :    7 - 0x7
    "01000100", --  448 - 0x1c0  :   68 - 0x44 -- Sprite 0x38
    "01000100", --  449 - 0x1c1  :   68 - 0x44
    "01000100", --  450 - 0x1c2  :   68 - 0x44
    "01000100", --  451 - 0x1c3  :   68 - 0x44
    "01000100", --  452 - 0x1c4  :   68 - 0x44
    "01011000", --  453 - 0x1c5  :   88 - 0x58
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00010000", --  456 - 0x1c8  :   16 - 0x10 -- Sprite 0x39
    "00111000", --  457 - 0x1c9  :   56 - 0x38
    "01111100", --  458 - 0x1ca  :  124 - 0x7c
    "11111000", --  459 - 0x1cb  :  248 - 0xf8
    "01110000", --  460 - 0x1cc  :  112 - 0x70
    "00100010", --  461 - 0x1cd  :   34 - 0x22
    "00000100", --  462 - 0x1ce  :    4 - 0x4
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "01000100", --  464 - 0x1d0  :   68 - 0x44 -- Sprite 0x3a
    "01000100", --  465 - 0x1d1  :   68 - 0x44
    "01000100", --  466 - 0x1d2  :   68 - 0x44
    "01000100", --  467 - 0x1d3  :   68 - 0x44
    "01000100", --  468 - 0x1d4  :   68 - 0x44
    "01011000", --  469 - 0x1d5  :   88 - 0x58
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "01000000", --  472 - 0x1d8  :   64 - 0x40 -- Sprite 0x3b
    "01000111", --  473 - 0x1d9  :   71 - 0x47
    "01000111", --  474 - 0x1da  :   71 - 0x47
    "01000111", --  475 - 0x1db  :   71 - 0x47
    "01000111", --  476 - 0x1dc  :   71 - 0x47
    "01011111", --  477 - 0x1dd  :   95 - 0x5f
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "11111111", --  481 - 0x1e1  :  255 - 0xff
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000111", --  488 - 0x1e8  :    7 - 0x7 -- Sprite 0x3d
    "11111111", --  489 - 0x1e9  :  255 - 0xff
    "11111111", --  490 - 0x1ea  :  255 - 0xff
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "11111111", --  492 - 0x1ec  :  255 - 0xff
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00010000", --  496 - 0x1f0  :   16 - 0x10 -- Sprite 0x3e
    "00111000", --  497 - 0x1f1  :   56 - 0x38
    "01110001", --  498 - 0x1f2  :  113 - 0x71
    "11100010", --  499 - 0x1f3  :  226 - 0xe2
    "01100010", --  500 - 0x1f4  :   98 - 0x62
    "00100001", --  501 - 0x1f5  :   33 - 0x21
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "10000111", --  504 - 0x1f8  :  135 - 0x87 -- Sprite 0x3f
    "10000111", --  505 - 0x1f9  :  135 - 0x87
    "00000111", --  506 - 0x1fa  :    7 - 0x7
    "00001111", --  507 - 0x1fb  :   15 - 0xf
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "00011111", --  509 - 0x1fd  :   31 - 0x1f
    "10011111", --  510 - 0x1fe  :  159 - 0x9f
    "10001111", --  511 - 0x1ff  :  143 - 0x8f
    "01000100", --  512 - 0x200  :   68 - 0x44 -- Sprite 0x40
    "01000100", --  513 - 0x201  :   68 - 0x44
    "01000100", --  514 - 0x202  :   68 - 0x44
    "01000100", --  515 - 0x203  :   68 - 0x44
    "01000100", --  516 - 0x204  :   68 - 0x44
    "01000110", --  517 - 0x205  :   70 - 0x46
    "01000110", --  518 - 0x206  :   70 - 0x46
    "01000111", --  519 - 0x207  :   71 - 0x47
    "00010000", --  520 - 0x208  :   16 - 0x10 -- Sprite 0x41
    "00111000", --  521 - 0x209  :   56 - 0x38
    "01111100", --  522 - 0x20a  :  124 - 0x7c
    "01111000", --  523 - 0x20b  :  120 - 0x78
    "00110000", --  524 - 0x20c  :   48 - 0x30
    "00000010", --  525 - 0x20d  :    2 - 0x2
    "00000101", --  526 - 0x20e  :    5 - 0x5
    "00000010", --  527 - 0x20f  :    2 - 0x2
    "00010000", --  528 - 0x210  :   16 - 0x10 -- Sprite 0x42
    "00111000", --  529 - 0x211  :   56 - 0x38
    "01111100", --  530 - 0x212  :  124 - 0x7c
    "11111000", --  531 - 0x213  :  248 - 0xf8
    "01110000", --  532 - 0x214  :  112 - 0x70
    "00100000", --  533 - 0x215  :   32 - 0x20
    "00000001", --  534 - 0x216  :    1 - 0x1
    "00000010", --  535 - 0x217  :    2 - 0x2
    "01000100", --  536 - 0x218  :   68 - 0x44 -- Sprite 0x43
    "01000100", --  537 - 0x219  :   68 - 0x44
    "01000100", --  538 - 0x21a  :   68 - 0x44
    "01000100", --  539 - 0x21b  :   68 - 0x44
    "10000100", --  540 - 0x21c  :  132 - 0x84
    "10000100", --  541 - 0x21d  :  132 - 0x84
    "00000100", --  542 - 0x21e  :    4 - 0x4
    "00001100", --  543 - 0x21f  :   12 - 0xc
    "00010000", --  544 - 0x220  :   16 - 0x10 -- Sprite 0x44
    "00111000", --  545 - 0x221  :   56 - 0x38
    "01111100", --  546 - 0x222  :  124 - 0x7c
    "11111000", --  547 - 0x223  :  248 - 0xf8
    "01110000", --  548 - 0x224  :  112 - 0x70
    "00100010", --  549 - 0x225  :   34 - 0x22
    "00000101", --  550 - 0x226  :    5 - 0x5
    "00000010", --  551 - 0x227  :    2 - 0x2
    "01001111", --  552 - 0x228  :   79 - 0x4f -- Sprite 0x45
    "01000111", --  553 - 0x229  :   71 - 0x47
    "01000111", --  554 - 0x22a  :   71 - 0x47
    "01000111", --  555 - 0x22b  :   71 - 0x47
    "01000111", --  556 - 0x22c  :   71 - 0x47
    "01000111", --  557 - 0x22d  :   71 - 0x47
    "01000111", --  558 - 0x22e  :   71 - 0x47
    "01000111", --  559 - 0x22f  :   71 - 0x47
    "10100000", --  560 - 0x230  :  160 - 0xa0 -- Sprite 0x46
    "10011111", --  561 - 0x231  :  159 - 0x9f
    "11000000", --  562 - 0x232  :  192 - 0xc0
    "11100000", --  563 - 0x233  :  224 - 0xe0
    "11111000", --  564 - 0x234  :  248 - 0xf8
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "11111111", --  567 - 0x237  :  255 - 0xff
    "00001100", --  568 - 0x238  :   12 - 0xc -- Sprite 0x47
    "11110000", --  569 - 0x239  :  240 - 0xf0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000001", --  572 - 0x23c  :    1 - 0x1
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11111111", --  574 - 0x23e  :  255 - 0xff
    "11111111", --  575 - 0x23f  :  255 - 0xff
    "00001100", --  576 - 0x240  :   12 - 0xc -- Sprite 0x48
    "00011101", --  577 - 0x241  :   29 - 0x1d
    "00111000", --  578 - 0x242  :   56 - 0x38
    "01111110", --  579 - 0x243  :  126 - 0x7e
    "11111110", --  580 - 0x244  :  254 - 0xfe
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "11111111", --  584 - 0x248  :  255 - 0xff -- Sprite 0x49
    "11111111", --  585 - 0x249  :  255 - 0xff
    "11111111", --  586 - 0x24a  :  255 - 0xff
    "11111111", --  587 - 0x24b  :  255 - 0xff
    "11111111", --  588 - 0x24c  :  255 - 0xff
    "11111111", --  589 - 0x24d  :  255 - 0xff
    "11111111", --  590 - 0x24e  :  255 - 0xff
    "11111111", --  591 - 0x24f  :  255 - 0xff
    "11111111", --  592 - 0x250  :  255 - 0xff -- Sprite 0x4a
    "11101111", --  593 - 0x251  :  239 - 0xef
    "11111101", --  594 - 0x252  :  253 - 0xfd
    "11111111", --  595 - 0x253  :  255 - 0xff
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11101111", --  597 - 0x255  :  239 - 0xef
    "11111110", --  598 - 0x256  :  254 - 0xfe
    "11111111", --  599 - 0x257  :  255 - 0xff
    "11111111", --  600 - 0x258  :  255 - 0xff -- Sprite 0x4b
    "11101010", --  601 - 0x259  :  234 - 0xea
    "11111111", --  602 - 0x25a  :  255 - 0xff
    "10101111", --  603 - 0x25b  :  175 - 0xaf
    "11111111", --  604 - 0x25c  :  255 - 0xff
    "11111111", --  605 - 0x25d  :  255 - 0xff
    "11111010", --  606 - 0x25e  :  250 - 0xfa
    "11111111", --  607 - 0x25f  :  255 - 0xff
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x4c
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111110", --  614 - 0x266  :  254 - 0xfe
    "11111111", --  615 - 0x267  :  255 - 0xff
    "11111111", --  616 - 0x268  :  255 - 0xff -- Sprite 0x4d
    "10111111", --  617 - 0x269  :  191 - 0xbf
    "11111110", --  618 - 0x26a  :  254 - 0xfe
    "10101111", --  619 - 0x26b  :  175 - 0xaf
    "11111111", --  620 - 0x26c  :  255 - 0xff
    "11111111", --  621 - 0x26d  :  255 - 0xff
    "11101111", --  622 - 0x26e  :  239 - 0xef
    "11111111", --  623 - 0x26f  :  255 - 0xff
    "11111111", --  624 - 0x270  :  255 - 0xff -- Sprite 0x4e
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11111011", --  626 - 0x272  :  251 - 0xfb
    "11111111", --  627 - 0x273  :  255 - 0xff
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111111", --  629 - 0x275  :  255 - 0xff
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11111111", --  632 - 0x278  :  255 - 0xff -- Sprite 0x4f
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11110111", --  634 - 0x27a  :  247 - 0xf7
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "11111011", --  636 - 0x27c  :  251 - 0xfb
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11101111", --  638 - 0x27e  :  239 - 0xef
    "11111101", --  639 - 0x27f  :  253 - 0xfd
    "11111111", --  640 - 0x280  :  255 - 0xff -- Sprite 0x50
    "11111111", --  641 - 0x281  :  255 - 0xff
    "00000011", --  642 - 0x282  :    3 - 0x3
    "00000001", --  643 - 0x283  :    1 - 0x1
    "11101110", --  644 - 0x284  :  238 - 0xee
    "00000000", --  645 - 0x285  :    0 - 0x0
    "11101110", --  646 - 0x286  :  238 - 0xee
    "11101110", --  647 - 0x287  :  238 - 0xee
    "11111111", --  648 - 0x288  :  255 - 0xff -- Sprite 0x51
    "11111111", --  649 - 0x289  :  255 - 0xff
    "00000011", --  650 - 0x28a  :    3 - 0x3
    "00000001", --  651 - 0x28b  :    1 - 0x1
    "11101110", --  652 - 0x28c  :  238 - 0xee
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "11101110", --  654 - 0x28e  :  238 - 0xee
    "11101110", --  655 - 0x28f  :  238 - 0xee
    "11111111", --  656 - 0x290  :  255 - 0xff -- Sprite 0x52
    "11111111", --  657 - 0x291  :  255 - 0xff
    "00000001", --  658 - 0x292  :    1 - 0x1
    "00000000", --  659 - 0x293  :    0 - 0x0
    "11100000", --  660 - 0x294  :  224 - 0xe0
    "00001111", --  661 - 0x295  :   15 - 0xf
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111011", --  663 - 0x297  :  251 - 0xfb
    "11111111", --  664 - 0x298  :  255 - 0xff -- Sprite 0x53
    "11111111", --  665 - 0x299  :  255 - 0xff
    "10000011", --  666 - 0x29a  :  131 - 0x83
    "00000001", --  667 - 0x29b  :    1 - 0x1
    "11101110", --  668 - 0x29c  :  238 - 0xee
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "11111111", --  670 - 0x29e  :  255 - 0xff
    "11111111", --  671 - 0x29f  :  255 - 0xff
    "11111111", --  672 - 0x2a0  :  255 - 0xff -- Sprite 0x54
    "11111111", --  673 - 0x2a1  :  255 - 0xff
    "00000001", --  674 - 0x2a2  :    1 - 0x1
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "10111000", --  676 - 0x2a4  :  184 - 0xb8
    "11000011", --  677 - 0x2a5  :  195 - 0xc3
    "11111011", --  678 - 0x2a6  :  251 - 0xfb
    "11111011", --  679 - 0x2a7  :  251 - 0xfb
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Sprite 0x55
    "11111111", --  681 - 0x2a9  :  255 - 0xff
    "10000011", --  682 - 0x2aa  :  131 - 0x83
    "00000001", --  683 - 0x2ab  :    1 - 0x1
    "11101110", --  684 - 0x2ac  :  238 - 0xee
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "11101110", --  686 - 0x2ae  :  238 - 0xee
    "11101110", --  687 - 0x2af  :  238 - 0xee
    "11111111", --  688 - 0x2b0  :  255 - 0xff -- Sprite 0x56
    "11111111", --  689 - 0x2b1  :  255 - 0xff
    "00011111", --  690 - 0x2b2  :   31 - 0x1f
    "00001111", --  691 - 0x2b3  :   15 - 0xf
    "11101111", --  692 - 0x2b4  :  239 - 0xef
    "00001111", --  693 - 0x2b5  :   15 - 0xf
    "11101111", --  694 - 0x2b6  :  239 - 0xef
    "11101111", --  695 - 0x2b7  :  239 - 0xef
    "11111111", --  696 - 0x2b8  :  255 - 0xff -- Sprite 0x57
    "11111111", --  697 - 0x2b9  :  255 - 0xff
    "00010001", --  698 - 0x2ba  :   17 - 0x11
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "11101110", --  700 - 0x2bc  :  238 - 0xee
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "11101110", --  702 - 0x2be  :  238 - 0xee
    "11101110", --  703 - 0x2bf  :  238 - 0xee
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Sprite 0x58
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "01110001", --  706 - 0x2c2  :  113 - 0x71
    "00110000", --  707 - 0x2c3  :   48 - 0x30
    "11111110", --  708 - 0x2c4  :  254 - 0xfe
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "11111110", --  710 - 0x2c6  :  254 - 0xfe
    "11101110", --  711 - 0x2c7  :  238 - 0xee
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- Sprite 0x59
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "00000011", --  714 - 0x2ca  :    3 - 0x3
    "00000001", --  715 - 0x2cb  :    1 - 0x1
    "11101110", --  716 - 0x2cc  :  238 - 0xee
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "11101110", --  718 - 0x2ce  :  238 - 0xee
    "11101110", --  719 - 0x2cf  :  238 - 0xee
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Sprite 0x5a
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "10000011", --  722 - 0x2d2  :  131 - 0x83
    "00000001", --  723 - 0x2d3  :    1 - 0x1
    "11101110", --  724 - 0x2d4  :  238 - 0xee
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "11101110", --  726 - 0x2d6  :  238 - 0xee
    "11101110", --  727 - 0x2d7  :  238 - 0xee
    "11111111", --  728 - 0x2d8  :  255 - 0xff -- Sprite 0x5b
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "00000001", --  730 - 0x2da  :    1 - 0x1
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "11100000", --  732 - 0x2dc  :  224 - 0xe0
    "00001111", --  733 - 0x2dd  :   15 - 0xf
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111011", --  735 - 0x2df  :  251 - 0xfb
    "11111111", --  736 - 0x2e0  :  255 - 0xff -- Sprite 0x5c
    "11111111", --  737 - 0x2e1  :  255 - 0xff
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11011101", --  743 - 0x2e7  :  221 - 0xdd
    "11111111", --  744 - 0x2e8  :  255 - 0xff -- Sprite 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "00000001", --  746 - 0x2ea  :    1 - 0x1
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "11100000", --  748 - 0x2ec  :  224 - 0xe0
    "00001111", --  749 - 0x2ed  :   15 - 0xf
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111011", --  751 - 0x2ef  :  251 - 0xfb
    "11111111", --  752 - 0x2f0  :  255 - 0xff -- Sprite 0x5e
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "00010001", --  754 - 0x2f2  :   17 - 0x11
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "11101110", --  756 - 0x2f4  :  238 - 0xee
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "11101110", --  758 - 0x2f6  :  238 - 0xee
    "11101110", --  759 - 0x2f7  :  238 - 0xee
    "10111101", --  760 - 0x2f8  :  189 - 0xbd -- Sprite 0x5f
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111111", --  763 - 0x2fb  :  255 - 0xff
    "11111111", --  764 - 0x2fc  :  255 - 0xff
    "11111111", --  765 - 0x2fd  :  255 - 0xff
    "11111111", --  766 - 0x2fe  :  255 - 0xff
    "11111111", --  767 - 0x2ff  :  255 - 0xff
    "11101110", --  768 - 0x300  :  238 - 0xee -- Sprite 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "11111110", --  770 - 0x302  :  254 - 0xfe
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000001", --  772 - 0x304  :    1 - 0x1
    "00001111", --  773 - 0x305  :   15 - 0xf
    "10001111", --  774 - 0x306  :  143 - 0x8f
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11101110", --  776 - 0x308  :  238 - 0xee -- Sprite 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "11111100", --  778 - 0x30a  :  252 - 0xfc
    "00000001", --  779 - 0x30b  :    1 - 0x1
    "00000001", --  780 - 0x30c  :    1 - 0x1
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "10001000", --  782 - 0x30e  :  136 - 0x88
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11100011", --  784 - 0x310  :  227 - 0xe3 -- Sprite 0x62
    "00001111", --  785 - 0x311  :   15 - 0xf
    "11101111", --  786 - 0x312  :  239 - 0xef
    "00001111", --  787 - 0x313  :   15 - 0xf
    "00000001", --  788 - 0x314  :    1 - 0x1
    "00000000", --  789 - 0x315  :    0 - 0x0
    "10000000", --  790 - 0x316  :  128 - 0x80
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11001110", --  792 - 0x318  :  206 - 0xce -- Sprite 0x63
    "11110000", --  793 - 0x319  :  240 - 0xf0
    "11111110", --  794 - 0x31a  :  254 - 0xfe
    "00010000", --  795 - 0x31b  :   16 - 0x10
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "10000000", --  797 - 0x31d  :  128 - 0x80
    "11000001", --  798 - 0x31e  :  193 - 0xc1
    "11111111", --  799 - 0x31f  :  255 - 0xff
    "11111011", --  800 - 0x320  :  251 - 0xfb -- Sprite 0x64
    "11000011", --  801 - 0x321  :  195 - 0xc3
    "11111011", --  802 - 0x322  :  251 - 0xfb
    "11000011", --  803 - 0x323  :  195 - 0xc3
    "11000011", --  804 - 0x324  :  195 - 0xc3
    "11000011", --  805 - 0x325  :  195 - 0xc3
    "11100011", --  806 - 0x326  :  227 - 0xe3
    "11111111", --  807 - 0x327  :  255 - 0xff
    "11101110", --  808 - 0x328  :  238 - 0xee -- Sprite 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "11111110", --  810 - 0x32a  :  254 - 0xfe
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "10001000", --  814 - 0x32e  :  136 - 0x88
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11101111", --  816 - 0x330  :  239 - 0xef -- Sprite 0x66
    "00001111", --  817 - 0x331  :   15 - 0xf
    "11101111", --  818 - 0x332  :  239 - 0xef
    "00000001", --  819 - 0x333  :    1 - 0x1
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "10000000", --  822 - 0x336  :  128 - 0x80
    "11111111", --  823 - 0x337  :  255 - 0xff
    "11101110", --  824 - 0x338  :  238 - 0xee -- Sprite 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "11111110", --  826 - 0x33a  :  254 - 0xfe
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00001000", --  829 - 0x33d  :    8 - 0x8
    "10011100", --  830 - 0x33e  :  156 - 0x9c
    "11111111", --  831 - 0x33f  :  255 - 0xff
    "11101110", --  832 - 0x340  :  238 - 0xee -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "11101110", --  834 - 0x342  :  238 - 0xee
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "10001000", --  838 - 0x346  :  136 - 0x88
    "11111111", --  839 - 0x347  :  255 - 0xff
    "11101110", --  840 - 0x348  :  238 - 0xee -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "11101110", --  842 - 0x34a  :  238 - 0xee
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "10000001", --  846 - 0x34e  :  129 - 0x81
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "11101110", --  848 - 0x350  :  238 - 0xee -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "11101110", --  850 - 0x352  :  238 - 0xee
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "10000000", --  853 - 0x355  :  128 - 0x80
    "11000001", --  854 - 0x356  :  193 - 0xc1
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11100011", --  856 - 0x358  :  227 - 0xe3 -- Sprite 0x6b
    "00001111", --  857 - 0x359  :   15 - 0xf
    "11101111", --  858 - 0x35a  :  239 - 0xef
    "00001111", --  859 - 0x35b  :   15 - 0xf
    "00000001", --  860 - 0x35c  :    1 - 0x1
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "10000000", --  862 - 0x35e  :  128 - 0x80
    "11111111", --  863 - 0x35f  :  255 - 0xff
    "10011001", --  864 - 0x360  :  153 - 0x99 -- Sprite 0x6c
    "11100011", --  865 - 0x361  :  227 - 0xe3
    "11110011", --  866 - 0x362  :  243 - 0xf3
    "11000111", --  867 - 0x363  :  199 - 0xc7
    "10000001", --  868 - 0x364  :  129 - 0x81
    "10001000", --  869 - 0x365  :  136 - 0x88
    "11001100", --  870 - 0x366  :  204 - 0xcc
    "11111111", --  871 - 0x367  :  255 - 0xff
    "11100011", --  872 - 0x368  :  227 - 0xe3 -- Sprite 0x6d
    "00001111", --  873 - 0x369  :   15 - 0xf
    "11101111", --  874 - 0x36a  :  239 - 0xef
    "00001111", --  875 - 0x36b  :   15 - 0xf
    "00001111", --  876 - 0x36c  :   15 - 0xf
    "00001111", --  877 - 0x36d  :   15 - 0xf
    "10001111", --  878 - 0x36e  :  143 - 0x8f
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11101110", --  880 - 0x370  :  238 - 0xee -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "11101110", --  882 - 0x372  :  238 - 0xee
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "10000000", --  885 - 0x375  :  128 - 0x80
    "11000001", --  886 - 0x376  :  193 - 0xc1
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff -- Sprite 0x6f
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "10111101", --  891 - 0x37b  :  189 - 0xbd
    "11111111", --  892 - 0x37c  :  255 - 0xff
    "11011011", --  893 - 0x37d  :  219 - 0xdb
    "11111111", --  894 - 0x37e  :  255 - 0xff
    "11111111", --  895 - 0x37f  :  255 - 0xff
    "11111011", --  896 - 0x380  :  251 - 0xfb -- Sprite 0x70
    "11101111", --  897 - 0x381  :  239 - 0xef
    "11011111", --  898 - 0x382  :  223 - 0xdf
    "11111111", --  899 - 0x383  :  255 - 0xff
    "10111111", --  900 - 0x384  :  191 - 0xbf
    "10111111", --  901 - 0x385  :  191 - 0xbf
    "11111110", --  902 - 0x386  :  254 - 0xfe
    "11111111", --  903 - 0x387  :  255 - 0xff
    "11011111", --  904 - 0x388  :  223 - 0xdf -- Sprite 0x71
    "11110111", --  905 - 0x389  :  247 - 0xf7
    "11111011", --  906 - 0x38a  :  251 - 0xfb
    "11111111", --  907 - 0x38b  :  255 - 0xff
    "11111101", --  908 - 0x38c  :  253 - 0xfd
    "11111101", --  909 - 0x38d  :  253 - 0xfd
    "01111111", --  910 - 0x38e  :  127 - 0x7f
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "11111111", --  912 - 0x390  :  255 - 0xff -- Sprite 0x72
    "11111111", --  913 - 0x391  :  255 - 0xff
    "11111111", --  914 - 0x392  :  255 - 0xff
    "11111111", --  915 - 0x393  :  255 - 0xff
    "11111111", --  916 - 0x394  :  255 - 0xff
    "11111111", --  917 - 0x395  :  255 - 0xff
    "11111111", --  918 - 0x396  :  255 - 0xff
    "11111111", --  919 - 0x397  :  255 - 0xff
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111110", --  921 - 0x399  :  254 - 0xfe
    "10111111", --  922 - 0x39a  :  191 - 0xbf
    "10111111", --  923 - 0x39b  :  191 - 0xbf
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11011111", --  925 - 0x39d  :  223 - 0xdf
    "11101111", --  926 - 0x39e  :  239 - 0xef
    "11111011", --  927 - 0x39f  :  251 - 0xfb
    "11111111", --  928 - 0x3a0  :  255 - 0xff -- Sprite 0x74
    "01111111", --  929 - 0x3a1  :  127 - 0x7f
    "11111101", --  930 - 0x3a2  :  253 - 0xfd
    "11111101", --  931 - 0x3a3  :  253 - 0xfd
    "11111111", --  932 - 0x3a4  :  255 - 0xff
    "11111011", --  933 - 0x3a5  :  251 - 0xfb
    "11110111", --  934 - 0x3a6  :  247 - 0xf7
    "11011111", --  935 - 0x3a7  :  223 - 0xdf
    "11111111", --  936 - 0x3a8  :  255 - 0xff -- Sprite 0x75
    "11111111", --  937 - 0x3a9  :  255 - 0xff
    "11111111", --  938 - 0x3aa  :  255 - 0xff
    "11111111", --  939 - 0x3ab  :  255 - 0xff
    "11111111", --  940 - 0x3ac  :  255 - 0xff
    "11111111", --  941 - 0x3ad  :  255 - 0xff
    "11111111", --  942 - 0x3ae  :  255 - 0xff
    "11111111", --  943 - 0x3af  :  255 - 0xff
    "11111111", --  944 - 0x3b0  :  255 - 0xff -- Sprite 0x76
    "11111111", --  945 - 0x3b1  :  255 - 0xff
    "11111111", --  946 - 0x3b2  :  255 - 0xff
    "11111111", --  947 - 0x3b3  :  255 - 0xff
    "11111111", --  948 - 0x3b4  :  255 - 0xff
    "11111111", --  949 - 0x3b5  :  255 - 0xff
    "11111111", --  950 - 0x3b6  :  255 - 0xff
    "11111111", --  951 - 0x3b7  :  255 - 0xff
    "11111111", --  952 - 0x3b8  :  255 - 0xff -- Sprite 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111111", --  954 - 0x3ba  :  255 - 0xff
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "11111111", --  956 - 0x3bc  :  255 - 0xff
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Sprite 0x78
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "11111111", --  966 - 0x3c6  :  255 - 0xff
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Sprite 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "11111111", --  971 - 0x3cb  :  255 - 0xff
    "11111111", --  972 - 0x3cc  :  255 - 0xff
    "11111111", --  973 - 0x3cd  :  255 - 0xff
    "11111111", --  974 - 0x3ce  :  255 - 0xff
    "11111111", --  975 - 0x3cf  :  255 - 0xff
    "11111111", --  976 - 0x3d0  :  255 - 0xff -- Sprite 0x7a
    "11111111", --  977 - 0x3d1  :  255 - 0xff
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "11111111", --  980 - 0x3d4  :  255 - 0xff
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "11111111", --  982 - 0x3d6  :  255 - 0xff
    "11111111", --  983 - 0x3d7  :  255 - 0xff
    "11111111", --  984 - 0x3d8  :  255 - 0xff -- Sprite 0x7b
    "11111111", --  985 - 0x3d9  :  255 - 0xff
    "11111111", --  986 - 0x3da  :  255 - 0xff
    "11111111", --  987 - 0x3db  :  255 - 0xff
    "11111111", --  988 - 0x3dc  :  255 - 0xff
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "11111111", --  991 - 0x3df  :  255 - 0xff
    "11111111", --  992 - 0x3e0  :  255 - 0xff -- Sprite 0x7c
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111111", --  996 - 0x3e4  :  255 - 0xff
    "11111111", --  997 - 0x3e5  :  255 - 0xff
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "11111111", -- 1000 - 0x3e8  :  255 - 0xff -- Sprite 0x7d
    "11111111", -- 1001 - 0x3e9  :  255 - 0xff
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111111", -- 1004 - 0x3ec  :  255 - 0xff
    "11111111", -- 1005 - 0x3ed  :  255 - 0xff
    "11111111", -- 1006 - 0x3ee  :  255 - 0xff
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "11111111", -- 1008 - 0x3f0  :  255 - 0xff -- Sprite 0x7e
    "11111111", -- 1009 - 0x3f1  :  255 - 0xff
    "11111111", -- 1010 - 0x3f2  :  255 - 0xff
    "11111111", -- 1011 - 0x3f3  :  255 - 0xff
    "11111111", -- 1012 - 0x3f4  :  255 - 0xff
    "11111111", -- 1013 - 0x3f5  :  255 - 0xff
    "11111111", -- 1014 - 0x3f6  :  255 - 0xff
    "11111111", -- 1015 - 0x3f7  :  255 - 0xff
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Sprite 0x7f
    "11111111", -- 1017 - 0x3f9  :  255 - 0xff
    "11111111", -- 1018 - 0x3fa  :  255 - 0xff
    "11111111", -- 1019 - 0x3fb  :  255 - 0xff
    "11111111", -- 1020 - 0x3fc  :  255 - 0xff
    "11111111", -- 1021 - 0x3fd  :  255 - 0xff
    "11111111", -- 1022 - 0x3fe  :  255 - 0xff
    "11111111", -- 1023 - 0x3ff  :  255 - 0xff
    "10111111", -- 1024 - 0x400  :  191 - 0xbf -- Sprite 0x80
    "11110111", -- 1025 - 0x401  :  247 - 0xf7
    "11111101", -- 1026 - 0x402  :  253 - 0xfd
    "11011111", -- 1027 - 0x403  :  223 - 0xdf
    "11111011", -- 1028 - 0x404  :  251 - 0xfb
    "10111111", -- 1029 - 0x405  :  191 - 0xbf
    "11111110", -- 1030 - 0x406  :  254 - 0xfe
    "11101111", -- 1031 - 0x407  :  239 - 0xef
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Sprite 0x81
    "11101110", -- 1033 - 0x409  :  238 - 0xee
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11011111", -- 1035 - 0x40b  :  223 - 0xdf
    "01110111", -- 1036 - 0x40c  :  119 - 0x77
    "11111101", -- 1037 - 0x40d  :  253 - 0xfd
    "11011111", -- 1038 - 0x40e  :  223 - 0xdf
    "10111111", -- 1039 - 0x40f  :  191 - 0xbf
    "11111110", -- 1040 - 0x410  :  254 - 0xfe -- Sprite 0x82
    "11101111", -- 1041 - 0x411  :  239 - 0xef
    "10111111", -- 1042 - 0x412  :  191 - 0xbf
    "11110111", -- 1043 - 0x413  :  247 - 0xf7
    "11111101", -- 1044 - 0x414  :  253 - 0xfd
    "11011111", -- 1045 - 0x415  :  223 - 0xdf
    "11111011", -- 1046 - 0x416  :  251 - 0xfb
    "10111111", -- 1047 - 0x417  :  191 - 0xbf
    "11101111", -- 1048 - 0x418  :  239 - 0xef -- Sprite 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "10111011", -- 1050 - 0x41a  :  187 - 0xbb
    "11111111", -- 1051 - 0x41b  :  255 - 0xff
    "11110111", -- 1052 - 0x41c  :  247 - 0xf7
    "11011101", -- 1053 - 0x41d  :  221 - 0xdd
    "01111111", -- 1054 - 0x41e  :  127 - 0x7f
    "11110111", -- 1055 - 0x41f  :  247 - 0xf7
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Sprite 0x84
    "11101110", -- 1057 - 0x421  :  238 - 0xee
    "11111011", -- 1058 - 0x422  :  251 - 0xfb
    "10111111", -- 1059 - 0x423  :  191 - 0xbf
    "01111111", -- 1060 - 0x424  :  127 - 0x7f
    "11101101", -- 1061 - 0x425  :  237 - 0xed
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "10111111", -- 1063 - 0x427  :  191 - 0xbf
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "10111111", -- 1065 - 0x429  :  191 - 0xbf
    "01111101", -- 1066 - 0x42a  :  125 - 0x7d
    "11110111", -- 1067 - 0x42b  :  247 - 0xf7
    "11011011", -- 1068 - 0x42c  :  219 - 0xdb
    "11111101", -- 1069 - 0x42d  :  253 - 0xfd
    "01111110", -- 1070 - 0x42e  :  126 - 0x7e
    "11111011", -- 1071 - 0x42f  :  251 - 0xfb
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Sprite 0x86
    "11110111", -- 1073 - 0x431  :  247 - 0xf7
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11011101", -- 1075 - 0x433  :  221 - 0xdd
    "01111111", -- 1076 - 0x434  :  127 - 0x7f
    "11110111", -- 1077 - 0x435  :  247 - 0xf7
    "11101111", -- 1078 - 0x436  :  239 - 0xef
    "10111101", -- 1079 - 0x437  :  189 - 0xbd
    "01011111", -- 1080 - 0x438  :   95 - 0x5f -- Sprite 0x87
    "11111101", -- 1081 - 0x439  :  253 - 0xfd
    "11110110", -- 1082 - 0x43a  :  246 - 0xf6
    "01111111", -- 1083 - 0x43b  :  127 - 0x7f
    "10011111", -- 1084 - 0x43c  :  159 - 0x9f
    "11111110", -- 1085 - 0x43d  :  254 - 0xfe
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "11101111", -- 1087 - 0x43f  :  239 - 0xef
    "11111111", -- 1088 - 0x440  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "10011111", -- 1090 - 0x442  :  159 - 0x9f
    "10110011", -- 1091 - 0x443  :  179 - 0xb3
    "11110011", -- 1092 - 0x444  :  243 - 0xf3
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- Sprite 0x89
    "11001111", -- 1097 - 0x449  :  207 - 0xcf
    "11011111", -- 1098 - 0x44a  :  223 - 0xdf
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11110011", -- 1100 - 0x44c  :  243 - 0xf3
    "11110011", -- 1101 - 0x44d  :  243 - 0xf3
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "10111111", -- 1104 - 0x450  :  191 - 0xbf -- Sprite 0x8a
    "11110111", -- 1105 - 0x451  :  247 - 0xf7
    "11111101", -- 1106 - 0x452  :  253 - 0xfd
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "11111011", -- 1108 - 0x454  :  251 - 0xfb
    "10111111", -- 1109 - 0x455  :  191 - 0xbf
    "11111110", -- 1110 - 0x456  :  254 - 0xfe
    "11101111", -- 1111 - 0x457  :  239 - 0xef
    "10111111", -- 1112 - 0x458  :  191 - 0xbf -- Sprite 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11101110", -- 1114 - 0x45a  :  238 - 0xee
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11011111", -- 1116 - 0x45c  :  223 - 0xdf
    "01111101", -- 1117 - 0x45d  :  125 - 0x7d
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11011111", -- 1119 - 0x45f  :  223 - 0xdf
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Sprite 0x8c
    "11111000", -- 1121 - 0x461  :  248 - 0xf8
    "11100010", -- 1122 - 0x462  :  226 - 0xe2
    "11010111", -- 1123 - 0x463  :  215 - 0xd7
    "11001111", -- 1124 - 0x464  :  207 - 0xcf
    "10011111", -- 1125 - 0x465  :  159 - 0x9f
    "10111110", -- 1126 - 0x466  :  190 - 0xbe
    "10011101", -- 1127 - 0x467  :  157 - 0x9d
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- Sprite 0x8d
    "00011111", -- 1129 - 0x469  :   31 - 0x1f
    "10100111", -- 1130 - 0x46a  :  167 - 0xa7
    "11000011", -- 1131 - 0x46b  :  195 - 0xc3
    "11100011", -- 1132 - 0x46c  :  227 - 0xe3
    "01000001", -- 1133 - 0x46d  :   65 - 0x41
    "10100001", -- 1134 - 0x46e  :  161 - 0xa1
    "00000001", -- 1135 - 0x46f  :    1 - 0x1
    "10111110", -- 1136 - 0x470  :  190 - 0xbe -- Sprite 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11011111", -- 1138 - 0x472  :  223 - 0xdf
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11101111", -- 1140 - 0x474  :  239 - 0xef
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11110111", -- 1142 - 0x476  :  247 - 0xf7
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "01111101", -- 1144 - 0x478  :  125 - 0x7d -- Sprite 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111011", -- 1146 - 0x47a  :  251 - 0xfb
    "11111111", -- 1147 - 0x47b  :  255 - 0xff
    "11110111", -- 1148 - 0x47c  :  247 - 0xf7
    "11111111", -- 1149 - 0x47d  :  255 - 0xff
    "11101111", -- 1150 - 0x47e  :  239 - 0xef
    "11111111", -- 1151 - 0x47f  :  255 - 0xff
    "10111110", -- 1152 - 0x480  :  190 - 0xbe -- Sprite 0x90
    "11110111", -- 1153 - 0x481  :  247 - 0xf7
    "11111111", -- 1154 - 0x482  :  255 - 0xff
    "11011111", -- 1155 - 0x483  :  223 - 0xdf
    "11111011", -- 1156 - 0x484  :  251 - 0xfb
    "11111110", -- 1157 - 0x485  :  254 - 0xfe
    "10111111", -- 1158 - 0x486  :  191 - 0xbf
    "11110111", -- 1159 - 0x487  :  247 - 0xf7
    "11101110", -- 1160 - 0x488  :  238 - 0xee -- Sprite 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "01111011", -- 1162 - 0x48a  :  123 - 0x7b
    "11111101", -- 1163 - 0x48b  :  253 - 0xfd
    "11101111", -- 1164 - 0x48c  :  239 - 0xef
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "10111101", -- 1166 - 0x48e  :  189 - 0xbd
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11111011", -- 1168 - 0x490  :  251 - 0xfb -- Sprite 0x92
    "10111111", -- 1169 - 0x491  :  191 - 0xbf
    "11101111", -- 1170 - 0x492  :  239 - 0xef
    "11111101", -- 1171 - 0x493  :  253 - 0xfd
    "11111111", -- 1172 - 0x494  :  255 - 0xff
    "10111111", -- 1173 - 0x495  :  191 - 0xbf
    "11111011", -- 1174 - 0x496  :  251 - 0xfb
    "11011111", -- 1175 - 0x497  :  223 - 0xdf
    "10111101", -- 1176 - 0x498  :  189 - 0xbd -- Sprite 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "01110111", -- 1178 - 0x49a  :  119 - 0x77
    "11111110", -- 1179 - 0x49b  :  254 - 0xfe
    "11011111", -- 1180 - 0x49c  :  223 - 0xdf
    "11111011", -- 1181 - 0x49d  :  251 - 0xfb
    "11101111", -- 1182 - 0x49e  :  239 - 0xef
    "01111111", -- 1183 - 0x49f  :  127 - 0x7f
    "01111111", -- 1184 - 0x4a0  :  127 - 0x7f -- Sprite 0x94
    "11110111", -- 1185 - 0x4a1  :  247 - 0xf7
    "11011101", -- 1186 - 0x4a2  :  221 - 0xdd
    "01111011", -- 1187 - 0x4a3  :  123 - 0x7b
    "11111111", -- 1188 - 0x4a4  :  255 - 0xff
    "11101110", -- 1189 - 0x4a5  :  238 - 0xee
    "10111011", -- 1190 - 0x4a6  :  187 - 0xbb
    "11111101", -- 1191 - 0x4a7  :  253 - 0xfd
    "11010111", -- 1192 - 0x4a8  :  215 - 0xd7 -- Sprite 0x95
    "01111111", -- 1193 - 0x4a9  :  127 - 0x7f
    "11111101", -- 1194 - 0x4aa  :  253 - 0xfd
    "11101110", -- 1195 - 0x4ab  :  238 - 0xee
    "11110111", -- 1196 - 0x4ac  :  247 - 0xf7
    "10111011", -- 1197 - 0x4ad  :  187 - 0xbb
    "11101111", -- 1198 - 0x4ae  :  239 - 0xef
    "11110111", -- 1199 - 0x4af  :  247 - 0xf7
    "10111111", -- 1200 - 0x4b0  :  191 - 0xbf -- Sprite 0x96
    "11101110", -- 1201 - 0x4b1  :  238 - 0xee
    "11011011", -- 1202 - 0x4b2  :  219 - 0xdb
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "01110111", -- 1204 - 0x4b4  :  119 - 0x77
    "11011101", -- 1205 - 0x4b5  :  221 - 0xdd
    "11101111", -- 1206 - 0x4b6  :  239 - 0xef
    "11111011", -- 1207 - 0x4b7  :  251 - 0xfb
    "11111101", -- 1208 - 0x4b8  :  253 - 0xfd -- Sprite 0x97
    "11101110", -- 1209 - 0x4b9  :  238 - 0xee
    "11111011", -- 1210 - 0x4ba  :  251 - 0xfb
    "11111101", -- 1211 - 0x4bb  :  253 - 0xfd
    "11110101", -- 1212 - 0x4bc  :  245 - 0xf5
    "11011111", -- 1213 - 0x4bd  :  223 - 0xdf
    "01111111", -- 1214 - 0x4be  :  127 - 0x7f
    "10111011", -- 1215 - 0x4bf  :  187 - 0xbb
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x98
    "11001111", -- 1217 - 0x4c1  :  207 - 0xcf
    "11011111", -- 1218 - 0x4c2  :  223 - 0xdf
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11110011", -- 1220 - 0x4c4  :  243 - 0xf3
    "11110011", -- 1221 - 0x4c5  :  243 - 0xf3
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "10011111", -- 1226 - 0x4ca  :  159 - 0x9f
    "10110011", -- 1227 - 0x4cb  :  179 - 0xb3
    "11110011", -- 1228 - 0x4cc  :  243 - 0xf3
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "10111111", -- 1232 - 0x4d0  :  191 - 0xbf -- Sprite 0x9a
    "11110111", -- 1233 - 0x4d1  :  247 - 0xf7
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11011111", -- 1235 - 0x4d3  :  223 - 0xdf
    "11111011", -- 1236 - 0x4d4  :  251 - 0xfb
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "10111111", -- 1238 - 0x4d6  :  191 - 0xbf
    "11110111", -- 1239 - 0x4d7  :  247 - 0xf7
    "11011111", -- 1240 - 0x4d8  :  223 - 0xdf -- Sprite 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "01111011", -- 1242 - 0x4da  :  123 - 0x7b
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11101111", -- 1244 - 0x4dc  :  239 - 0xef
    "11111101", -- 1245 - 0x4dd  :  253 - 0xfd
    "10111111", -- 1246 - 0x4de  :  191 - 0xbf
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "10111010", -- 1248 - 0x4e0  :  186 - 0xba -- Sprite 0x9c
    "10011100", -- 1249 - 0x4e1  :  156 - 0x9c
    "10101010", -- 1250 - 0x4e2  :  170 - 0xaa
    "11000000", -- 1251 - 0x4e3  :  192 - 0xc0
    "11000000", -- 1252 - 0x4e4  :  192 - 0xc0
    "11100000", -- 1253 - 0x4e5  :  224 - 0xe0
    "11111000", -- 1254 - 0x4e6  :  248 - 0xf8
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000001", -- 1256 - 0x4e8  :    1 - 0x1 -- Sprite 0x9d
    "00000001", -- 1257 - 0x4e9  :    1 - 0x1
    "00000001", -- 1258 - 0x4ea  :    1 - 0x1
    "00000011", -- 1259 - 0x4eb  :    3 - 0x3
    "00000011", -- 1260 - 0x4ec  :    3 - 0x3
    "00000111", -- 1261 - 0x4ed  :    7 - 0x7
    "00011111", -- 1262 - 0x4ee  :   31 - 0x1f
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "01111101", -- 1264 - 0x4f0  :  125 - 0x7d -- Sprite 0x9e
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11111011", -- 1266 - 0x4f2  :  251 - 0xfb
    "11111111", -- 1267 - 0x4f3  :  255 - 0xff
    "11111111", -- 1268 - 0x4f4  :  255 - 0xff
    "11111011", -- 1269 - 0x4f5  :  251 - 0xfb
    "11111111", -- 1270 - 0x4f6  :  255 - 0xff
    "01111101", -- 1271 - 0x4f7  :  125 - 0x7d
    "11111111", -- 1272 - 0x4f8  :  255 - 0xff -- Sprite 0x9f
    "11111111", -- 1273 - 0x4f9  :  255 - 0xff
    "10111101", -- 1274 - 0x4fa  :  189 - 0xbd
    "11111111", -- 1275 - 0x4fb  :  255 - 0xff
    "11111111", -- 1276 - 0x4fc  :  255 - 0xff
    "11111111", -- 1277 - 0x4fd  :  255 - 0xff
    "11111111", -- 1278 - 0x4fe  :  255 - 0xff
    "10111101", -- 1279 - 0x4ff  :  189 - 0xbd
    "11101111", -- 1280 - 0x500  :  239 - 0xef -- Sprite 0xa0
    "11000111", -- 1281 - 0x501  :  199 - 0xc7
    "10000011", -- 1282 - 0x502  :  131 - 0x83
    "00000111", -- 1283 - 0x503  :    7 - 0x7
    "10001111", -- 1284 - 0x504  :  143 - 0x8f
    "11011101", -- 1285 - 0x505  :  221 - 0xdd
    "11111010", -- 1286 - 0x506  :  250 - 0xfa
    "11111101", -- 1287 - 0x507  :  253 - 0xfd
    "11101111", -- 1288 - 0x508  :  239 - 0xef -- Sprite 0xa1
    "11000111", -- 1289 - 0x509  :  199 - 0xc7
    "10000011", -- 1290 - 0x50a  :  131 - 0x83
    "00011111", -- 1291 - 0x50b  :   31 - 0x1f
    "10010000", -- 1292 - 0x50c  :  144 - 0x90
    "11010100", -- 1293 - 0x50d  :  212 - 0xd4
    "11110011", -- 1294 - 0x50e  :  243 - 0xf3
    "11110010", -- 1295 - 0x50f  :  242 - 0xf2
    "11101111", -- 1296 - 0x510  :  239 - 0xef -- Sprite 0xa2
    "11000111", -- 1297 - 0x511  :  199 - 0xc7
    "10000011", -- 1298 - 0x512  :  131 - 0x83
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "01010101", -- 1302 - 0x516  :   85 - 0x55
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "11110000", -- 1304 - 0x518  :  240 - 0xf0 -- Sprite 0xa3
    "11010010", -- 1305 - 0x519  :  210 - 0xd2
    "10010000", -- 1306 - 0x51a  :  144 - 0x90
    "00010010", -- 1307 - 0x51b  :   18 - 0x12
    "10010000", -- 1308 - 0x51c  :  144 - 0x90
    "11010010", -- 1309 - 0x51d  :  210 - 0xd2
    "11110000", -- 1310 - 0x51e  :  240 - 0xf0
    "11110010", -- 1311 - 0x51f  :  242 - 0xf2
    "11110000", -- 1312 - 0x520  :  240 - 0xf0 -- Sprite 0xa4
    "11010011", -- 1313 - 0x521  :  211 - 0xd3
    "10010100", -- 1314 - 0x522  :  148 - 0x94
    "00011000", -- 1315 - 0x523  :   24 - 0x18
    "10011111", -- 1316 - 0x524  :  159 - 0x9f
    "11011101", -- 1317 - 0x525  :  221 - 0xdd
    "11111010", -- 1318 - 0x526  :  250 - 0xfa
    "11111101", -- 1319 - 0x527  :  253 - 0xfd
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11011101", -- 1325 - 0x52d  :  221 - 0xdd
    "11111010", -- 1326 - 0x52e  :  250 - 0xfa
    "11111101", -- 1327 - 0x52f  :  253 - 0xfd
    "11101111", -- 1328 - 0x530  :  239 - 0xef -- Sprite 0xa6
    "11000111", -- 1329 - 0x531  :  199 - 0xc7
    "10000011", -- 1330 - 0x532  :  131 - 0x83
    "11111111", -- 1331 - 0x533  :  255 - 0xff
    "00011111", -- 1332 - 0x534  :   31 - 0x1f
    "00101101", -- 1333 - 0x535  :   45 - 0x2d
    "01001010", -- 1334 - 0x536  :   74 - 0x4a
    "01001101", -- 1335 - 0x537  :   77 - 0x4d
    "01001111", -- 1336 - 0x538  :   79 - 0x4f -- Sprite 0xa7
    "01001111", -- 1337 - 0x539  :   79 - 0x4f
    "01001011", -- 1338 - 0x53a  :   75 - 0x4b
    "01001111", -- 1339 - 0x53b  :   79 - 0x4f
    "01001111", -- 1340 - 0x53c  :   79 - 0x4f
    "01001101", -- 1341 - 0x53d  :   77 - 0x4d
    "01001010", -- 1342 - 0x53e  :   74 - 0x4a
    "01001101", -- 1343 - 0x53f  :   77 - 0x4d
    "01001111", -- 1344 - 0x540  :   79 - 0x4f -- Sprite 0xa8
    "11001111", -- 1345 - 0x541  :  207 - 0xcf
    "00001011", -- 1346 - 0x542  :   11 - 0xb
    "00001111", -- 1347 - 0x543  :   15 - 0xf
    "11111111", -- 1348 - 0x544  :  255 - 0xff
    "11011101", -- 1349 - 0x545  :  221 - 0xdd
    "11111010", -- 1350 - 0x546  :  250 - 0xfa
    "11111101", -- 1351 - 0x547  :  253 - 0xfd
    "11111111", -- 1352 - 0x548  :  255 - 0xff -- Sprite 0xa9
    "11111111", -- 1353 - 0x549  :  255 - 0xff
    "11111111", -- 1354 - 0x54a  :  255 - 0xff
    "11111111", -- 1355 - 0x54b  :  255 - 0xff
    "11111111", -- 1356 - 0x54c  :  255 - 0xff
    "11111111", -- 1357 - 0x54d  :  255 - 0xff
    "11111111", -- 1358 - 0x54e  :  255 - 0xff
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Sprite 0xaa
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "10101111", -- 1362 - 0x552  :  175 - 0xaf
    "01010111", -- 1363 - 0x553  :   87 - 0x57
    "10001111", -- 1364 - 0x554  :  143 - 0x8f
    "11011101", -- 1365 - 0x555  :  221 - 0xdd
    "11111010", -- 1366 - 0x556  :  250 - 0xfa
    "11111101", -- 1367 - 0x557  :  253 - 0xfd
    "11111111", -- 1368 - 0x558  :  255 - 0xff -- Sprite 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Sprite 0xad
    "11111111", -- 1385 - 0x569  :  255 - 0xff
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "11111111", -- 1388 - 0x56c  :  255 - 0xff
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Sprite 0xae
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "11111111", -- 1394 - 0x572  :  255 - 0xff
    "11111111", -- 1395 - 0x573  :  255 - 0xff
    "11111111", -- 1396 - 0x574  :  255 - 0xff
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "11111111", -- 1398 - 0x576  :  255 - 0xff
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "11111111", -- 1400 - 0x578  :  255 - 0xff -- Sprite 0xaf
    "11111111", -- 1401 - 0x579  :  255 - 0xff
    "11111111", -- 1402 - 0x57a  :  255 - 0xff
    "11111111", -- 1403 - 0x57b  :  255 - 0xff
    "11111111", -- 1404 - 0x57c  :  255 - 0xff
    "11111111", -- 1405 - 0x57d  :  255 - 0xff
    "11111111", -- 1406 - 0x57e  :  255 - 0xff
    "11111111", -- 1407 - 0x57f  :  255 - 0xff
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00011111", -- 1409 - 0x581  :   31 - 0x1f
    "00010000", -- 1410 - 0x582  :   16 - 0x10
    "00010000", -- 1411 - 0x583  :   16 - 0x10
    "00010000", -- 1412 - 0x584  :   16 - 0x10
    "00010000", -- 1413 - 0x585  :   16 - 0x10
    "00010000", -- 1414 - 0x586  :   16 - 0x10
    "00010000", -- 1415 - 0x587  :   16 - 0x10
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- Sprite 0xb1
    "11111000", -- 1417 - 0x589  :  248 - 0xf8
    "00001000", -- 1418 - 0x58a  :    8 - 0x8
    "00001000", -- 1419 - 0x58b  :    8 - 0x8
    "00001000", -- 1420 - 0x58c  :    8 - 0x8
    "00001000", -- 1421 - 0x58d  :    8 - 0x8
    "00001000", -- 1422 - 0x58e  :    8 - 0x8
    "00001000", -- 1423 - 0x58f  :    8 - 0x8
    "00010000", -- 1424 - 0x590  :   16 - 0x10 -- Sprite 0xb2
    "00010000", -- 1425 - 0x591  :   16 - 0x10
    "00010000", -- 1426 - 0x592  :   16 - 0x10
    "00010000", -- 1427 - 0x593  :   16 - 0x10
    "00011111", -- 1428 - 0x594  :   31 - 0x1f
    "00011111", -- 1429 - 0x595  :   31 - 0x1f
    "00001111", -- 1430 - 0x596  :   15 - 0xf
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00001000", -- 1432 - 0x598  :    8 - 0x8 -- Sprite 0xb3
    "00001000", -- 1433 - 0x599  :    8 - 0x8
    "00001000", -- 1434 - 0x59a  :    8 - 0x8
    "00001000", -- 1435 - 0x59b  :    8 - 0x8
    "11111000", -- 1436 - 0x59c  :  248 - 0xf8
    "11111000", -- 1437 - 0x59d  :  248 - 0xf8
    "11110000", -- 1438 - 0x59e  :  240 - 0xf0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00111111", -- 1442 - 0x5a2  :   63 - 0x3f
    "01100000", -- 1443 - 0x5a3  :   96 - 0x60
    "01100000", -- 1444 - 0x5a4  :   96 - 0x60
    "01100000", -- 1445 - 0x5a5  :   96 - 0x60
    "01100000", -- 1446 - 0x5a6  :   96 - 0x60
    "01100000", -- 1447 - 0x5a7  :   96 - 0x60
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- Sprite 0xb5
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "11111100", -- 1450 - 0x5aa  :  252 - 0xfc
    "00000110", -- 1451 - 0x5ab  :    6 - 0x6
    "00000110", -- 1452 - 0x5ac  :    6 - 0x6
    "00000110", -- 1453 - 0x5ad  :    6 - 0x6
    "00000110", -- 1454 - 0x5ae  :    6 - 0x6
    "00000110", -- 1455 - 0x5af  :    6 - 0x6
    "01100000", -- 1456 - 0x5b0  :   96 - 0x60 -- Sprite 0xb6
    "01100000", -- 1457 - 0x5b1  :   96 - 0x60
    "01100000", -- 1458 - 0x5b2  :   96 - 0x60
    "01111111", -- 1459 - 0x5b3  :  127 - 0x7f
    "01111111", -- 1460 - 0x5b4  :  127 - 0x7f
    "00111111", -- 1461 - 0x5b5  :   63 - 0x3f
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000110", -- 1464 - 0x5b8  :    6 - 0x6 -- Sprite 0xb7
    "00000110", -- 1465 - 0x5b9  :    6 - 0x6
    "00000110", -- 1466 - 0x5ba  :    6 - 0x6
    "11111110", -- 1467 - 0x5bb  :  254 - 0xfe
    "11111110", -- 1468 - 0x5bc  :  254 - 0xfe
    "11111100", -- 1469 - 0x5bd  :  252 - 0xfc
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "01100000", -- 1472 - 0x5c0  :   96 - 0x60 -- Sprite 0xb8
    "11110011", -- 1473 - 0x5c1  :  243 - 0xf3
    "11000111", -- 1474 - 0x5c2  :  199 - 0xc7
    "10000110", -- 1475 - 0x5c3  :  134 - 0x86
    "00000100", -- 1476 - 0x5c4  :    4 - 0x4
    "00000100", -- 1477 - 0x5c5  :    4 - 0x4
    "00000111", -- 1478 - 0x5c6  :    7 - 0x7
    "00000111", -- 1479 - 0x5c7  :    7 - 0x7
    "00000110", -- 1480 - 0x5c8  :    6 - 0x6 -- Sprite 0xb9
    "10001111", -- 1481 - 0x5c9  :  143 - 0x8f
    "11000101", -- 1482 - 0x5ca  :  197 - 0xc5
    "00100011", -- 1483 - 0x5cb  :   35 - 0x23
    "00101110", -- 1484 - 0x5cc  :   46 - 0x2e
    "01100000", -- 1485 - 0x5cd  :   96 - 0x60
    "11100001", -- 1486 - 0x5ce  :  225 - 0xe1
    "11100001", -- 1487 - 0x5cf  :  225 - 0xe1
    "11001000", -- 1488 - 0x5d0  :  200 - 0xc8 -- Sprite 0xba
    "11111000", -- 1489 - 0x5d1  :  248 - 0xf8
    "10110000", -- 1490 - 0x5d2  :  176 - 0xb0
    "00010000", -- 1491 - 0x5d3  :   16 - 0x10
    "00110000", -- 1492 - 0x5d4  :   48 - 0x30
    "11001000", -- 1493 - 0x5d5  :  200 - 0xc8
    "11111000", -- 1494 - 0x5d6  :  248 - 0xf8
    "10000000", -- 1495 - 0x5d7  :  128 - 0x80
    "00000011", -- 1496 - 0x5d8  :    3 - 0x3 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "01100000", -- 1499 - 0x5db  :   96 - 0x60
    "11110000", -- 1500 - 0x5dc  :  240 - 0xf0
    "11010000", -- 1501 - 0x5dd  :  208 - 0xd0
    "10010000", -- 1502 - 0x5de  :  144 - 0x90
    "01100000", -- 1503 - 0x5df  :   96 - 0x60
    "11000011", -- 1504 - 0x5e0  :  195 - 0xc3 -- Sprite 0xbc
    "00001110", -- 1505 - 0x5e1  :   14 - 0xe
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000110", -- 1507 - 0x5e3  :    6 - 0x6
    "00001111", -- 1508 - 0x5e4  :   15 - 0xf
    "00001101", -- 1509 - 0x5e5  :   13 - 0xd
    "00001001", -- 1510 - 0x5e6  :    9 - 0x9
    "00000110", -- 1511 - 0x5e7  :    6 - 0x6
    "11100000", -- 1512 - 0x5e8  :  224 - 0xe0 -- Sprite 0xbd
    "01100011", -- 1513 - 0x5e9  :   99 - 0x63
    "11100111", -- 1514 - 0x5ea  :  231 - 0xe7
    "11100110", -- 1515 - 0x5eb  :  230 - 0xe6
    "00000100", -- 1516 - 0x5ec  :    4 - 0x4
    "00000100", -- 1517 - 0x5ed  :    4 - 0x4
    "00000111", -- 1518 - 0x5ee  :    7 - 0x7
    "00000111", -- 1519 - 0x5ef  :    7 - 0x7
    "00000111", -- 1520 - 0x5f0  :    7 - 0x7 -- Sprite 0xbe
    "10000011", -- 1521 - 0x5f1  :  131 - 0x83
    "11000111", -- 1522 - 0x5f2  :  199 - 0xc7
    "00100111", -- 1523 - 0x5f3  :   39 - 0x27
    "00100000", -- 1524 - 0x5f4  :   32 - 0x20
    "01100000", -- 1525 - 0x5f5  :   96 - 0x60
    "11100000", -- 1526 - 0x5f6  :  224 - 0xe0
    "11100000", -- 1527 - 0x5f7  :  224 - 0xe0
    "00000011", -- 1528 - 0x5f8  :    3 - 0x3 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00001100", -- 1530 - 0x5fa  :   12 - 0xc
    "00001100", -- 1531 - 0x5fb  :   12 - 0xc
    "11100100", -- 1532 - 0x5fc  :  228 - 0xe4
    "01101100", -- 1533 - 0x5fd  :  108 - 0x6c
    "11101101", -- 1534 - 0x5fe  :  237 - 0xed
    "11100111", -- 1535 - 0x5ff  :  231 - 0xe7
    "11000000", -- 1536 - 0x600  :  192 - 0xc0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00110000", -- 1538 - 0x602  :   48 - 0x30
    "00110000", -- 1539 - 0x603  :   48 - 0x30
    "00010111", -- 1540 - 0x604  :   23 - 0x17
    "00110011", -- 1541 - 0x605  :   51 - 0x33
    "01110111", -- 1542 - 0x606  :  119 - 0x77
    "11010111", -- 1543 - 0x607  :  215 - 0xd7
    "00001100", -- 1544 - 0x608  :   12 - 0xc -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00110000", -- 1552 - 0x610  :   48 - 0x30 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000100", -- 1562 - 0x61a  :    4 - 0x4
    "00001101", -- 1563 - 0x61b  :   13 - 0xd
    "00001111", -- 1564 - 0x61c  :   15 - 0xf
    "00001100", -- 1565 - 0x61d  :   12 - 0xc
    "00001100", -- 1566 - 0x61e  :   12 - 0xc
    "00000100", -- 1567 - 0x61f  :    4 - 0x4
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00010000", -- 1570 - 0x622  :   16 - 0x10
    "01110000", -- 1571 - 0x623  :  112 - 0x70
    "11110000", -- 1572 - 0x624  :  240 - 0xf0
    "00110000", -- 1573 - 0x625  :   48 - 0x30
    "00110000", -- 1574 - 0x626  :   48 - 0x30
    "00010000", -- 1575 - 0x627  :   16 - 0x10
    "11100100", -- 1576 - 0x628  :  228 - 0xe4 -- Sprite 0xc5
    "00100100", -- 1577 - 0x629  :   36 - 0x24
    "11101111", -- 1578 - 0x62a  :  239 - 0xef
    "11100111", -- 1579 - 0x62b  :  231 - 0xe7
    "00000110", -- 1580 - 0x62c  :    6 - 0x6
    "00000100", -- 1581 - 0x62d  :    4 - 0x4
    "00000100", -- 1582 - 0x62e  :    4 - 0x4
    "00000111", -- 1583 - 0x62f  :    7 - 0x7
    "00010111", -- 1584 - 0x630  :   23 - 0x17 -- Sprite 0xc6
    "00010001", -- 1585 - 0x631  :   17 - 0x11
    "10110111", -- 1586 - 0x632  :  183 - 0xb7
    "11000111", -- 1587 - 0x633  :  199 - 0xc7
    "00100000", -- 1588 - 0x634  :   32 - 0x20
    "00100000", -- 1589 - 0x635  :   32 - 0x20
    "01100000", -- 1590 - 0x636  :   96 - 0x60
    "11100000", -- 1591 - 0x637  :  224 - 0xe0
    "00000111", -- 1592 - 0x638  :    7 - 0x7 -- Sprite 0xc7
    "00000011", -- 1593 - 0x639  :    3 - 0x3
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "11100000", -- 1596 - 0x63c  :  224 - 0xe0
    "00100000", -- 1597 - 0x63d  :   32 - 0x20
    "11100000", -- 1598 - 0x63e  :  224 - 0xe0
    "11100000", -- 1599 - 0x63f  :  224 - 0xe0
    "11100000", -- 1600 - 0x640  :  224 - 0xe0 -- Sprite 0xc8
    "11000000", -- 1601 - 0x641  :  192 - 0xc0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000111", -- 1604 - 0x644  :    7 - 0x7
    "00000001", -- 1605 - 0x645  :    1 - 0x1
    "00000111", -- 1606 - 0x646  :    7 - 0x7
    "00000111", -- 1607 - 0x647  :    7 - 0x7
    "00010011", -- 1608 - 0x648  :   19 - 0x13 -- Sprite 0xc9
    "00011111", -- 1609 - 0x649  :   31 - 0x1f
    "00001101", -- 1610 - 0x64a  :   13 - 0xd
    "00000100", -- 1611 - 0x64b  :    4 - 0x4
    "00001100", -- 1612 - 0x64c  :   12 - 0xc
    "00010011", -- 1613 - 0x64d  :   19 - 0x13
    "00011111", -- 1614 - 0x64e  :   31 - 0x1f
    "00000001", -- 1615 - 0x64f  :    1 - 0x1
    "01100000", -- 1616 - 0x650  :   96 - 0x60 -- Sprite 0xca
    "11110011", -- 1617 - 0x651  :  243 - 0xf3
    "10100111", -- 1618 - 0x652  :  167 - 0xa7
    "11000110", -- 1619 - 0x653  :  198 - 0xc6
    "01110100", -- 1620 - 0x654  :  116 - 0x74
    "00000100", -- 1621 - 0x655  :    4 - 0x4
    "10000111", -- 1622 - 0x656  :  135 - 0x87
    "10000111", -- 1623 - 0x657  :  135 - 0x87
    "00000110", -- 1624 - 0x658  :    6 - 0x6 -- Sprite 0xcb
    "10001111", -- 1625 - 0x659  :  143 - 0x8f
    "11000011", -- 1626 - 0x65a  :  195 - 0xc3
    "00100001", -- 1627 - 0x65b  :   33 - 0x21
    "00100000", -- 1628 - 0x65c  :   32 - 0x20
    "01100000", -- 1629 - 0x65d  :   96 - 0x60
    "11100000", -- 1630 - 0x65e  :  224 - 0xe0
    "11100000", -- 1631 - 0x65f  :  224 - 0xe0
    "11000011", -- 1632 - 0x660  :  195 - 0xc3 -- Sprite 0xcc
    "01110000", -- 1633 - 0x661  :  112 - 0x70
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "01100000", -- 1635 - 0x663  :   96 - 0x60
    "11110000", -- 1636 - 0x664  :  240 - 0xf0
    "11010000", -- 1637 - 0x665  :  208 - 0xd0
    "10010000", -- 1638 - 0x666  :  144 - 0x90
    "01100000", -- 1639 - 0x667  :   96 - 0x60
    "11000000", -- 1640 - 0x668  :  192 - 0xc0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000110", -- 1643 - 0x66b  :    6 - 0x6
    "00001111", -- 1644 - 0x66c  :   15 - 0xf
    "00001101", -- 1645 - 0x66d  :   13 - 0xd
    "00001001", -- 1646 - 0x66e  :    9 - 0x9
    "00000110", -- 1647 - 0x66f  :    6 - 0x6
    "11111100", -- 1648 - 0x670  :  252 - 0xfc -- Sprite 0xce
    "11000000", -- 1649 - 0x671  :  192 - 0xc0
    "11010001", -- 1650 - 0x672  :  209 - 0xd1
    "11000010", -- 1651 - 0x673  :  194 - 0xc2
    "10011110", -- 1652 - 0x674  :  158 - 0x9e
    "10111111", -- 1653 - 0x675  :  191 - 0xbf
    "10110000", -- 1654 - 0x676  :  176 - 0xb0
    "10110011", -- 1655 - 0x677  :  179 - 0xb3
    "00000111", -- 1656 - 0x678  :    7 - 0x7 -- Sprite 0xcf
    "11110011", -- 1657 - 0x679  :  243 - 0xf3
    "00001011", -- 1658 - 0x67a  :   11 - 0xb
    "01111011", -- 1659 - 0x67b  :  123 - 0x7b
    "01111011", -- 1660 - 0x67c  :  123 - 0x7b
    "11111001", -- 1661 - 0x67d  :  249 - 0xf9
    "00001101", -- 1662 - 0x67e  :   13 - 0xd
    "11101101", -- 1663 - 0x67f  :  237 - 0xed
    "11111111", -- 1664 - 0x680  :  255 - 0xff -- Sprite 0xd0
    "11111111", -- 1665 - 0x681  :  255 - 0xff
    "11111111", -- 1666 - 0x682  :  255 - 0xff
    "11111111", -- 1667 - 0x683  :  255 - 0xff
    "11101110", -- 1668 - 0x684  :  238 - 0xee
    "11101110", -- 1669 - 0x685  :  238 - 0xee
    "11101110", -- 1670 - 0x686  :  238 - 0xee
    "11101110", -- 1671 - 0x687  :  238 - 0xee
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Sprite 0xd1
    "11111111", -- 1673 - 0x689  :  255 - 0xff
    "11111111", -- 1674 - 0x68a  :  255 - 0xff
    "11111011", -- 1675 - 0x68b  :  251 - 0xfb
    "11111011", -- 1676 - 0x68c  :  251 - 0xfb
    "11111011", -- 1677 - 0x68d  :  251 - 0xfb
    "11111011", -- 1678 - 0x68e  :  251 - 0xfb
    "11111011", -- 1679 - 0x68f  :  251 - 0xfb
    "11111111", -- 1680 - 0x690  :  255 - 0xff -- Sprite 0xd2
    "11111111", -- 1681 - 0x691  :  255 - 0xff
    "11111111", -- 1682 - 0x692  :  255 - 0xff
    "11111111", -- 1683 - 0x693  :  255 - 0xff
    "11101110", -- 1684 - 0x694  :  238 - 0xee
    "10001110", -- 1685 - 0x695  :  142 - 0x8e
    "11111110", -- 1686 - 0x696  :  254 - 0xfe
    "11111110", -- 1687 - 0x697  :  254 - 0xfe
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11101110", -- 1692 - 0x69c  :  238 - 0xee
    "10001110", -- 1693 - 0x69d  :  142 - 0x8e
    "11111100", -- 1694 - 0x69e  :  252 - 0xfc
    "11111101", -- 1695 - 0x69f  :  253 - 0xfd
    "11111111", -- 1696 - 0x6a0  :  255 - 0xff -- Sprite 0xd4
    "11111111", -- 1697 - 0x6a1  :  255 - 0xff
    "11111111", -- 1698 - 0x6a2  :  255 - 0xff
    "11111110", -- 1699 - 0x6a3  :  254 - 0xfe
    "11101110", -- 1700 - 0x6a4  :  238 - 0xee
    "11101110", -- 1701 - 0x6a5  :  238 - 0xee
    "11101110", -- 1702 - 0x6a6  :  238 - 0xee
    "11101110", -- 1703 - 0x6a7  :  238 - 0xee
    "11111111", -- 1704 - 0x6a8  :  255 - 0xff -- Sprite 0xd5
    "11111111", -- 1705 - 0x6a9  :  255 - 0xff
    "11111111", -- 1706 - 0x6aa  :  255 - 0xff
    "11111101", -- 1707 - 0x6ab  :  253 - 0xfd
    "11100001", -- 1708 - 0x6ac  :  225 - 0xe1
    "11101111", -- 1709 - 0x6ad  :  239 - 0xef
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "11111111", -- 1712 - 0x6b0  :  255 - 0xff -- Sprite 0xd6
    "11111111", -- 1713 - 0x6b1  :  255 - 0xff
    "11111111", -- 1714 - 0x6b2  :  255 - 0xff
    "11111101", -- 1715 - 0x6b3  :  253 - 0xfd
    "11100001", -- 1716 - 0x6b4  :  225 - 0xe1
    "11101111", -- 1717 - 0x6b5  :  239 - 0xef
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111110", -- 1723 - 0x6bb  :  254 - 0xfe
    "11101110", -- 1724 - 0x6bc  :  238 - 0xee
    "10001110", -- 1725 - 0x6bd  :  142 - 0x8e
    "11111110", -- 1726 - 0x6be  :  254 - 0xfe
    "11111100", -- 1727 - 0x6bf  :  252 - 0xfc
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11101110", -- 1732 - 0x6c4  :  238 - 0xee
    "11101110", -- 1733 - 0x6c5  :  238 - 0xee
    "11111100", -- 1734 - 0x6c6  :  252 - 0xfc
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- Sprite 0xd9
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11101110", -- 1740 - 0x6cc  :  238 - 0xee
    "11101110", -- 1741 - 0x6cd  :  238 - 0xee
    "11101110", -- 1742 - 0x6ce  :  238 - 0xee
    "11101110", -- 1743 - 0x6cf  :  238 - 0xee
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "10000000", -- 1747 - 0x6d3  :  128 - 0x80
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000100", -- 1750 - 0x6d6  :    4 - 0x4
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Sprite 0xdb
    "00000100", -- 1753 - 0x6d9  :    4 - 0x4
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00010001", -- 1755 - 0x6db  :   17 - 0x11
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00100000", -- 1759 - 0x6df  :   32 - 0x20
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00100000", -- 1763 - 0x6e3  :   32 - 0x20
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000100", -- 1767 - 0x6e7  :    4 - 0x4
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00010001", -- 1770 - 0x6ea  :   17 - 0x11
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "10000000", -- 1773 - 0x6ed  :  128 - 0x80
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "10110011", -- 1776 - 0x6f0  :  179 - 0xb3 -- Sprite 0xde
    "10110011", -- 1777 - 0x6f1  :  179 - 0xb3
    "10110011", -- 1778 - 0x6f2  :  179 - 0xb3
    "10110011", -- 1779 - 0x6f3  :  179 - 0xb3
    "10110000", -- 1780 - 0x6f4  :  176 - 0xb0
    "10101111", -- 1781 - 0x6f5  :  175 - 0xaf
    "10011111", -- 1782 - 0x6f6  :  159 - 0x9f
    "11000000", -- 1783 - 0x6f7  :  192 - 0xc0
    "11101101", -- 1784 - 0x6f8  :  237 - 0xed -- Sprite 0xdf
    "11001101", -- 1785 - 0x6f9  :  205 - 0xcd
    "11001101", -- 1786 - 0x6fa  :  205 - 0xcd
    "00001101", -- 1787 - 0x6fb  :   13 - 0xd
    "00001101", -- 1788 - 0x6fc  :   13 - 0xd
    "11111101", -- 1789 - 0x6fd  :  253 - 0xfd
    "11111101", -- 1790 - 0x6fe  :  253 - 0xfd
    "00000011", -- 1791 - 0x6ff  :    3 - 0x3
    "11101110", -- 1792 - 0x700  :  238 - 0xee -- Sprite 0xe0
    "11101110", -- 1793 - 0x701  :  238 - 0xee
    "11101110", -- 1794 - 0x702  :  238 - 0xee
    "11101110", -- 1795 - 0x703  :  238 - 0xee
    "11111110", -- 1796 - 0x704  :  254 - 0xfe
    "11111100", -- 1797 - 0x705  :  252 - 0xfc
    "11000001", -- 1798 - 0x706  :  193 - 0xc1
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111011", -- 1800 - 0x708  :  251 - 0xfb -- Sprite 0xe1
    "11111011", -- 1801 - 0x709  :  251 - 0xfb
    "11111011", -- 1802 - 0x70a  :  251 - 0xfb
    "11111011", -- 1803 - 0x70b  :  251 - 0xfb
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111101", -- 1805 - 0x70d  :  253 - 0xfd
    "11000001", -- 1806 - 0x70e  :  193 - 0xc1
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111100", -- 1808 - 0x710  :  252 - 0xfc -- Sprite 0xe2
    "11100001", -- 1809 - 0x711  :  225 - 0xe1
    "11101111", -- 1810 - 0x712  :  239 - 0xef
    "11101111", -- 1811 - 0x713  :  239 - 0xef
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111110", -- 1813 - 0x715  :  254 - 0xfe
    "10000000", -- 1814 - 0x716  :  128 - 0x80
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11101110", -- 1816 - 0x718  :  238 - 0xee -- Sprite 0xe3
    "11111110", -- 1817 - 0x719  :  254 - 0xfe
    "11111110", -- 1818 - 0x71a  :  254 - 0xfe
    "11111110", -- 1819 - 0x71b  :  254 - 0xfe
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111100", -- 1821 - 0x71d  :  252 - 0xfc
    "11000001", -- 1822 - 0x71e  :  193 - 0xc1
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "11101110", -- 1824 - 0x720  :  238 - 0xee -- Sprite 0xe4
    "11101110", -- 1825 - 0x721  :  238 - 0xee
    "11111110", -- 1826 - 0x722  :  254 - 0xfe
    "11111110", -- 1827 - 0x723  :  254 - 0xfe
    "10001110", -- 1828 - 0x724  :  142 - 0x8e
    "11111110", -- 1829 - 0x725  :  254 - 0xfe
    "11111000", -- 1830 - 0x726  :  248 - 0xf8
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "10001110", -- 1832 - 0x728  :  142 - 0x8e -- Sprite 0xe5
    "11111110", -- 1833 - 0x729  :  254 - 0xfe
    "11111110", -- 1834 - 0x72a  :  254 - 0xfe
    "11111110", -- 1835 - 0x72b  :  254 - 0xfe
    "11111110", -- 1836 - 0x72c  :  254 - 0xfe
    "11111100", -- 1837 - 0x72d  :  252 - 0xfc
    "11000001", -- 1838 - 0x72e  :  193 - 0xc1
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11101110", -- 1840 - 0x730  :  238 - 0xee -- Sprite 0xe6
    "11101110", -- 1841 - 0x731  :  238 - 0xee
    "11101110", -- 1842 - 0x732  :  238 - 0xee
    "11101110", -- 1843 - 0x733  :  238 - 0xee
    "11111110", -- 1844 - 0x734  :  254 - 0xfe
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11000001", -- 1846 - 0x736  :  193 - 0xc1
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111101", -- 1848 - 0x738  :  253 - 0xfd -- Sprite 0xe7
    "11111101", -- 1849 - 0x739  :  253 - 0xfd
    "11111001", -- 1850 - 0x73a  :  249 - 0xf9
    "11111011", -- 1851 - 0x73b  :  251 - 0xfb
    "11111011", -- 1852 - 0x73c  :  251 - 0xfb
    "11111011", -- 1853 - 0x73d  :  251 - 0xfb
    "11100011", -- 1854 - 0x73e  :  227 - 0xe3
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "11101110", -- 1856 - 0x740  :  238 - 0xee -- Sprite 0xe8
    "11101110", -- 1857 - 0x741  :  238 - 0xee
    "11101110", -- 1858 - 0x742  :  238 - 0xee
    "11101110", -- 1859 - 0x743  :  238 - 0xee
    "11111110", -- 1860 - 0x744  :  254 - 0xfe
    "11111100", -- 1861 - 0x745  :  252 - 0xfc
    "11000001", -- 1862 - 0x746  :  193 - 0xc1
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11111110", -- 1864 - 0x748  :  254 - 0xfe -- Sprite 0xe9
    "11111110", -- 1865 - 0x749  :  254 - 0xfe
    "11001110", -- 1866 - 0x74a  :  206 - 0xce
    "11111110", -- 1867 - 0x74b  :  254 - 0xfe
    "11111110", -- 1868 - 0x74c  :  254 - 0xfe
    "11111100", -- 1869 - 0x74d  :  252 - 0xfc
    "11000001", -- 1870 - 0x74e  :  193 - 0xc1
    "11111111", -- 1871 - 0x74f  :  255 - 0xff
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0xea
    "01110000", -- 1873 - 0x751  :  112 - 0x70
    "00111000", -- 1874 - 0x752  :   56 - 0x38
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000010", -- 1876 - 0x754  :    2 - 0x2
    "00000111", -- 1877 - 0x755  :    7 - 0x7
    "00000011", -- 1878 - 0x756  :    3 - 0x3
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00001100", -- 1881 - 0x759  :   12 - 0xc
    "00000110", -- 1882 - 0x75a  :    6 - 0x6
    "00000110", -- 1883 - 0x75b  :    6 - 0x6
    "01100000", -- 1884 - 0x75c  :   96 - 0x60
    "01110000", -- 1885 - 0x75d  :  112 - 0x70
    "00110000", -- 1886 - 0x75e  :   48 - 0x30
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "11000000", -- 1889 - 0x761  :  192 - 0xc0
    "11100000", -- 1890 - 0x762  :  224 - 0xe0
    "01100000", -- 1891 - 0x763  :   96 - 0x60
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00001100", -- 1893 - 0x765  :   12 - 0xc
    "00001110", -- 1894 - 0x766  :   14 - 0xe
    "00000110", -- 1895 - 0x767  :    6 - 0x6
    "01100000", -- 1896 - 0x768  :   96 - 0x60 -- Sprite 0xed
    "01110000", -- 1897 - 0x769  :  112 - 0x70
    "00110000", -- 1898 - 0x76a  :   48 - 0x30
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00001100", -- 1901 - 0x76d  :   12 - 0xc
    "00001110", -- 1902 - 0x76e  :   14 - 0xe
    "00000110", -- 1903 - 0x76f  :    6 - 0x6
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Sprite 0xee
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "10111101", -- 1906 - 0x772  :  189 - 0xbd
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111011", -- 1909 - 0x775  :  251 - 0xfb
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "11111111", -- 1912 - 0x778  :  255 - 0xff -- Sprite 0xef
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111011", -- 1914 - 0x77a  :  251 - 0xfb
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11011111", -- 1916 - 0x77c  :  223 - 0xdf
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11111111", -- 1919 - 0x77f  :  255 - 0xff
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Sprite 0xf1
    "10000000", -- 1929 - 0x789  :  128 - 0x80
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "11000000", -- 1937 - 0x791  :  192 - 0xc0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Sprite 0xf3
    "11100000", -- 1945 - 0x799  :  224 - 0xe0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "11110000", -- 1953 - 0x7a1  :  240 - 0xf0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Sprite 0xf5
    "11111000", -- 1961 - 0x7a9  :  248 - 0xf8
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "11111100", -- 1969 - 0x7b1  :  252 - 0xfc
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "11111110", -- 1977 - 0x7b9  :  254 - 0xfe
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "10000000", -- 1996 - 0x7cc  :  128 - 0x80
    "10000000", -- 1997 - 0x7cd  :  128 - 0x80
    "11000000", -- 1998 - 0x7ce  :  192 - 0xc0
    "11000000", -- 1999 - 0x7cf  :  192 - 0xc0
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "00000001", -- 2012 - 0x7dc  :    1 - 0x1
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000010", -- 2014 - 0x7de  :    2 - 0x2
    "00000010", -- 2015 - 0x7df  :    2 - 0x2
    "11000000", -- 2016 - 0x7e0  :  192 - 0xc0 -- Sprite 0xfc
    "11000000", -- 2017 - 0x7e1  :  192 - 0xc0
    "10000000", -- 2018 - 0x7e2  :  128 - 0x80
    "10000000", -- 2019 - 0x7e3  :  128 - 0x80
    "11000000", -- 2020 - 0x7e4  :  192 - 0xc0
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "00000010", -- 2032 - 0x7f0  :    2 - 0x2 -- Sprite 0xfe
    "00000010", -- 2033 - 0x7f1  :    2 - 0x2
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
