------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : img_128.pgm 
--- Filas    : 128 
--- Columnas : 128 
--- Color    :  8 bits



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM8b_img_128 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(14-1 downto 0);
    dout : out std_logic_vector(8-1 downto 0) 
  );
end ROM8b_img_128;


architecture BEHAVIORAL of ROM8b_img_128 is
  signal addr_int  : natural range 0 to 2**14-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
       "11111111",
       "11101001",
       "11111111",
       "11000110",
       "11111111",
       "10010010",
       "11111111",
       "01010010",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "00111110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "01100100",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "01100100",
       "11111111",
       "10100000",
       "11111111",
       "11010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "01110100",
       "01110100",
       "01110100",
       "11111111",
       "11111111",
       "10101101",
       "10101101",
       "10101101",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "10100000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11101001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11011110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01010011",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "01100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "01111001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "00100111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000",
       "11111111",
       "00000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

