//-   Background Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_BG_PLN0
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 0
      11'h0: dout  = 8'b00111000; //    0 :  56 - 0x38 -- Background 0x0
      11'h1: dout  = 8'b01001100; //    1 :  76 - 0x4c
      11'h2: dout  = 8'b11000110; //    2 : 198 - 0xc6
      11'h3: dout  = 8'b11000110; //    3 : 198 - 0xc6
      11'h4: dout  = 8'b11000110; //    4 : 198 - 0xc6
      11'h5: dout  = 8'b01100100; //    5 : 100 - 0x64
      11'h6: dout  = 8'b00111000; //    6 :  56 - 0x38
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00011000; //    8 :  24 - 0x18 -- Background 0x1
      11'h9: dout  = 8'b00111000; //    9 :  56 - 0x38
      11'hA: dout  = 8'b00011000; //   10 :  24 - 0x18
      11'hB: dout  = 8'b00011000; //   11 :  24 - 0x18
      11'hC: dout  = 8'b00011000; //   12 :  24 - 0x18
      11'hD: dout  = 8'b00011000; //   13 :  24 - 0x18
      11'hE: dout  = 8'b01111110; //   14 : 126 - 0x7e
      11'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout  = 8'b01111100; //   16 : 124 - 0x7c -- Background 0x2
      11'h11: dout  = 8'b11000110; //   17 : 198 - 0xc6
      11'h12: dout  = 8'b00001110; //   18 :  14 - 0xe
      11'h13: dout  = 8'b00111100; //   19 :  60 - 0x3c
      11'h14: dout  = 8'b01111000; //   20 : 120 - 0x78
      11'h15: dout  = 8'b11100000; //   21 : 224 - 0xe0
      11'h16: dout  = 8'b11111110; //   22 : 254 - 0xfe
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b01111110; //   24 : 126 - 0x7e -- Background 0x3
      11'h19: dout  = 8'b00001100; //   25 :  12 - 0xc
      11'h1A: dout  = 8'b00011000; //   26 :  24 - 0x18
      11'h1B: dout  = 8'b00111100; //   27 :  60 - 0x3c
      11'h1C: dout  = 8'b00000110; //   28 :   6 - 0x6
      11'h1D: dout  = 8'b11000110; //   29 : 198 - 0xc6
      11'h1E: dout  = 8'b01111100; //   30 : 124 - 0x7c
      11'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout  = 8'b00011100; //   32 :  28 - 0x1c -- Background 0x4
      11'h21: dout  = 8'b00111100; //   33 :  60 - 0x3c
      11'h22: dout  = 8'b01101100; //   34 : 108 - 0x6c
      11'h23: dout  = 8'b11001100; //   35 : 204 - 0xcc
      11'h24: dout  = 8'b11111110; //   36 : 254 - 0xfe
      11'h25: dout  = 8'b00001100; //   37 :  12 - 0xc
      11'h26: dout  = 8'b00001100; //   38 :  12 - 0xc
      11'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout  = 8'b11111100; //   40 : 252 - 0xfc -- Background 0x5
      11'h29: dout  = 8'b11000000; //   41 : 192 - 0xc0
      11'h2A: dout  = 8'b11111100; //   42 : 252 - 0xfc
      11'h2B: dout  = 8'b00000110; //   43 :   6 - 0x6
      11'h2C: dout  = 8'b00000110; //   44 :   6 - 0x6
      11'h2D: dout  = 8'b11000110; //   45 : 198 - 0xc6
      11'h2E: dout  = 8'b01111100; //   46 : 124 - 0x7c
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00111100; //   48 :  60 - 0x3c -- Background 0x6
      11'h31: dout  = 8'b01100000; //   49 :  96 - 0x60
      11'h32: dout  = 8'b11000000; //   50 : 192 - 0xc0
      11'h33: dout  = 8'b11111100; //   51 : 252 - 0xfc
      11'h34: dout  = 8'b11000110; //   52 : 198 - 0xc6
      11'h35: dout  = 8'b11000110; //   53 : 198 - 0xc6
      11'h36: dout  = 8'b01111100; //   54 : 124 - 0x7c
      11'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout  = 8'b11111110; //   56 : 254 - 0xfe -- Background 0x7
      11'h39: dout  = 8'b11000110; //   57 : 198 - 0xc6
      11'h3A: dout  = 8'b00001100; //   58 :  12 - 0xc
      11'h3B: dout  = 8'b00011000; //   59 :  24 - 0x18
      11'h3C: dout  = 8'b00110000; //   60 :  48 - 0x30
      11'h3D: dout  = 8'b00110000; //   61 :  48 - 0x30
      11'h3E: dout  = 8'b00110000; //   62 :  48 - 0x30
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b01111100; //   64 : 124 - 0x7c -- Background 0x8
      11'h41: dout  = 8'b11000110; //   65 : 198 - 0xc6
      11'h42: dout  = 8'b11000110; //   66 : 198 - 0xc6
      11'h43: dout  = 8'b01111100; //   67 : 124 - 0x7c
      11'h44: dout  = 8'b11000110; //   68 : 198 - 0xc6
      11'h45: dout  = 8'b11000110; //   69 : 198 - 0xc6
      11'h46: dout  = 8'b01111100; //   70 : 124 - 0x7c
      11'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout  = 8'b01111100; //   72 : 124 - 0x7c -- Background 0x9
      11'h49: dout  = 8'b11000110; //   73 : 198 - 0xc6
      11'h4A: dout  = 8'b11000110; //   74 : 198 - 0xc6
      11'h4B: dout  = 8'b01111110; //   75 : 126 - 0x7e
      11'h4C: dout  = 8'b00000110; //   76 :   6 - 0x6
      11'h4D: dout  = 8'b00001100; //   77 :  12 - 0xc
      11'h4E: dout  = 8'b01111000; //   78 : 120 - 0x78
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00111000; //   80 :  56 - 0x38 -- Background 0xa
      11'h51: dout  = 8'b01101100; //   81 : 108 - 0x6c
      11'h52: dout  = 8'b11000110; //   82 : 198 - 0xc6
      11'h53: dout  = 8'b11000110; //   83 : 198 - 0xc6
      11'h54: dout  = 8'b11111110; //   84 : 254 - 0xfe
      11'h55: dout  = 8'b11000110; //   85 : 198 - 0xc6
      11'h56: dout  = 8'b11000110; //   86 : 198 - 0xc6
      11'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout  = 8'b11111100; //   88 : 252 - 0xfc -- Background 0xb
      11'h59: dout  = 8'b11000110; //   89 : 198 - 0xc6
      11'h5A: dout  = 8'b11000110; //   90 : 198 - 0xc6
      11'h5B: dout  = 8'b11111100; //   91 : 252 - 0xfc
      11'h5C: dout  = 8'b11000110; //   92 : 198 - 0xc6
      11'h5D: dout  = 8'b11000110; //   93 : 198 - 0xc6
      11'h5E: dout  = 8'b11111100; //   94 : 252 - 0xfc
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00111100; //   96 :  60 - 0x3c -- Background 0xc
      11'h61: dout  = 8'b01100110; //   97 : 102 - 0x66
      11'h62: dout  = 8'b11000000; //   98 : 192 - 0xc0
      11'h63: dout  = 8'b11000000; //   99 : 192 - 0xc0
      11'h64: dout  = 8'b11000000; //  100 : 192 - 0xc0
      11'h65: dout  = 8'b01100110; //  101 : 102 - 0x66
      11'h66: dout  = 8'b00111100; //  102 :  60 - 0x3c
      11'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout  = 8'b11111000; //  104 : 248 - 0xf8 -- Background 0xd
      11'h69: dout  = 8'b11001100; //  105 : 204 - 0xcc
      11'h6A: dout  = 8'b11000110; //  106 : 198 - 0xc6
      11'h6B: dout  = 8'b11000110; //  107 : 198 - 0xc6
      11'h6C: dout  = 8'b11000110; //  108 : 198 - 0xc6
      11'h6D: dout  = 8'b11001100; //  109 : 204 - 0xcc
      11'h6E: dout  = 8'b11111000; //  110 : 248 - 0xf8
      11'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout  = 8'b11111110; //  112 : 254 - 0xfe -- Background 0xe
      11'h71: dout  = 8'b11000000; //  113 : 192 - 0xc0
      11'h72: dout  = 8'b11000000; //  114 : 192 - 0xc0
      11'h73: dout  = 8'b11111100; //  115 : 252 - 0xfc
      11'h74: dout  = 8'b11000000; //  116 : 192 - 0xc0
      11'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      11'h76: dout  = 8'b11111110; //  118 : 254 - 0xfe
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b11111110; //  120 : 254 - 0xfe -- Background 0xf
      11'h79: dout  = 8'b11000000; //  121 : 192 - 0xc0
      11'h7A: dout  = 8'b11000000; //  122 : 192 - 0xc0
      11'h7B: dout  = 8'b11111100; //  123 : 252 - 0xfc
      11'h7C: dout  = 8'b11000000; //  124 : 192 - 0xc0
      11'h7D: dout  = 8'b11000000; //  125 : 192 - 0xc0
      11'h7E: dout  = 8'b11000000; //  126 : 192 - 0xc0
      11'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout  = 8'b00111110; //  128 :  62 - 0x3e -- Background 0x10
      11'h81: dout  = 8'b01100000; //  129 :  96 - 0x60
      11'h82: dout  = 8'b11000000; //  130 : 192 - 0xc0
      11'h83: dout  = 8'b11001110; //  131 : 206 - 0xce
      11'h84: dout  = 8'b11000110; //  132 : 198 - 0xc6
      11'h85: dout  = 8'b01100110; //  133 : 102 - 0x66
      11'h86: dout  = 8'b00111110; //  134 :  62 - 0x3e
      11'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout  = 8'b11000110; //  136 : 198 - 0xc6 -- Background 0x11
      11'h89: dout  = 8'b11000110; //  137 : 198 - 0xc6
      11'h8A: dout  = 8'b11000110; //  138 : 198 - 0xc6
      11'h8B: dout  = 8'b11111110; //  139 : 254 - 0xfe
      11'h8C: dout  = 8'b11000110; //  140 : 198 - 0xc6
      11'h8D: dout  = 8'b11000110; //  141 : 198 - 0xc6
      11'h8E: dout  = 8'b11000110; //  142 : 198 - 0xc6
      11'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout  = 8'b01111110; //  144 : 126 - 0x7e -- Background 0x12
      11'h91: dout  = 8'b00011000; //  145 :  24 - 0x18
      11'h92: dout  = 8'b00011000; //  146 :  24 - 0x18
      11'h93: dout  = 8'b00011000; //  147 :  24 - 0x18
      11'h94: dout  = 8'b00011000; //  148 :  24 - 0x18
      11'h95: dout  = 8'b00011000; //  149 :  24 - 0x18
      11'h96: dout  = 8'b01111110; //  150 : 126 - 0x7e
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b00011110; //  152 :  30 - 0x1e -- Background 0x13
      11'h99: dout  = 8'b00000110; //  153 :   6 - 0x6
      11'h9A: dout  = 8'b00000110; //  154 :   6 - 0x6
      11'h9B: dout  = 8'b00000110; //  155 :   6 - 0x6
      11'h9C: dout  = 8'b11000110; //  156 : 198 - 0xc6
      11'h9D: dout  = 8'b11000110; //  157 : 198 - 0xc6
      11'h9E: dout  = 8'b01111100; //  158 : 124 - 0x7c
      11'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout  = 8'b11000110; //  160 : 198 - 0xc6 -- Background 0x14
      11'hA1: dout  = 8'b11001100; //  161 : 204 - 0xcc
      11'hA2: dout  = 8'b11011000; //  162 : 216 - 0xd8
      11'hA3: dout  = 8'b11110000; //  163 : 240 - 0xf0
      11'hA4: dout  = 8'b11111000; //  164 : 248 - 0xf8
      11'hA5: dout  = 8'b11011100; //  165 : 220 - 0xdc
      11'hA6: dout  = 8'b11001110; //  166 : 206 - 0xce
      11'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout  = 8'b01100000; //  168 :  96 - 0x60 -- Background 0x15
      11'hA9: dout  = 8'b01100000; //  169 :  96 - 0x60
      11'hAA: dout  = 8'b01100000; //  170 :  96 - 0x60
      11'hAB: dout  = 8'b01100000; //  171 :  96 - 0x60
      11'hAC: dout  = 8'b01100000; //  172 :  96 - 0x60
      11'hAD: dout  = 8'b01100000; //  173 :  96 - 0x60
      11'hAE: dout  = 8'b01111110; //  174 : 126 - 0x7e
      11'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout  = 8'b11000110; //  176 : 198 - 0xc6 -- Background 0x16
      11'hB1: dout  = 8'b11101110; //  177 : 238 - 0xee
      11'hB2: dout  = 8'b11111110; //  178 : 254 - 0xfe
      11'hB3: dout  = 8'b11111110; //  179 : 254 - 0xfe
      11'hB4: dout  = 8'b11010110; //  180 : 214 - 0xd6
      11'hB5: dout  = 8'b11000110; //  181 : 198 - 0xc6
      11'hB6: dout  = 8'b11000110; //  182 : 198 - 0xc6
      11'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout  = 8'b11000110; //  184 : 198 - 0xc6 -- Background 0x17
      11'hB9: dout  = 8'b11100110; //  185 : 230 - 0xe6
      11'hBA: dout  = 8'b11110110; //  186 : 246 - 0xf6
      11'hBB: dout  = 8'b11111110; //  187 : 254 - 0xfe
      11'hBC: dout  = 8'b11011110; //  188 : 222 - 0xde
      11'hBD: dout  = 8'b11001110; //  189 : 206 - 0xce
      11'hBE: dout  = 8'b11000110; //  190 : 198 - 0xc6
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b01111100; //  192 : 124 - 0x7c -- Background 0x18
      11'hC1: dout  = 8'b11000110; //  193 : 198 - 0xc6
      11'hC2: dout  = 8'b11000110; //  194 : 198 - 0xc6
      11'hC3: dout  = 8'b11000110; //  195 : 198 - 0xc6
      11'hC4: dout  = 8'b11000110; //  196 : 198 - 0xc6
      11'hC5: dout  = 8'b11000110; //  197 : 198 - 0xc6
      11'hC6: dout  = 8'b01111100; //  198 : 124 - 0x7c
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b11111100; //  200 : 252 - 0xfc -- Background 0x19
      11'hC9: dout  = 8'b11000110; //  201 : 198 - 0xc6
      11'hCA: dout  = 8'b11000110; //  202 : 198 - 0xc6
      11'hCB: dout  = 8'b11000110; //  203 : 198 - 0xc6
      11'hCC: dout  = 8'b11111100; //  204 : 252 - 0xfc
      11'hCD: dout  = 8'b11000000; //  205 : 192 - 0xc0
      11'hCE: dout  = 8'b11000000; //  206 : 192 - 0xc0
      11'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout  = 8'b01111100; //  208 : 124 - 0x7c -- Background 0x1a
      11'hD1: dout  = 8'b11000110; //  209 : 198 - 0xc6
      11'hD2: dout  = 8'b11000110; //  210 : 198 - 0xc6
      11'hD3: dout  = 8'b11000110; //  211 : 198 - 0xc6
      11'hD4: dout  = 8'b11011110; //  212 : 222 - 0xde
      11'hD5: dout  = 8'b11001100; //  213 : 204 - 0xcc
      11'hD6: dout  = 8'b01111010; //  214 : 122 - 0x7a
      11'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout  = 8'b11111100; //  216 : 252 - 0xfc -- Background 0x1b
      11'hD9: dout  = 8'b11000110; //  217 : 198 - 0xc6
      11'hDA: dout  = 8'b11000110; //  218 : 198 - 0xc6
      11'hDB: dout  = 8'b11001110; //  219 : 206 - 0xce
      11'hDC: dout  = 8'b11111000; //  220 : 248 - 0xf8
      11'hDD: dout  = 8'b11011100; //  221 : 220 - 0xdc
      11'hDE: dout  = 8'b11001110; //  222 : 206 - 0xce
      11'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout  = 8'b01111000; //  224 : 120 - 0x78 -- Background 0x1c
      11'hE1: dout  = 8'b11001100; //  225 : 204 - 0xcc
      11'hE2: dout  = 8'b11000000; //  226 : 192 - 0xc0
      11'hE3: dout  = 8'b01111100; //  227 : 124 - 0x7c
      11'hE4: dout  = 8'b00000110; //  228 :   6 - 0x6
      11'hE5: dout  = 8'b11000110; //  229 : 198 - 0xc6
      11'hE6: dout  = 8'b01111100; //  230 : 124 - 0x7c
      11'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout  = 8'b01111110; //  232 : 126 - 0x7e -- Background 0x1d
      11'hE9: dout  = 8'b00011000; //  233 :  24 - 0x18
      11'hEA: dout  = 8'b00011000; //  234 :  24 - 0x18
      11'hEB: dout  = 8'b00011000; //  235 :  24 - 0x18
      11'hEC: dout  = 8'b00011000; //  236 :  24 - 0x18
      11'hED: dout  = 8'b00011000; //  237 :  24 - 0x18
      11'hEE: dout  = 8'b00011000; //  238 :  24 - 0x18
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b11000110; //  240 : 198 - 0xc6 -- Background 0x1e
      11'hF1: dout  = 8'b11000110; //  241 : 198 - 0xc6
      11'hF2: dout  = 8'b11000110; //  242 : 198 - 0xc6
      11'hF3: dout  = 8'b11000110; //  243 : 198 - 0xc6
      11'hF4: dout  = 8'b11000110; //  244 : 198 - 0xc6
      11'hF5: dout  = 8'b11000110; //  245 : 198 - 0xc6
      11'hF6: dout  = 8'b01111100; //  246 : 124 - 0x7c
      11'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout  = 8'b11000110; //  248 : 198 - 0xc6 -- Background 0x1f
      11'hF9: dout  = 8'b11000110; //  249 : 198 - 0xc6
      11'hFA: dout  = 8'b11000110; //  250 : 198 - 0xc6
      11'hFB: dout  = 8'b11101110; //  251 : 238 - 0xee
      11'hFC: dout  = 8'b01111100; //  252 : 124 - 0x7c
      11'hFD: dout  = 8'b00111000; //  253 :  56 - 0x38
      11'hFE: dout  = 8'b00010000; //  254 :  16 - 0x10
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b11000110; //  256 : 198 - 0xc6 -- Background 0x20
      11'h101: dout  = 8'b11000110; //  257 : 198 - 0xc6
      11'h102: dout  = 8'b11010110; //  258 : 214 - 0xd6
      11'h103: dout  = 8'b11111110; //  259 : 254 - 0xfe
      11'h104: dout  = 8'b11111110; //  260 : 254 - 0xfe
      11'h105: dout  = 8'b11101110; //  261 : 238 - 0xee
      11'h106: dout  = 8'b11000110; //  262 : 198 - 0xc6
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b11000110; //  264 : 198 - 0xc6 -- Background 0x21
      11'h109: dout  = 8'b11101110; //  265 : 238 - 0xee
      11'h10A: dout  = 8'b01111100; //  266 : 124 - 0x7c
      11'h10B: dout  = 8'b00111000; //  267 :  56 - 0x38
      11'h10C: dout  = 8'b01111100; //  268 : 124 - 0x7c
      11'h10D: dout  = 8'b11101110; //  269 : 238 - 0xee
      11'h10E: dout  = 8'b11000110; //  270 : 198 - 0xc6
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b01100110; //  272 : 102 - 0x66 -- Background 0x22
      11'h111: dout  = 8'b01100110; //  273 : 102 - 0x66
      11'h112: dout  = 8'b01100110; //  274 : 102 - 0x66
      11'h113: dout  = 8'b00111100; //  275 :  60 - 0x3c
      11'h114: dout  = 8'b00011000; //  276 :  24 - 0x18
      11'h115: dout  = 8'b00011000; //  277 :  24 - 0x18
      11'h116: dout  = 8'b00011000; //  278 :  24 - 0x18
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b11111110; //  280 : 254 - 0xfe -- Background 0x23
      11'h119: dout  = 8'b00001110; //  281 :  14 - 0xe
      11'h11A: dout  = 8'b00011100; //  282 :  28 - 0x1c
      11'h11B: dout  = 8'b00111000; //  283 :  56 - 0x38
      11'h11C: dout  = 8'b01110000; //  284 : 112 - 0x70
      11'h11D: dout  = 8'b11100000; //  285 : 224 - 0xe0
      11'h11E: dout  = 8'b11111110; //  286 : 254 - 0xfe
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Background 0x24
      11'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b11111111; //  296 : 255 - 0xff -- Background 0x25
      11'h129: dout  = 8'b11111111; //  297 : 255 - 0xff
      11'h12A: dout  = 8'b11111111; //  298 : 255 - 0xff
      11'h12B: dout  = 8'b11111111; //  299 : 255 - 0xff
      11'h12C: dout  = 8'b11111111; //  300 : 255 - 0xff
      11'h12D: dout  = 8'b11111111; //  301 : 255 - 0xff
      11'h12E: dout  = 8'b11111111; //  302 : 255 - 0xff
      11'h12F: dout  = 8'b11111111; //  303 : 255 - 0xff
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Background 0x26
      11'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      11'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      11'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      11'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout  = 8'b11111111; //  312 : 255 - 0xff -- Background 0x27
      11'h139: dout  = 8'b11111111; //  313 : 255 - 0xff
      11'h13A: dout  = 8'b11111111; //  314 : 255 - 0xff
      11'h13B: dout  = 8'b11111111; //  315 : 255 - 0xff
      11'h13C: dout  = 8'b11111111; //  316 : 255 - 0xff
      11'h13D: dout  = 8'b11111111; //  317 : 255 - 0xff
      11'h13E: dout  = 8'b11111111; //  318 : 255 - 0xff
      11'h13F: dout  = 8'b11111111; //  319 : 255 - 0xff
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout  = 8'b01111110; //  323 : 126 - 0x7e
      11'h144: dout  = 8'b01111110; //  324 : 126 - 0x7e
      11'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Background 0x29
      11'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      11'h14A: dout  = 8'b01000100; //  330 :  68 - 0x44
      11'h14B: dout  = 8'b00101000; //  331 :  40 - 0x28
      11'h14C: dout  = 8'b00010000; //  332 :  16 - 0x10
      11'h14D: dout  = 8'b00101000; //  333 :  40 - 0x28
      11'h14E: dout  = 8'b01000100; //  334 :  68 - 0x44
      11'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout  = 8'b11111111; //  336 : 255 - 0xff -- Background 0x2a
      11'h151: dout  = 8'b11111111; //  337 : 255 - 0xff
      11'h152: dout  = 8'b11111111; //  338 : 255 - 0xff
      11'h153: dout  = 8'b11111111; //  339 : 255 - 0xff
      11'h154: dout  = 8'b11111111; //  340 : 255 - 0xff
      11'h155: dout  = 8'b11111111; //  341 : 255 - 0xff
      11'h156: dout  = 8'b11111111; //  342 : 255 - 0xff
      11'h157: dout  = 8'b11111111; //  343 : 255 - 0xff
      11'h158: dout  = 8'b00011000; //  344 :  24 - 0x18 -- Background 0x2b
      11'h159: dout  = 8'b00111100; //  345 :  60 - 0x3c
      11'h15A: dout  = 8'b00111100; //  346 :  60 - 0x3c
      11'h15B: dout  = 8'b00111100; //  347 :  60 - 0x3c
      11'h15C: dout  = 8'b00011000; //  348 :  24 - 0x18
      11'h15D: dout  = 8'b00011000; //  349 :  24 - 0x18
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00011000; //  351 :  24 - 0x18
      11'h160: dout  = 8'b11111111; //  352 : 255 - 0xff -- Background 0x2c
      11'h161: dout  = 8'b01111111; //  353 : 127 - 0x7f
      11'h162: dout  = 8'b01111111; //  354 : 127 - 0x7f
      11'h163: dout  = 8'b01111111; //  355 : 127 - 0x7f
      11'h164: dout  = 8'b01111111; //  356 : 127 - 0x7f
      11'h165: dout  = 8'b11111111; //  357 : 255 - 0xff
      11'h166: dout  = 8'b11100011; //  358 : 227 - 0xe3
      11'h167: dout  = 8'b11000001; //  359 : 193 - 0xc1
      11'h168: dout  = 8'b10000000; //  360 : 128 - 0x80 -- Background 0x2d
      11'h169: dout  = 8'b10000000; //  361 : 128 - 0x80
      11'h16A: dout  = 8'b10000000; //  362 : 128 - 0x80
      11'h16B: dout  = 8'b11000001; //  363 : 193 - 0xc1
      11'h16C: dout  = 8'b11100011; //  364 : 227 - 0xe3
      11'h16D: dout  = 8'b11111111; //  365 : 255 - 0xff
      11'h16E: dout  = 8'b11111111; //  366 : 255 - 0xff
      11'h16F: dout  = 8'b11111111; //  367 : 255 - 0xff
      11'h170: dout  = 8'b00111000; //  368 :  56 - 0x38 -- Background 0x2e
      11'h171: dout  = 8'b01111100; //  369 : 124 - 0x7c
      11'h172: dout  = 8'b01111100; //  370 : 124 - 0x7c
      11'h173: dout  = 8'b01111100; //  371 : 124 - 0x7c
      11'h174: dout  = 8'b01111100; //  372 : 124 - 0x7c
      11'h175: dout  = 8'b01111100; //  373 : 124 - 0x7c
      11'h176: dout  = 8'b00111000; //  374 :  56 - 0x38
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b00000011; //  376 :   3 - 0x3 -- Background 0x2f
      11'h179: dout  = 8'b00000110; //  377 :   6 - 0x6
      11'h17A: dout  = 8'b00001100; //  378 :  12 - 0xc
      11'h17B: dout  = 8'b00001100; //  379 :  12 - 0xc
      11'h17C: dout  = 8'b00001000; //  380 :   8 - 0x8
      11'h17D: dout  = 8'b00001000; //  381 :   8 - 0x8
      11'h17E: dout  = 8'b00000100; //  382 :   4 - 0x4
      11'h17F: dout  = 8'b00000011; //  383 :   3 - 0x3
      11'h180: dout  = 8'b00000001; //  384 :   1 - 0x1 -- Background 0x30
      11'h181: dout  = 8'b00000010; //  385 :   2 - 0x2
      11'h182: dout  = 8'b00000100; //  386 :   4 - 0x4
      11'h183: dout  = 8'b00001000; //  387 :   8 - 0x8
      11'h184: dout  = 8'b00010000; //  388 :  16 - 0x10
      11'h185: dout  = 8'b00100000; //  389 :  32 - 0x20
      11'h186: dout  = 8'b01000000; //  390 :  64 - 0x40
      11'h187: dout  = 8'b10000000; //  391 : 128 - 0x80
      11'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- Background 0x31
      11'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      11'h18D: dout  = 8'b00000111; //  397 :   7 - 0x7
      11'h18E: dout  = 8'b00111000; //  398 :  56 - 0x38
      11'h18F: dout  = 8'b11000000; //  399 : 192 - 0xc0
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Background 0x32
      11'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout  = 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout  = 8'b00000000; //  404 :   0 - 0x0
      11'h195: dout  = 8'b11100000; //  405 : 224 - 0xe0
      11'h196: dout  = 8'b00011100; //  406 :  28 - 0x1c
      11'h197: dout  = 8'b00000011; //  407 :   3 - 0x3
      11'h198: dout  = 8'b10000000; //  408 : 128 - 0x80 -- Background 0x33
      11'h199: dout  = 8'b01000000; //  409 :  64 - 0x40
      11'h19A: dout  = 8'b00100000; //  410 :  32 - 0x20
      11'h19B: dout  = 8'b00010000; //  411 :  16 - 0x10
      11'h19C: dout  = 8'b00001000; //  412 :   8 - 0x8
      11'h19D: dout  = 8'b00000100; //  413 :   4 - 0x4
      11'h19E: dout  = 8'b00000010; //  414 :   2 - 0x2
      11'h19F: dout  = 8'b00000001; //  415 :   1 - 0x1
      11'h1A0: dout  = 8'b00000100; //  416 :   4 - 0x4 -- Background 0x34
      11'h1A1: dout  = 8'b00001110; //  417 :  14 - 0xe
      11'h1A2: dout  = 8'b00001110; //  418 :  14 - 0xe
      11'h1A3: dout  = 8'b00001110; //  419 :  14 - 0xe
      11'h1A4: dout  = 8'b01101110; //  420 : 110 - 0x6e
      11'h1A5: dout  = 8'b01100100; //  421 : 100 - 0x64
      11'h1A6: dout  = 8'b01100000; //  422 :  96 - 0x60
      11'h1A7: dout  = 8'b01100000; //  423 :  96 - 0x60
      11'h1A8: dout  = 8'b00000111; //  424 :   7 - 0x7 -- Background 0x35
      11'h1A9: dout  = 8'b00001111; //  425 :  15 - 0xf
      11'h1AA: dout  = 8'b00011111; //  426 :  31 - 0x1f
      11'h1AB: dout  = 8'b00011111; //  427 :  31 - 0x1f
      11'h1AC: dout  = 8'b01111111; //  428 : 127 - 0x7f
      11'h1AD: dout  = 8'b11111111; //  429 : 255 - 0xff
      11'h1AE: dout  = 8'b11111111; //  430 : 255 - 0xff
      11'h1AF: dout  = 8'b01111111; //  431 : 127 - 0x7f
      11'h1B0: dout  = 8'b00000011; //  432 :   3 - 0x3 -- Background 0x36
      11'h1B1: dout  = 8'b00000111; //  433 :   7 - 0x7
      11'h1B2: dout  = 8'b00011111; //  434 :  31 - 0x1f
      11'h1B3: dout  = 8'b00111111; //  435 :  63 - 0x3f
      11'h1B4: dout  = 8'b00111111; //  436 :  63 - 0x3f
      11'h1B5: dout  = 8'b00111111; //  437 :  63 - 0x3f
      11'h1B6: dout  = 8'b01111001; //  438 : 121 - 0x79
      11'h1B7: dout  = 8'b11110111; //  439 : 247 - 0xf7
      11'h1B8: dout  = 8'b11000000; //  440 : 192 - 0xc0 -- Background 0x37
      11'h1B9: dout  = 8'b11100000; //  441 : 224 - 0xe0
      11'h1BA: dout  = 8'b11110000; //  442 : 240 - 0xf0
      11'h1BB: dout  = 8'b11110100; //  443 : 244 - 0xf4
      11'h1BC: dout  = 8'b11111110; //  444 : 254 - 0xfe
      11'h1BD: dout  = 8'b10111111; //  445 : 191 - 0xbf
      11'h1BE: dout  = 8'b11011111; //  446 : 223 - 0xdf
      11'h1BF: dout  = 8'b11111111; //  447 : 255 - 0xff
      11'h1C0: dout  = 8'b10010000; //  448 : 144 - 0x90 -- Background 0x38
      11'h1C1: dout  = 8'b10111000; //  449 : 184 - 0xb8
      11'h1C2: dout  = 8'b11111000; //  450 : 248 - 0xf8
      11'h1C3: dout  = 8'b11111010; //  451 : 250 - 0xfa
      11'h1C4: dout  = 8'b11111111; //  452 : 255 - 0xff
      11'h1C5: dout  = 8'b11111111; //  453 : 255 - 0xff
      11'h1C6: dout  = 8'b11111111; //  454 : 255 - 0xff
      11'h1C7: dout  = 8'b11111110; //  455 : 254 - 0xfe
      11'h1C8: dout  = 8'b00111011; //  456 :  59 - 0x3b -- Background 0x39
      11'h1C9: dout  = 8'b00011101; //  457 :  29 - 0x1d
      11'h1CA: dout  = 8'b00001110; //  458 :  14 - 0xe
      11'h1CB: dout  = 8'b00001111; //  459 :  15 - 0xf
      11'h1CC: dout  = 8'b00000111; //  460 :   7 - 0x7
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b11111111; //  464 : 255 - 0xff -- Background 0x3a
      11'h1D1: dout  = 8'b10111111; //  465 : 191 - 0xbf
      11'h1D2: dout  = 8'b00011100; //  466 :  28 - 0x1c
      11'h1D3: dout  = 8'b11000000; //  467 : 192 - 0xc0
      11'h1D4: dout  = 8'b11110011; //  468 : 243 - 0xf3
      11'h1D5: dout  = 8'b11111111; //  469 : 255 - 0xff
      11'h1D6: dout  = 8'b01111110; //  470 : 126 - 0x7e
      11'h1D7: dout  = 8'b00011100; //  471 :  28 - 0x1c
      11'h1D8: dout  = 8'b10111111; //  472 : 191 - 0xbf -- Background 0x3b
      11'h1D9: dout  = 8'b01111111; //  473 : 127 - 0x7f
      11'h1DA: dout  = 8'b00111101; //  474 :  61 - 0x3d
      11'h1DB: dout  = 8'b10000011; //  475 : 131 - 0x83
      11'h1DC: dout  = 8'b11000111; //  476 : 199 - 0xc7
      11'h1DD: dout  = 8'b11111111; //  477 : 255 - 0xff
      11'h1DE: dout  = 8'b11111111; //  478 : 255 - 0xff
      11'h1DF: dout  = 8'b00111100; //  479 :  60 - 0x3c
      11'h1E0: dout  = 8'b11111100; //  480 : 252 - 0xfc -- Background 0x3c
      11'h1E1: dout  = 8'b11111110; //  481 : 254 - 0xfe
      11'h1E2: dout  = 8'b11111111; //  482 : 255 - 0xff
      11'h1E3: dout  = 8'b11111110; //  483 : 254 - 0xfe
      11'h1E4: dout  = 8'b11111110; //  484 : 254 - 0xfe
      11'h1E5: dout  = 8'b11111000; //  485 : 248 - 0xf8
      11'h1E6: dout  = 8'b01100000; //  486 :  96 - 0x60
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b11000000; //  488 : 192 - 0xc0 -- Background 0x3d
      11'h1E9: dout  = 8'b00100000; //  489 :  32 - 0x20
      11'h1EA: dout  = 8'b00010000; //  490 :  16 - 0x10
      11'h1EB: dout  = 8'b00010000; //  491 :  16 - 0x10
      11'h1EC: dout  = 8'b00010000; //  492 :  16 - 0x10
      11'h1ED: dout  = 8'b00010000; //  493 :  16 - 0x10
      11'h1EE: dout  = 8'b00100000; //  494 :  32 - 0x20
      11'h1EF: dout  = 8'b11000000; //  495 : 192 - 0xc0
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout  = 8'b00111111; //  500 :  63 - 0x3f
      11'h1F5: dout  = 8'b01111111; //  501 : 127 - 0x7f
      11'h1F6: dout  = 8'b11100000; //  502 : 224 - 0xe0
      11'h1F7: dout  = 8'b11000000; //  503 : 192 - 0xc0
      11'h1F8: dout  = 8'b10001000; //  504 : 136 - 0x88 -- Background 0x3f
      11'h1F9: dout  = 8'b10011100; //  505 : 156 - 0x9c
      11'h1FA: dout  = 8'b10001000; //  506 : 136 - 0x88
      11'h1FB: dout  = 8'b10000000; //  507 : 128 - 0x80
      11'h1FC: dout  = 8'b10000000; //  508 : 128 - 0x80
      11'h1FD: dout  = 8'b10000000; //  509 : 128 - 0x80
      11'h1FE: dout  = 8'b10000000; //  510 : 128 - 0x80
      11'h1FF: dout  = 8'b10000000; //  511 : 128 - 0x80
      11'h200: dout  = 8'b11111110; //  512 : 254 - 0xfe -- Background 0x40
      11'h201: dout  = 8'b11111110; //  513 : 254 - 0xfe
      11'h202: dout  = 8'b11111110; //  514 : 254 - 0xfe
      11'h203: dout  = 8'b11111110; //  515 : 254 - 0xfe
      11'h204: dout  = 8'b11111110; //  516 : 254 - 0xfe
      11'h205: dout  = 8'b11111110; //  517 : 254 - 0xfe
      11'h206: dout  = 8'b11111110; //  518 : 254 - 0xfe
      11'h207: dout  = 8'b11111110; //  519 : 254 - 0xfe
      11'h208: dout  = 8'b00001000; //  520 :   8 - 0x8 -- Background 0x41
      11'h209: dout  = 8'b00010100; //  521 :  20 - 0x14
      11'h20A: dout  = 8'b00100100; //  522 :  36 - 0x24
      11'h20B: dout  = 8'b11000100; //  523 : 196 - 0xc4
      11'h20C: dout  = 8'b00000011; //  524 :   3 - 0x3
      11'h20D: dout  = 8'b01000000; //  525 :  64 - 0x40
      11'h20E: dout  = 8'b10100001; //  526 : 161 - 0xa1
      11'h20F: dout  = 8'b00100110; //  527 :  38 - 0x26
      11'h210: dout  = 8'b11111111; //  528 : 255 - 0xff -- Background 0x42
      11'h211: dout  = 8'b11111111; //  529 : 255 - 0xff
      11'h212: dout  = 8'b11111111; //  530 : 255 - 0xff
      11'h213: dout  = 8'b11111111; //  531 : 255 - 0xff
      11'h214: dout  = 8'b01111111; //  532 : 127 - 0x7f
      11'h215: dout  = 8'b01111111; //  533 : 127 - 0x7f
      11'h216: dout  = 8'b01111111; //  534 : 127 - 0x7f
      11'h217: dout  = 8'b01111111; //  535 : 127 - 0x7f
      11'h218: dout  = 8'b11111111; //  536 : 255 - 0xff -- Background 0x43
      11'h219: dout  = 8'b11111111; //  537 : 255 - 0xff
      11'h21A: dout  = 8'b11111111; //  538 : 255 - 0xff
      11'h21B: dout  = 8'b11111111; //  539 : 255 - 0xff
      11'h21C: dout  = 8'b11111111; //  540 : 255 - 0xff
      11'h21D: dout  = 8'b11111111; //  541 : 255 - 0xff
      11'h21E: dout  = 8'b11111111; //  542 : 255 - 0xff
      11'h21F: dout  = 8'b11111111; //  543 : 255 - 0xff
      11'h220: dout  = 8'b01111111; //  544 : 127 - 0x7f -- Background 0x44
      11'h221: dout  = 8'b10000000; //  545 : 128 - 0x80
      11'h222: dout  = 8'b10000000; //  546 : 128 - 0x80
      11'h223: dout  = 8'b10011000; //  547 : 152 - 0x98
      11'h224: dout  = 8'b10011100; //  548 : 156 - 0x9c
      11'h225: dout  = 8'b10001100; //  549 : 140 - 0x8c
      11'h226: dout  = 8'b10000000; //  550 : 128 - 0x80
      11'h227: dout  = 8'b10000000; //  551 : 128 - 0x80
      11'h228: dout  = 8'b11111111; //  552 : 255 - 0xff -- Background 0x45
      11'h229: dout  = 8'b00000001; //  553 :   1 - 0x1
      11'h22A: dout  = 8'b00000001; //  554 :   1 - 0x1
      11'h22B: dout  = 8'b11111111; //  555 : 255 - 0xff
      11'h22C: dout  = 8'b00010000; //  556 :  16 - 0x10
      11'h22D: dout  = 8'b00010000; //  557 :  16 - 0x10
      11'h22E: dout  = 8'b00010000; //  558 :  16 - 0x10
      11'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      11'h230: dout  = 8'b10000000; //  560 : 128 - 0x80 -- Background 0x46
      11'h231: dout  = 8'b10000000; //  561 : 128 - 0x80
      11'h232: dout  = 8'b10000000; //  562 : 128 - 0x80
      11'h233: dout  = 8'b10000000; //  563 : 128 - 0x80
      11'h234: dout  = 8'b10000000; //  564 : 128 - 0x80
      11'h235: dout  = 8'b10000000; //  565 : 128 - 0x80
      11'h236: dout  = 8'b10000000; //  566 : 128 - 0x80
      11'h237: dout  = 8'b10000000; //  567 : 128 - 0x80
      11'h238: dout  = 8'b00000001; //  568 :   1 - 0x1 -- Background 0x47
      11'h239: dout  = 8'b00000001; //  569 :   1 - 0x1
      11'h23A: dout  = 8'b00000001; //  570 :   1 - 0x1
      11'h23B: dout  = 8'b11111111; //  571 : 255 - 0xff
      11'h23C: dout  = 8'b00010000; //  572 :  16 - 0x10
      11'h23D: dout  = 8'b00010000; //  573 :  16 - 0x10
      11'h23E: dout  = 8'b00010000; //  574 :  16 - 0x10
      11'h23F: dout  = 8'b11111111; //  575 : 255 - 0xff
      11'h240: dout  = 8'b11111111; //  576 : 255 - 0xff -- Background 0x48
      11'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      11'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      11'h243: dout  = 8'b00000000; //  579 :   0 - 0x0
      11'h244: dout  = 8'b00000000; //  580 :   0 - 0x0
      11'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      11'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b11111110; //  584 : 254 - 0xfe -- Background 0x49
      11'h249: dout  = 8'b00000001; //  585 :   1 - 0x1
      11'h24A: dout  = 8'b00000001; //  586 :   1 - 0x1
      11'h24B: dout  = 8'b00011001; //  587 :  25 - 0x19
      11'h24C: dout  = 8'b00011101; //  588 :  29 - 0x1d
      11'h24D: dout  = 8'b00001101; //  589 :  13 - 0xd
      11'h24E: dout  = 8'b00000001; //  590 :   1 - 0x1
      11'h24F: dout  = 8'b00000001; //  591 :   1 - 0x1
      11'h250: dout  = 8'b00000001; //  592 :   1 - 0x1 -- Background 0x4a
      11'h251: dout  = 8'b00000001; //  593 :   1 - 0x1
      11'h252: dout  = 8'b00000001; //  594 :   1 - 0x1
      11'h253: dout  = 8'b00000001; //  595 :   1 - 0x1
      11'h254: dout  = 8'b00000001; //  596 :   1 - 0x1
      11'h255: dout  = 8'b00000001; //  597 :   1 - 0x1
      11'h256: dout  = 8'b00000001; //  598 :   1 - 0x1
      11'h257: dout  = 8'b00000001; //  599 :   1 - 0x1
      11'h258: dout  = 8'b00111111; //  600 :  63 - 0x3f -- Background 0x4b
      11'h259: dout  = 8'b01111111; //  601 : 127 - 0x7f
      11'h25A: dout  = 8'b01111111; //  602 : 127 - 0x7f
      11'h25B: dout  = 8'b11111111; //  603 : 255 - 0xff
      11'h25C: dout  = 8'b11111111; //  604 : 255 - 0xff
      11'h25D: dout  = 8'b11111111; //  605 : 255 - 0xff
      11'h25E: dout  = 8'b11111111; //  606 : 255 - 0xff
      11'h25F: dout  = 8'b11111111; //  607 : 255 - 0xff
      11'h260: dout  = 8'b11111111; //  608 : 255 - 0xff -- Background 0x4c
      11'h261: dout  = 8'b11111111; //  609 : 255 - 0xff
      11'h262: dout  = 8'b11111111; //  610 : 255 - 0xff
      11'h263: dout  = 8'b11111111; //  611 : 255 - 0xff
      11'h264: dout  = 8'b11111111; //  612 : 255 - 0xff
      11'h265: dout  = 8'b11111111; //  613 : 255 - 0xff
      11'h266: dout  = 8'b01111110; //  614 : 126 - 0x7e
      11'h267: dout  = 8'b00111100; //  615 :  60 - 0x3c
      11'h268: dout  = 8'b11111111; //  616 : 255 - 0xff -- Background 0x4d
      11'h269: dout  = 8'b11111111; //  617 : 255 - 0xff
      11'h26A: dout  = 8'b11111111; //  618 : 255 - 0xff
      11'h26B: dout  = 8'b11111111; //  619 : 255 - 0xff
      11'h26C: dout  = 8'b11111111; //  620 : 255 - 0xff
      11'h26D: dout  = 8'b11111111; //  621 : 255 - 0xff
      11'h26E: dout  = 8'b11111111; //  622 : 255 - 0xff
      11'h26F: dout  = 8'b11111111; //  623 : 255 - 0xff
      11'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Background 0x4e
      11'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      11'h272: dout  = 8'b11111111; //  626 : 255 - 0xff
      11'h273: dout  = 8'b11111111; //  627 : 255 - 0xff
      11'h274: dout  = 8'b11111111; //  628 : 255 - 0xff
      11'h275: dout  = 8'b11111111; //  629 : 255 - 0xff
      11'h276: dout  = 8'b11111110; //  630 : 254 - 0xfe
      11'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      11'h278: dout  = 8'b11111111; //  632 : 255 - 0xff -- Background 0x4f
      11'h279: dout  = 8'b11111111; //  633 : 255 - 0xff
      11'h27A: dout  = 8'b11111111; //  634 : 255 - 0xff
      11'h27B: dout  = 8'b11111111; //  635 : 255 - 0xff
      11'h27C: dout  = 8'b11111111; //  636 : 255 - 0xff
      11'h27D: dout  = 8'b11111111; //  637 : 255 - 0xff
      11'h27E: dout  = 8'b11111110; //  638 : 254 - 0xfe
      11'h27F: dout  = 8'b01111100; //  639 : 124 - 0x7c
      11'h280: dout  = 8'b11111000; //  640 : 248 - 0xf8 -- Background 0x50
      11'h281: dout  = 8'b11111100; //  641 : 252 - 0xfc
      11'h282: dout  = 8'b11111110; //  642 : 254 - 0xfe
      11'h283: dout  = 8'b11111110; //  643 : 254 - 0xfe
      11'h284: dout  = 8'b11111111; //  644 : 255 - 0xff
      11'h285: dout  = 8'b11111111; //  645 : 255 - 0xff
      11'h286: dout  = 8'b11111111; //  646 : 255 - 0xff
      11'h287: dout  = 8'b11111111; //  647 : 255 - 0xff
      11'h288: dout  = 8'b11111111; //  648 : 255 - 0xff -- Background 0x51
      11'h289: dout  = 8'b11111111; //  649 : 255 - 0xff
      11'h28A: dout  = 8'b11111111; //  650 : 255 - 0xff
      11'h28B: dout  = 8'b11111111; //  651 : 255 - 0xff
      11'h28C: dout  = 8'b11111111; //  652 : 255 - 0xff
      11'h28D: dout  = 8'b11111111; //  653 : 255 - 0xff
      11'h28E: dout  = 8'b01111110; //  654 : 126 - 0x7e
      11'h28F: dout  = 8'b00111100; //  655 :  60 - 0x3c
      11'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Background 0x52
      11'h291: dout  = 8'b00001000; //  657 :   8 - 0x8
      11'h292: dout  = 8'b00001000; //  658 :   8 - 0x8
      11'h293: dout  = 8'b00001000; //  659 :   8 - 0x8
      11'h294: dout  = 8'b00010000; //  660 :  16 - 0x10
      11'h295: dout  = 8'b00010000; //  661 :  16 - 0x10
      11'h296: dout  = 8'b00010000; //  662 :  16 - 0x10
      11'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      11'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Background 0x53
      11'h299: dout  = 8'b01111111; //  665 : 127 - 0x7f
      11'h29A: dout  = 8'b01111111; //  666 : 127 - 0x7f
      11'h29B: dout  = 8'b01111000; //  667 : 120 - 0x78
      11'h29C: dout  = 8'b01110011; //  668 : 115 - 0x73
      11'h29D: dout  = 8'b01110011; //  669 : 115 - 0x73
      11'h29E: dout  = 8'b01110011; //  670 : 115 - 0x73
      11'h29F: dout  = 8'b01111111; //  671 : 127 - 0x7f
      11'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Background 0x54
      11'h2A1: dout  = 8'b11111111; //  673 : 255 - 0xff
      11'h2A2: dout  = 8'b11111111; //  674 : 255 - 0xff
      11'h2A3: dout  = 8'b00111111; //  675 :  63 - 0x3f
      11'h2A4: dout  = 8'b10011111; //  676 : 159 - 0x9f
      11'h2A5: dout  = 8'b10011111; //  677 : 159 - 0x9f
      11'h2A6: dout  = 8'b10011111; //  678 : 159 - 0x9f
      11'h2A7: dout  = 8'b00011111; //  679 :  31 - 0x1f
      11'h2A8: dout  = 8'b01111110; //  680 : 126 - 0x7e -- Background 0x55
      11'h2A9: dout  = 8'b01111110; //  681 : 126 - 0x7e
      11'h2AA: dout  = 8'b01111111; //  682 : 127 - 0x7f
      11'h2AB: dout  = 8'b01111110; //  683 : 126 - 0x7e
      11'h2AC: dout  = 8'b01111110; //  684 : 126 - 0x7e
      11'h2AD: dout  = 8'b01111111; //  685 : 127 - 0x7f
      11'h2AE: dout  = 8'b01111111; //  686 : 127 - 0x7f
      11'h2AF: dout  = 8'b11111111; //  687 : 255 - 0xff
      11'h2B0: dout  = 8'b01111111; //  688 : 127 - 0x7f -- Background 0x56
      11'h2B1: dout  = 8'b01111111; //  689 : 127 - 0x7f
      11'h2B2: dout  = 8'b11111111; //  690 : 255 - 0xff
      11'h2B3: dout  = 8'b01111111; //  691 : 127 - 0x7f
      11'h2B4: dout  = 8'b01111111; //  692 : 127 - 0x7f
      11'h2B5: dout  = 8'b11111111; //  693 : 255 - 0xff
      11'h2B6: dout  = 8'b11111111; //  694 : 255 - 0xff
      11'h2B7: dout  = 8'b11111111; //  695 : 255 - 0xff
      11'h2B8: dout  = 8'b01111111; //  696 : 127 - 0x7f -- Background 0x57
      11'h2B9: dout  = 8'b10000000; //  697 : 128 - 0x80
      11'h2BA: dout  = 8'b10100000; //  698 : 160 - 0xa0
      11'h2BB: dout  = 8'b10000000; //  699 : 128 - 0x80
      11'h2BC: dout  = 8'b10000000; //  700 : 128 - 0x80
      11'h2BD: dout  = 8'b10000000; //  701 : 128 - 0x80
      11'h2BE: dout  = 8'b10000000; //  702 : 128 - 0x80
      11'h2BF: dout  = 8'b10000000; //  703 : 128 - 0x80
      11'h2C0: dout  = 8'b11111110; //  704 : 254 - 0xfe -- Background 0x58
      11'h2C1: dout  = 8'b00000001; //  705 :   1 - 0x1
      11'h2C2: dout  = 8'b00000101; //  706 :   5 - 0x5
      11'h2C3: dout  = 8'b00000001; //  707 :   1 - 0x1
      11'h2C4: dout  = 8'b00000001; //  708 :   1 - 0x1
      11'h2C5: dout  = 8'b00000001; //  709 :   1 - 0x1
      11'h2C6: dout  = 8'b00000001; //  710 :   1 - 0x1
      11'h2C7: dout  = 8'b00000001; //  711 :   1 - 0x1
      11'h2C8: dout  = 8'b10000000; //  712 : 128 - 0x80 -- Background 0x59
      11'h2C9: dout  = 8'b10000000; //  713 : 128 - 0x80
      11'h2CA: dout  = 8'b10000000; //  714 : 128 - 0x80
      11'h2CB: dout  = 8'b10000000; //  715 : 128 - 0x80
      11'h2CC: dout  = 8'b10000000; //  716 : 128 - 0x80
      11'h2CD: dout  = 8'b10100000; //  717 : 160 - 0xa0
      11'h2CE: dout  = 8'b10000000; //  718 : 128 - 0x80
      11'h2CF: dout  = 8'b01111111; //  719 : 127 - 0x7f
      11'h2D0: dout  = 8'b00000001; //  720 :   1 - 0x1 -- Background 0x5a
      11'h2D1: dout  = 8'b00000001; //  721 :   1 - 0x1
      11'h2D2: dout  = 8'b00000001; //  722 :   1 - 0x1
      11'h2D3: dout  = 8'b00000001; //  723 :   1 - 0x1
      11'h2D4: dout  = 8'b00000001; //  724 :   1 - 0x1
      11'h2D5: dout  = 8'b00000101; //  725 :   5 - 0x5
      11'h2D6: dout  = 8'b00000001; //  726 :   1 - 0x1
      11'h2D7: dout  = 8'b11111110; //  727 : 254 - 0xfe
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Background 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout  = 8'b11111100; //  732 : 252 - 0xfc
      11'h2DD: dout  = 8'b11111110; //  733 : 254 - 0xfe
      11'h2DE: dout  = 8'b00000111; //  734 :   7 - 0x7
      11'h2DF: dout  = 8'b00000011; //  735 :   3 - 0x3
      11'h2E0: dout  = 8'b00010001; //  736 :  17 - 0x11 -- Background 0x5c
      11'h2E1: dout  = 8'b00111001; //  737 :  57 - 0x39
      11'h2E2: dout  = 8'b00010001; //  738 :  17 - 0x11
      11'h2E3: dout  = 8'b00000001; //  739 :   1 - 0x1
      11'h2E4: dout  = 8'b00000001; //  740 :   1 - 0x1
      11'h2E5: dout  = 8'b00000001; //  741 :   1 - 0x1
      11'h2E6: dout  = 8'b00000001; //  742 :   1 - 0x1
      11'h2E7: dout  = 8'b00000001; //  743 :   1 - 0x1
      11'h2E8: dout  = 8'b11101111; //  744 : 239 - 0xef -- Background 0x5d
      11'h2E9: dout  = 8'b00101000; //  745 :  40 - 0x28
      11'h2EA: dout  = 8'b00101000; //  746 :  40 - 0x28
      11'h2EB: dout  = 8'b00101000; //  747 :  40 - 0x28
      11'h2EC: dout  = 8'b00101000; //  748 :  40 - 0x28
      11'h2ED: dout  = 8'b00101000; //  749 :  40 - 0x28
      11'h2EE: dout  = 8'b11101111; //  750 : 239 - 0xef
      11'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      11'h2F0: dout  = 8'b11111110; //  752 : 254 - 0xfe -- Background 0x5e
      11'h2F1: dout  = 8'b10000010; //  753 : 130 - 0x82
      11'h2F2: dout  = 8'b10000010; //  754 : 130 - 0x82
      11'h2F3: dout  = 8'b10000010; //  755 : 130 - 0x82
      11'h2F4: dout  = 8'b10000010; //  756 : 130 - 0x82
      11'h2F5: dout  = 8'b10000010; //  757 : 130 - 0x82
      11'h2F6: dout  = 8'b11111110; //  758 : 254 - 0xfe
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b10000000; //  760 : 128 - 0x80 -- Background 0x5f
      11'h2F9: dout  = 8'b10000000; //  761 : 128 - 0x80
      11'h2FA: dout  = 8'b10000000; //  762 : 128 - 0x80
      11'h2FB: dout  = 8'b10011000; //  763 : 152 - 0x98
      11'h2FC: dout  = 8'b10011100; //  764 : 156 - 0x9c
      11'h2FD: dout  = 8'b10001100; //  765 : 140 - 0x8c
      11'h2FE: dout  = 8'b10000000; //  766 : 128 - 0x80
      11'h2FF: dout  = 8'b01111111; //  767 : 127 - 0x7f
      11'h300: dout  = 8'b11111111; //  768 : 255 - 0xff -- Background 0x60
      11'h301: dout  = 8'b11111111; //  769 : 255 - 0xff
      11'h302: dout  = 8'b10000011; //  770 : 131 - 0x83
      11'h303: dout  = 8'b11110011; //  771 : 243 - 0xf3
      11'h304: dout  = 8'b11110011; //  772 : 243 - 0xf3
      11'h305: dout  = 8'b11110011; //  773 : 243 - 0xf3
      11'h306: dout  = 8'b11110011; //  774 : 243 - 0xf3
      11'h307: dout  = 8'b11110011; //  775 : 243 - 0xf3
      11'h308: dout  = 8'b11111111; //  776 : 255 - 0xff -- Background 0x61
      11'h309: dout  = 8'b11111111; //  777 : 255 - 0xff
      11'h30A: dout  = 8'b11110000; //  778 : 240 - 0xf0
      11'h30B: dout  = 8'b11110110; //  779 : 246 - 0xf6
      11'h30C: dout  = 8'b11110110; //  780 : 246 - 0xf6
      11'h30D: dout  = 8'b11110110; //  781 : 246 - 0xf6
      11'h30E: dout  = 8'b11110110; //  782 : 246 - 0xf6
      11'h30F: dout  = 8'b11110110; //  783 : 246 - 0xf6
      11'h310: dout  = 8'b11111111; //  784 : 255 - 0xff -- Background 0x62
      11'h311: dout  = 8'b11111111; //  785 : 255 - 0xff
      11'h312: dout  = 8'b00000000; //  786 :   0 - 0x0
      11'h313: dout  = 8'b00000000; //  787 :   0 - 0x0
      11'h314: dout  = 8'b00000000; //  788 :   0 - 0x0
      11'h315: dout  = 8'b00000000; //  789 :   0 - 0x0
      11'h316: dout  = 8'b00000000; //  790 :   0 - 0x0
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b11111111; //  792 : 255 - 0xff -- Background 0x63
      11'h319: dout  = 8'b11111111; //  793 : 255 - 0xff
      11'h31A: dout  = 8'b00000001; //  794 :   1 - 0x1
      11'h31B: dout  = 8'b01010111; //  795 :  87 - 0x57
      11'h31C: dout  = 8'b00101111; //  796 :  47 - 0x2f
      11'h31D: dout  = 8'b01010111; //  797 :  87 - 0x57
      11'h31E: dout  = 8'b00101111; //  798 :  47 - 0x2f
      11'h31F: dout  = 8'b01010111; //  799 :  87 - 0x57
      11'h320: dout  = 8'b11110011; //  800 : 243 - 0xf3 -- Background 0x64
      11'h321: dout  = 8'b11110011; //  801 : 243 - 0xf3
      11'h322: dout  = 8'b11110011; //  802 : 243 - 0xf3
      11'h323: dout  = 8'b11110011; //  803 : 243 - 0xf3
      11'h324: dout  = 8'b11110011; //  804 : 243 - 0xf3
      11'h325: dout  = 8'b11110011; //  805 : 243 - 0xf3
      11'h326: dout  = 8'b11111111; //  806 : 255 - 0xff
      11'h327: dout  = 8'b00111111; //  807 :  63 - 0x3f
      11'h328: dout  = 8'b11110110; //  808 : 246 - 0xf6 -- Background 0x65
      11'h329: dout  = 8'b11110110; //  809 : 246 - 0xf6
      11'h32A: dout  = 8'b11110110; //  810 : 246 - 0xf6
      11'h32B: dout  = 8'b11110110; //  811 : 246 - 0xf6
      11'h32C: dout  = 8'b11110110; //  812 : 246 - 0xf6
      11'h32D: dout  = 8'b11110110; //  813 : 246 - 0xf6
      11'h32E: dout  = 8'b11111111; //  814 : 255 - 0xff
      11'h32F: dout  = 8'b11111111; //  815 : 255 - 0xff
      11'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Background 0x66
      11'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      11'h332: dout  = 8'b00000000; //  818 :   0 - 0x0
      11'h333: dout  = 8'b00000000; //  819 :   0 - 0x0
      11'h334: dout  = 8'b00000000; //  820 :   0 - 0x0
      11'h335: dout  = 8'b00000000; //  821 :   0 - 0x0
      11'h336: dout  = 8'b11111111; //  822 : 255 - 0xff
      11'h337: dout  = 8'b11111111; //  823 : 255 - 0xff
      11'h338: dout  = 8'b00101111; //  824 :  47 - 0x2f -- Background 0x67
      11'h339: dout  = 8'b01010111; //  825 :  87 - 0x57
      11'h33A: dout  = 8'b00101111; //  826 :  47 - 0x2f
      11'h33B: dout  = 8'b01010111; //  827 :  87 - 0x57
      11'h33C: dout  = 8'b00101111; //  828 :  47 - 0x2f
      11'h33D: dout  = 8'b01010111; //  829 :  87 - 0x57
      11'h33E: dout  = 8'b11111111; //  830 : 255 - 0xff
      11'h33F: dout  = 8'b11111100; //  831 : 252 - 0xfc
      11'h340: dout  = 8'b00111100; //  832 :  60 - 0x3c -- Background 0x68
      11'h341: dout  = 8'b00111100; //  833 :  60 - 0x3c
      11'h342: dout  = 8'b00111100; //  834 :  60 - 0x3c
      11'h343: dout  = 8'b00111100; //  835 :  60 - 0x3c
      11'h344: dout  = 8'b00111100; //  836 :  60 - 0x3c
      11'h345: dout  = 8'b00111100; //  837 :  60 - 0x3c
      11'h346: dout  = 8'b00111100; //  838 :  60 - 0x3c
      11'h347: dout  = 8'b00111100; //  839 :  60 - 0x3c
      11'h348: dout  = 8'b11111011; //  840 : 251 - 0xfb -- Background 0x69
      11'h349: dout  = 8'b11111011; //  841 : 251 - 0xfb
      11'h34A: dout  = 8'b11111011; //  842 : 251 - 0xfb
      11'h34B: dout  = 8'b11111011; //  843 : 251 - 0xfb
      11'h34C: dout  = 8'b11111011; //  844 : 251 - 0xfb
      11'h34D: dout  = 8'b11111011; //  845 : 251 - 0xfb
      11'h34E: dout  = 8'b11111011; //  846 : 251 - 0xfb
      11'h34F: dout  = 8'b11111011; //  847 : 251 - 0xfb
      11'h350: dout  = 8'b10111100; //  848 : 188 - 0xbc -- Background 0x6a
      11'h351: dout  = 8'b01011100; //  849 :  92 - 0x5c
      11'h352: dout  = 8'b10111100; //  850 : 188 - 0xbc
      11'h353: dout  = 8'b01011100; //  851 :  92 - 0x5c
      11'h354: dout  = 8'b10111100; //  852 : 188 - 0xbc
      11'h355: dout  = 8'b01011100; //  853 :  92 - 0x5c
      11'h356: dout  = 8'b10111100; //  854 : 188 - 0xbc
      11'h357: dout  = 8'b01011100; //  855 :  92 - 0x5c
      11'h358: dout  = 8'b00011111; //  856 :  31 - 0x1f -- Background 0x6b
      11'h359: dout  = 8'b00100000; //  857 :  32 - 0x20
      11'h35A: dout  = 8'b01000000; //  858 :  64 - 0x40
      11'h35B: dout  = 8'b01000000; //  859 :  64 - 0x40
      11'h35C: dout  = 8'b10000000; //  860 : 128 - 0x80
      11'h35D: dout  = 8'b10000000; //  861 : 128 - 0x80
      11'h35E: dout  = 8'b10000000; //  862 : 128 - 0x80
      11'h35F: dout  = 8'b10000001; //  863 : 129 - 0x81
      11'h360: dout  = 8'b11111111; //  864 : 255 - 0xff -- Background 0x6c
      11'h361: dout  = 8'b10000000; //  865 : 128 - 0x80
      11'h362: dout  = 8'b10000000; //  866 : 128 - 0x80
      11'h363: dout  = 8'b11000000; //  867 : 192 - 0xc0
      11'h364: dout  = 8'b11111111; //  868 : 255 - 0xff
      11'h365: dout  = 8'b11111111; //  869 : 255 - 0xff
      11'h366: dout  = 8'b11111110; //  870 : 254 - 0xfe
      11'h367: dout  = 8'b11111110; //  871 : 254 - 0xfe
      11'h368: dout  = 8'b11111111; //  872 : 255 - 0xff -- Background 0x6d
      11'h369: dout  = 8'b01111111; //  873 : 127 - 0x7f
      11'h36A: dout  = 8'b01111111; //  874 : 127 - 0x7f
      11'h36B: dout  = 8'b11111111; //  875 : 255 - 0xff
      11'h36C: dout  = 8'b11111111; //  876 : 255 - 0xff
      11'h36D: dout  = 8'b00000111; //  877 :   7 - 0x7
      11'h36E: dout  = 8'b00000011; //  878 :   3 - 0x3
      11'h36F: dout  = 8'b00000011; //  879 :   3 - 0x3
      11'h370: dout  = 8'b11111111; //  880 : 255 - 0xff -- Background 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout  = 8'b10000001; //  885 : 129 - 0x81
      11'h376: dout  = 8'b11000011; //  886 : 195 - 0xc3
      11'h377: dout  = 8'b11111111; //  887 : 255 - 0xff
      11'h378: dout  = 8'b11111000; //  888 : 248 - 0xf8 -- Background 0x6f
      11'h379: dout  = 8'b11111100; //  889 : 252 - 0xfc
      11'h37A: dout  = 8'b11111110; //  890 : 254 - 0xfe
      11'h37B: dout  = 8'b11111110; //  891 : 254 - 0xfe
      11'h37C: dout  = 8'b11100011; //  892 : 227 - 0xe3
      11'h37D: dout  = 8'b11000001; //  893 : 193 - 0xc1
      11'h37E: dout  = 8'b10000001; //  894 : 129 - 0x81
      11'h37F: dout  = 8'b10000001; //  895 : 129 - 0x81
      11'h380: dout  = 8'b10000011; //  896 : 131 - 0x83 -- Background 0x70
      11'h381: dout  = 8'b11111111; //  897 : 255 - 0xff
      11'h382: dout  = 8'b11111111; //  898 : 255 - 0xff
      11'h383: dout  = 8'b11111111; //  899 : 255 - 0xff
      11'h384: dout  = 8'b11111111; //  900 : 255 - 0xff
      11'h385: dout  = 8'b11111111; //  901 : 255 - 0xff
      11'h386: dout  = 8'b01111111; //  902 : 127 - 0x7f
      11'h387: dout  = 8'b00011111; //  903 :  31 - 0x1f
      11'h388: dout  = 8'b11111100; //  904 : 252 - 0xfc -- Background 0x71
      11'h389: dout  = 8'b11111100; //  905 : 252 - 0xfc
      11'h38A: dout  = 8'b11111100; //  906 : 252 - 0xfc
      11'h38B: dout  = 8'b11111100; //  907 : 252 - 0xfc
      11'h38C: dout  = 8'b11111110; //  908 : 254 - 0xfe
      11'h38D: dout  = 8'b11111110; //  909 : 254 - 0xfe
      11'h38E: dout  = 8'b11111111; //  910 : 255 - 0xff
      11'h38F: dout  = 8'b11111111; //  911 : 255 - 0xff
      11'h390: dout  = 8'b00000001; //  912 :   1 - 0x1 -- Background 0x72
      11'h391: dout  = 8'b00000001; //  913 :   1 - 0x1
      11'h392: dout  = 8'b00000001; //  914 :   1 - 0x1
      11'h393: dout  = 8'b00000001; //  915 :   1 - 0x1
      11'h394: dout  = 8'b00000011; //  916 :   3 - 0x3
      11'h395: dout  = 8'b00000011; //  917 :   3 - 0x3
      11'h396: dout  = 8'b00000111; //  918 :   7 - 0x7
      11'h397: dout  = 8'b11111111; //  919 : 255 - 0xff
      11'h398: dout  = 8'b11111111; //  920 : 255 - 0xff -- Background 0x73
      11'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout  = 8'b11111111; //  922 : 255 - 0xff
      11'h39B: dout  = 8'b11111111; //  923 : 255 - 0xff
      11'h39C: dout  = 8'b11111111; //  924 : 255 - 0xff
      11'h39D: dout  = 8'b11111111; //  925 : 255 - 0xff
      11'h39E: dout  = 8'b11111111; //  926 : 255 - 0xff
      11'h39F: dout  = 8'b11111111; //  927 : 255 - 0xff
      11'h3A0: dout  = 8'b10000001; //  928 : 129 - 0x81 -- Background 0x74
      11'h3A1: dout  = 8'b11000001; //  929 : 193 - 0xc1
      11'h3A2: dout  = 8'b11100011; //  930 : 227 - 0xe3
      11'h3A3: dout  = 8'b11111111; //  931 : 255 - 0xff
      11'h3A4: dout  = 8'b11111111; //  932 : 255 - 0xff
      11'h3A5: dout  = 8'b11111111; //  933 : 255 - 0xff
      11'h3A6: dout  = 8'b11111111; //  934 : 255 - 0xff
      11'h3A7: dout  = 8'b11111110; //  935 : 254 - 0xfe
      11'h3A8: dout  = 8'b11111111; //  936 : 255 - 0xff -- Background 0x75
      11'h3A9: dout  = 8'b11111111; //  937 : 255 - 0xff
      11'h3AA: dout  = 8'b11111111; //  938 : 255 - 0xff
      11'h3AB: dout  = 8'b11111111; //  939 : 255 - 0xff
      11'h3AC: dout  = 8'b11111111; //  940 : 255 - 0xff
      11'h3AD: dout  = 8'b11111011; //  941 : 251 - 0xfb
      11'h3AE: dout  = 8'b10110101; //  942 : 181 - 0xb5
      11'h3AF: dout  = 8'b11001110; //  943 : 206 - 0xce
      11'h3B0: dout  = 8'b11111111; //  944 : 255 - 0xff -- Background 0x76
      11'h3B1: dout  = 8'b11111111; //  945 : 255 - 0xff
      11'h3B2: dout  = 8'b11111111; //  946 : 255 - 0xff
      11'h3B3: dout  = 8'b11111111; //  947 : 255 - 0xff
      11'h3B4: dout  = 8'b11111111; //  948 : 255 - 0xff
      11'h3B5: dout  = 8'b11011111; //  949 : 223 - 0xdf
      11'h3B6: dout  = 8'b10101101; //  950 : 173 - 0xad
      11'h3B7: dout  = 8'b01110011; //  951 : 115 - 0x73
      11'h3B8: dout  = 8'b01110111; //  952 : 119 - 0x77 -- Background 0x77
      11'h3B9: dout  = 8'b01110111; //  953 : 119 - 0x77
      11'h3BA: dout  = 8'b01110111; //  954 : 119 - 0x77
      11'h3BB: dout  = 8'b01110111; //  955 : 119 - 0x77
      11'h3BC: dout  = 8'b01110111; //  956 : 119 - 0x77
      11'h3BD: dout  = 8'b01110111; //  957 : 119 - 0x77
      11'h3BE: dout  = 8'b01110111; //  958 : 119 - 0x77
      11'h3BF: dout  = 8'b01110111; //  959 : 119 - 0x77
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b11111111; //  967 : 255 - 0xff
      11'h3C8: dout  = 8'b01110111; //  968 : 119 - 0x77 -- Background 0x79
      11'h3C9: dout  = 8'b01110111; //  969 : 119 - 0x77
      11'h3CA: dout  = 8'b01110111; //  970 : 119 - 0x77
      11'h3CB: dout  = 8'b01110111; //  971 : 119 - 0x77
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b00000001; //  976 :   1 - 0x1 -- Background 0x7a
      11'h3D1: dout  = 8'b00000001; //  977 :   1 - 0x1
      11'h3D2: dout  = 8'b00000001; //  978 :   1 - 0x1
      11'h3D3: dout  = 8'b00011001; //  979 :  25 - 0x19
      11'h3D4: dout  = 8'b00011101; //  980 :  29 - 0x1d
      11'h3D5: dout  = 8'b00001101; //  981 :  13 - 0xd
      11'h3D6: dout  = 8'b00000001; //  982 :   1 - 0x1
      11'h3D7: dout  = 8'b11111110; //  983 : 254 - 0xfe
      11'h3D8: dout  = 8'b00100000; //  984 :  32 - 0x20 -- Background 0x7b
      11'h3D9: dout  = 8'b01111000; //  985 : 120 - 0x78
      11'h3DA: dout  = 8'b01111111; //  986 : 127 - 0x7f
      11'h3DB: dout  = 8'b11111110; //  987 : 254 - 0xfe
      11'h3DC: dout  = 8'b11111110; //  988 : 254 - 0xfe
      11'h3DD: dout  = 8'b11111110; //  989 : 254 - 0xfe
      11'h3DE: dout  = 8'b11111110; //  990 : 254 - 0xfe
      11'h3DF: dout  = 8'b11111110; //  991 : 254 - 0xfe
      11'h3E0: dout  = 8'b00000100; //  992 :   4 - 0x4 -- Background 0x7c
      11'h3E1: dout  = 8'b10011010; //  993 : 154 - 0x9a
      11'h3E2: dout  = 8'b11111010; //  994 : 250 - 0xfa
      11'h3E3: dout  = 8'b11111101; //  995 : 253 - 0xfd
      11'h3E4: dout  = 8'b11111101; //  996 : 253 - 0xfd
      11'h3E5: dout  = 8'b11111101; //  997 : 253 - 0xfd
      11'h3E6: dout  = 8'b11111101; //  998 : 253 - 0xfd
      11'h3E7: dout  = 8'b11111101; //  999 : 253 - 0xfd
      11'h3E8: dout  = 8'b01111110; // 1000 : 126 - 0x7e -- Background 0x7d
      11'h3E9: dout  = 8'b00111000; // 1001 :  56 - 0x38
      11'h3EA: dout  = 8'b00100001; // 1002 :  33 - 0x21
      11'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      11'h3EC: dout  = 8'b00000001; // 1004 :   1 - 0x1
      11'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      11'h3EE: dout  = 8'b00000001; // 1006 :   1 - 0x1
      11'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout  = 8'b11111010; // 1008 : 250 - 0xfa -- Background 0x7e
      11'h3F1: dout  = 8'b10001010; // 1009 : 138 - 0x8a
      11'h3F2: dout  = 8'b10000100; // 1010 : 132 - 0x84
      11'h3F3: dout  = 8'b10000000; // 1011 : 128 - 0x80
      11'h3F4: dout  = 8'b10000000; // 1012 : 128 - 0x80
      11'h3F5: dout  = 8'b10000000; // 1013 : 128 - 0x80
      11'h3F6: dout  = 8'b10000000; // 1014 : 128 - 0x80
      11'h3F7: dout  = 8'b10000000; // 1015 : 128 - 0x80
      11'h3F8: dout  = 8'b00000010; // 1016 :   2 - 0x2 -- Background 0x7f
      11'h3F9: dout  = 8'b00000100; // 1017 :   4 - 0x4
      11'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      11'h3FB: dout  = 8'b00010000; // 1019 :  16 - 0x10
      11'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      11'h3FD: dout  = 8'b01000000; // 1021 :  64 - 0x40
      11'h3FE: dout  = 8'b10000000; // 1022 : 128 - 0x80
      11'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      11'h400: dout  = 8'b00001011; // 1024 :  11 - 0xb -- Background 0x80
      11'h401: dout  = 8'b00001011; // 1025 :  11 - 0xb
      11'h402: dout  = 8'b00111011; // 1026 :  59 - 0x3b
      11'h403: dout  = 8'b00001011; // 1027 :  11 - 0xb
      11'h404: dout  = 8'b11111011; // 1028 : 251 - 0xfb
      11'h405: dout  = 8'b00001011; // 1029 :  11 - 0xb
      11'h406: dout  = 8'b00001011; // 1030 :  11 - 0xb
      11'h407: dout  = 8'b00001010; // 1031 :  10 - 0xa
      11'h408: dout  = 8'b10010000; // 1032 : 144 - 0x90 -- Background 0x81
      11'h409: dout  = 8'b00010000; // 1033 :  16 - 0x10
      11'h40A: dout  = 8'b00011111; // 1034 :  31 - 0x1f
      11'h40B: dout  = 8'b00010000; // 1035 :  16 - 0x10
      11'h40C: dout  = 8'b00011111; // 1036 :  31 - 0x1f
      11'h40D: dout  = 8'b00010000; // 1037 :  16 - 0x10
      11'h40E: dout  = 8'b00010000; // 1038 :  16 - 0x10
      11'h40F: dout  = 8'b10010000; // 1039 : 144 - 0x90
      11'h410: dout  = 8'b00111111; // 1040 :  63 - 0x3f -- Background 0x82
      11'h411: dout  = 8'b01111000; // 1041 : 120 - 0x78
      11'h412: dout  = 8'b11100111; // 1042 : 231 - 0xe7
      11'h413: dout  = 8'b11001111; // 1043 : 207 - 0xcf
      11'h414: dout  = 8'b01011000; // 1044 :  88 - 0x58
      11'h415: dout  = 8'b01011000; // 1045 :  88 - 0x58
      11'h416: dout  = 8'b01010000; // 1046 :  80 - 0x50
      11'h417: dout  = 8'b10010000; // 1047 : 144 - 0x90
      11'h418: dout  = 8'b10110000; // 1048 : 176 - 0xb0 -- Background 0x83
      11'h419: dout  = 8'b11111100; // 1049 : 252 - 0xfc
      11'h41A: dout  = 8'b11100010; // 1050 : 226 - 0xe2
      11'h41B: dout  = 8'b11000001; // 1051 : 193 - 0xc1
      11'h41C: dout  = 8'b11000001; // 1052 : 193 - 0xc1
      11'h41D: dout  = 8'b10000011; // 1053 : 131 - 0x83
      11'h41E: dout  = 8'b10001111; // 1054 : 143 - 0x8f
      11'h41F: dout  = 8'b01111110; // 1055 : 126 - 0x7e
      11'h420: dout  = 8'b11111110; // 1056 : 254 - 0xfe -- Background 0x84
      11'h421: dout  = 8'b00000011; // 1057 :   3 - 0x3
      11'h422: dout  = 8'b00001111; // 1058 :  15 - 0xf
      11'h423: dout  = 8'b10010001; // 1059 : 145 - 0x91
      11'h424: dout  = 8'b01110000; // 1060 : 112 - 0x70
      11'h425: dout  = 8'b01100000; // 1061 :  96 - 0x60
      11'h426: dout  = 8'b00100000; // 1062 :  32 - 0x20
      11'h427: dout  = 8'b00110001; // 1063 :  49 - 0x31
      11'h428: dout  = 8'b00111111; // 1064 :  63 - 0x3f -- Background 0x85
      11'h429: dout  = 8'b00111111; // 1065 :  63 - 0x3f
      11'h42A: dout  = 8'b00011101; // 1066 :  29 - 0x1d
      11'h42B: dout  = 8'b00111001; // 1067 :  57 - 0x39
      11'h42C: dout  = 8'b01111011; // 1068 : 123 - 0x7b
      11'h42D: dout  = 8'b11110011; // 1069 : 243 - 0xf3
      11'h42E: dout  = 8'b10000110; // 1070 : 134 - 0x86
      11'h42F: dout  = 8'b11111110; // 1071 : 254 - 0xfe
      11'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Background 0x86
      11'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      11'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      11'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      11'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      11'h435: dout  = 8'b10000000; // 1077 : 128 - 0x80
      11'h436: dout  = 8'b10000000; // 1078 : 128 - 0x80
      11'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      11'h438: dout  = 8'b11111110; // 1080 : 254 - 0xfe -- Background 0x87
      11'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout  = 8'b00000011; // 1085 :   3 - 0x3
      11'h43E: dout  = 8'b00000011; // 1086 :   3 - 0x3
      11'h43F: dout  = 8'b11111111; // 1087 : 255 - 0xff
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x88
      11'h441: dout  = 8'b11111111; // 1089 : 255 - 0xff
      11'h442: dout  = 8'b11111111; // 1090 : 255 - 0xff
      11'h443: dout  = 8'b11111111; // 1091 : 255 - 0xff
      11'h444: dout  = 8'b11111111; // 1092 : 255 - 0xff
      11'h445: dout  = 8'b11111111; // 1093 : 255 - 0xff
      11'h446: dout  = 8'b00000000; // 1094 :   0 - 0x0
      11'h447: dout  = 8'b00000000; // 1095 :   0 - 0x0
      11'h448: dout  = 8'b00111100; // 1096 :  60 - 0x3c -- Background 0x89
      11'h449: dout  = 8'b11111100; // 1097 : 252 - 0xfc
      11'h44A: dout  = 8'b11111100; // 1098 : 252 - 0xfc
      11'h44B: dout  = 8'b11111100; // 1099 : 252 - 0xfc
      11'h44C: dout  = 8'b11111100; // 1100 : 252 - 0xfc
      11'h44D: dout  = 8'b11111100; // 1101 : 252 - 0xfc
      11'h44E: dout  = 8'b00000100; // 1102 :   4 - 0x4
      11'h44F: dout  = 8'b00000100; // 1103 :   4 - 0x4
      11'h450: dout  = 8'b11111111; // 1104 : 255 - 0xff -- Background 0x8a
      11'h451: dout  = 8'b11111111; // 1105 : 255 - 0xff
      11'h452: dout  = 8'b11111111; // 1106 : 255 - 0xff
      11'h453: dout  = 8'b11111111; // 1107 : 255 - 0xff
      11'h454: dout  = 8'b10000000; // 1108 : 128 - 0x80
      11'h455: dout  = 8'b11111111; // 1109 : 255 - 0xff
      11'h456: dout  = 8'b11111111; // 1110 : 255 - 0xff
      11'h457: dout  = 8'b11111111; // 1111 : 255 - 0xff
      11'h458: dout  = 8'b11111111; // 1112 : 255 - 0xff -- Background 0x8b
      11'h459: dout  = 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout  = 8'b11111111; // 1114 : 255 - 0xff
      11'h45B: dout  = 8'b11111111; // 1115 : 255 - 0xff
      11'h45C: dout  = 8'b00000011; // 1116 :   3 - 0x3
      11'h45D: dout  = 8'b11111111; // 1117 : 255 - 0xff
      11'h45E: dout  = 8'b11111111; // 1118 : 255 - 0xff
      11'h45F: dout  = 8'b11111111; // 1119 : 255 - 0xff
      11'h460: dout  = 8'b11111111; // 1120 : 255 - 0xff -- Background 0x8c
      11'h461: dout  = 8'b11111111; // 1121 : 255 - 0xff
      11'h462: dout  = 8'b11111111; // 1122 : 255 - 0xff
      11'h463: dout  = 8'b11111111; // 1123 : 255 - 0xff
      11'h464: dout  = 8'b11111111; // 1124 : 255 - 0xff
      11'h465: dout  = 8'b00000000; // 1125 :   0 - 0x0
      11'h466: dout  = 8'b11111111; // 1126 : 255 - 0xff
      11'h467: dout  = 8'b11111111; // 1127 : 255 - 0xff
      11'h468: dout  = 8'b11111100; // 1128 : 252 - 0xfc -- Background 0x8d
      11'h469: dout  = 8'b11111100; // 1129 : 252 - 0xfc
      11'h46A: dout  = 8'b11111110; // 1130 : 254 - 0xfe
      11'h46B: dout  = 8'b11111110; // 1131 : 254 - 0xfe
      11'h46C: dout  = 8'b11111110; // 1132 : 254 - 0xfe
      11'h46D: dout  = 8'b00000010; // 1133 :   2 - 0x2
      11'h46E: dout  = 8'b11111110; // 1134 : 254 - 0xfe
      11'h46F: dout  = 8'b11111110; // 1135 : 254 - 0xfe
      11'h470: dout  = 8'b11111111; // 1136 : 255 - 0xff -- Background 0x8e
      11'h471: dout  = 8'b10000000; // 1137 : 128 - 0x80
      11'h472: dout  = 8'b10000000; // 1138 : 128 - 0x80
      11'h473: dout  = 8'b10000000; // 1139 : 128 - 0x80
      11'h474: dout  = 8'b10000000; // 1140 : 128 - 0x80
      11'h475: dout  = 8'b10000000; // 1141 : 128 - 0x80
      11'h476: dout  = 8'b10000000; // 1142 : 128 - 0x80
      11'h477: dout  = 8'b10000000; // 1143 : 128 - 0x80
      11'h478: dout  = 8'b11111111; // 1144 : 255 - 0xff -- Background 0x8f
      11'h479: dout  = 8'b00000011; // 1145 :   3 - 0x3
      11'h47A: dout  = 8'b00000011; // 1146 :   3 - 0x3
      11'h47B: dout  = 8'b00000011; // 1147 :   3 - 0x3
      11'h47C: dout  = 8'b00000011; // 1148 :   3 - 0x3
      11'h47D: dout  = 8'b00000011; // 1149 :   3 - 0x3
      11'h47E: dout  = 8'b00000011; // 1150 :   3 - 0x3
      11'h47F: dout  = 8'b00000011; // 1151 :   3 - 0x3
      11'h480: dout  = 8'b00000010; // 1152 :   2 - 0x2 -- Background 0x90
      11'h481: dout  = 8'b00000010; // 1153 :   2 - 0x2
      11'h482: dout  = 8'b00000010; // 1154 :   2 - 0x2
      11'h483: dout  = 8'b00000010; // 1155 :   2 - 0x2
      11'h484: dout  = 8'b00000010; // 1156 :   2 - 0x2
      11'h485: dout  = 8'b00000010; // 1157 :   2 - 0x2
      11'h486: dout  = 8'b00000100; // 1158 :   4 - 0x4
      11'h487: dout  = 8'b00000100; // 1159 :   4 - 0x4
      11'h488: dout  = 8'b10000000; // 1160 : 128 - 0x80 -- Background 0x91
      11'h489: dout  = 8'b10000000; // 1161 : 128 - 0x80
      11'h48A: dout  = 8'b10101010; // 1162 : 170 - 0xaa
      11'h48B: dout  = 8'b11010101; // 1163 : 213 - 0xd5
      11'h48C: dout  = 8'b10101010; // 1164 : 170 - 0xaa
      11'h48D: dout  = 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout  = 8'b11111111; // 1166 : 255 - 0xff
      11'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout  = 8'b00000011; // 1168 :   3 - 0x3 -- Background 0x92
      11'h491: dout  = 8'b00000011; // 1169 :   3 - 0x3
      11'h492: dout  = 8'b10101011; // 1170 : 171 - 0xab
      11'h493: dout  = 8'b01010111; // 1171 :  87 - 0x57
      11'h494: dout  = 8'b10101011; // 1172 : 171 - 0xab
      11'h495: dout  = 8'b11111111; // 1173 : 255 - 0xff
      11'h496: dout  = 8'b11111111; // 1174 : 255 - 0xff
      11'h497: dout  = 8'b11111110; // 1175 : 254 - 0xfe
      11'h498: dout  = 8'b00000000; // 1176 :   0 - 0x0 -- Background 0x93
      11'h499: dout  = 8'b01010101; // 1177 :  85 - 0x55
      11'h49A: dout  = 8'b10101010; // 1178 : 170 - 0xaa
      11'h49B: dout  = 8'b01010101; // 1179 :  85 - 0x55
      11'h49C: dout  = 8'b11111111; // 1180 : 255 - 0xff
      11'h49D: dout  = 8'b11111111; // 1181 : 255 - 0xff
      11'h49E: dout  = 8'b11111111; // 1182 : 255 - 0xff
      11'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout  = 8'b00000100; // 1184 :   4 - 0x4 -- Background 0x94
      11'h4A1: dout  = 8'b01010100; // 1185 :  84 - 0x54
      11'h4A2: dout  = 8'b10101100; // 1186 : 172 - 0xac
      11'h4A3: dout  = 8'b01011100; // 1187 :  92 - 0x5c
      11'h4A4: dout  = 8'b11111100; // 1188 : 252 - 0xfc
      11'h4A5: dout  = 8'b11111100; // 1189 : 252 - 0xfc
      11'h4A6: dout  = 8'b11111100; // 1190 : 252 - 0xfc
      11'h4A7: dout  = 8'b00111100; // 1191 :  60 - 0x3c
      11'h4A8: dout  = 8'b00111111; // 1192 :  63 - 0x3f -- Background 0x95
      11'h4A9: dout  = 8'b00111111; // 1193 :  63 - 0x3f
      11'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      11'h4AB: dout  = 8'b00111111; // 1195 :  63 - 0x3f
      11'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      11'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      11'h4AF: dout  = 8'b11111111; // 1199 : 255 - 0xff
      11'h4B0: dout  = 8'b01111110; // 1200 : 126 - 0x7e -- Background 0x96
      11'h4B1: dout  = 8'b01111100; // 1201 : 124 - 0x7c
      11'h4B2: dout  = 8'b01111100; // 1202 : 124 - 0x7c
      11'h4B3: dout  = 8'b01111000; // 1203 : 120 - 0x78
      11'h4B4: dout  = 8'b00000000; // 1204 :   0 - 0x0
      11'h4B5: dout  = 8'b00000000; // 1205 :   0 - 0x0
      11'h4B6: dout  = 8'b00000000; // 1206 :   0 - 0x0
      11'h4B7: dout  = 8'b11111111; // 1207 : 255 - 0xff
      11'h4B8: dout  = 8'b00011111; // 1208 :  31 - 0x1f -- Background 0x97
      11'h4B9: dout  = 8'b00001111; // 1209 :  15 - 0xf
      11'h4BA: dout  = 8'b00001111; // 1210 :  15 - 0xf
      11'h4BB: dout  = 8'b00000111; // 1211 :   7 - 0x7
      11'h4BC: dout  = 8'b00000000; // 1212 :   0 - 0x0
      11'h4BD: dout  = 8'b00000000; // 1213 :   0 - 0x0
      11'h4BE: dout  = 8'b00000000; // 1214 :   0 - 0x0
      11'h4BF: dout  = 8'b11111111; // 1215 : 255 - 0xff
      11'h4C0: dout  = 8'b11111110; // 1216 : 254 - 0xfe -- Background 0x98
      11'h4C1: dout  = 8'b11111100; // 1217 : 252 - 0xfc
      11'h4C2: dout  = 8'b11111100; // 1218 : 252 - 0xfc
      11'h4C3: dout  = 8'b11111000; // 1219 : 248 - 0xf8
      11'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      11'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      11'h4C6: dout  = 8'b00000000; // 1222 :   0 - 0x0
      11'h4C7: dout  = 8'b11111111; // 1223 : 255 - 0xff
      11'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- Background 0x99
      11'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      11'h4CA: dout  = 8'b00000000; // 1226 :   0 - 0x0
      11'h4CB: dout  = 8'b00000000; // 1227 :   0 - 0x0
      11'h4CC: dout  = 8'b11111111; // 1228 : 255 - 0xff
      11'h4CD: dout  = 8'b11111111; // 1229 : 255 - 0xff
      11'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      11'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout  = 8'b00011000; // 1232 :  24 - 0x18 -- Background 0x9a
      11'h4D1: dout  = 8'b00011000; // 1233 :  24 - 0x18
      11'h4D2: dout  = 8'b00011000; // 1234 :  24 - 0x18
      11'h4D3: dout  = 8'b00011000; // 1235 :  24 - 0x18
      11'h4D4: dout  = 8'b00011000; // 1236 :  24 - 0x18
      11'h4D5: dout  = 8'b00011000; // 1237 :  24 - 0x18
      11'h4D6: dout  = 8'b00011000; // 1238 :  24 - 0x18
      11'h4D7: dout  = 8'b00011000; // 1239 :  24 - 0x18
      11'h4D8: dout  = 8'b00000111; // 1240 :   7 - 0x7 -- Background 0x9b
      11'h4D9: dout  = 8'b00011111; // 1241 :  31 - 0x1f
      11'h4DA: dout  = 8'b00111111; // 1242 :  63 - 0x3f
      11'h4DB: dout  = 8'b11111111; // 1243 : 255 - 0xff
      11'h4DC: dout  = 8'b01111111; // 1244 : 127 - 0x7f
      11'h4DD: dout  = 8'b01111111; // 1245 : 127 - 0x7f
      11'h4DE: dout  = 8'b11111111; // 1246 : 255 - 0xff
      11'h4DF: dout  = 8'b11111111; // 1247 : 255 - 0xff
      11'h4E0: dout  = 8'b11100001; // 1248 : 225 - 0xe1 -- Background 0x9c
      11'h4E1: dout  = 8'b11111001; // 1249 : 249 - 0xf9
      11'h4E2: dout  = 8'b11111101; // 1250 : 253 - 0xfd
      11'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      11'h4E4: dout  = 8'b11111110; // 1252 : 254 - 0xfe
      11'h4E5: dout  = 8'b11111110; // 1253 : 254 - 0xfe
      11'h4E6: dout  = 8'b11111111; // 1254 : 255 - 0xff
      11'h4E7: dout  = 8'b11111111; // 1255 : 255 - 0xff
      11'h4E8: dout  = 8'b11110000; // 1256 : 240 - 0xf0 -- Background 0x9d
      11'h4E9: dout  = 8'b00010000; // 1257 :  16 - 0x10
      11'h4EA: dout  = 8'b00010000; // 1258 :  16 - 0x10
      11'h4EB: dout  = 8'b00010000; // 1259 :  16 - 0x10
      11'h4EC: dout  = 8'b00010000; // 1260 :  16 - 0x10
      11'h4ED: dout  = 8'b00010000; // 1261 :  16 - 0x10
      11'h4EE: dout  = 8'b00010000; // 1262 :  16 - 0x10
      11'h4EF: dout  = 8'b11111111; // 1263 : 255 - 0xff
      11'h4F0: dout  = 8'b00011111; // 1264 :  31 - 0x1f -- Background 0x9e
      11'h4F1: dout  = 8'b00010000; // 1265 :  16 - 0x10
      11'h4F2: dout  = 8'b00010000; // 1266 :  16 - 0x10
      11'h4F3: dout  = 8'b00010000; // 1267 :  16 - 0x10
      11'h4F4: dout  = 8'b00010000; // 1268 :  16 - 0x10
      11'h4F5: dout  = 8'b00010000; // 1269 :  16 - 0x10
      11'h4F6: dout  = 8'b00010000; // 1270 :  16 - 0x10
      11'h4F7: dout  = 8'b11111111; // 1271 : 255 - 0xff
      11'h4F8: dout  = 8'b10010010; // 1272 : 146 - 0x92 -- Background 0x9f
      11'h4F9: dout  = 8'b10010010; // 1273 : 146 - 0x92
      11'h4FA: dout  = 8'b10010010; // 1274 : 146 - 0x92
      11'h4FB: dout  = 8'b11111110; // 1275 : 254 - 0xfe
      11'h4FC: dout  = 8'b11111110; // 1276 : 254 - 0xfe
      11'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00001010; // 1280 :  10 - 0xa -- Background 0xa0
      11'h501: dout  = 8'b00001010; // 1281 :  10 - 0xa
      11'h502: dout  = 8'b00111010; // 1282 :  58 - 0x3a
      11'h503: dout  = 8'b00001010; // 1283 :  10 - 0xa
      11'h504: dout  = 8'b11111011; // 1284 : 251 - 0xfb
      11'h505: dout  = 8'b00001011; // 1285 :  11 - 0xb
      11'h506: dout  = 8'b00001011; // 1286 :  11 - 0xb
      11'h507: dout  = 8'b00001011; // 1287 :  11 - 0xb
      11'h508: dout  = 8'b10010000; // 1288 : 144 - 0x90 -- Background 0xa1
      11'h509: dout  = 8'b10010000; // 1289 : 144 - 0x90
      11'h50A: dout  = 8'b10011111; // 1290 : 159 - 0x9f
      11'h50B: dout  = 8'b10010000; // 1291 : 144 - 0x90
      11'h50C: dout  = 8'b10011111; // 1292 : 159 - 0x9f
      11'h50D: dout  = 8'b10010000; // 1293 : 144 - 0x90
      11'h50E: dout  = 8'b10010000; // 1294 : 144 - 0x90
      11'h50F: dout  = 8'b10010000; // 1295 : 144 - 0x90
      11'h510: dout  = 8'b00000001; // 1296 :   1 - 0x1 -- Background 0xa2
      11'h511: dout  = 8'b00000001; // 1297 :   1 - 0x1
      11'h512: dout  = 8'b00000001; // 1298 :   1 - 0x1
      11'h513: dout  = 8'b00000001; // 1299 :   1 - 0x1
      11'h514: dout  = 8'b00000001; // 1300 :   1 - 0x1
      11'h515: dout  = 8'b00000001; // 1301 :   1 - 0x1
      11'h516: dout  = 8'b00000001; // 1302 :   1 - 0x1
      11'h517: dout  = 8'b00000001; // 1303 :   1 - 0x1
      11'h518: dout  = 8'b10000000; // 1304 : 128 - 0x80 -- Background 0xa3
      11'h519: dout  = 8'b10000000; // 1305 : 128 - 0x80
      11'h51A: dout  = 8'b10000000; // 1306 : 128 - 0x80
      11'h51B: dout  = 8'b10000000; // 1307 : 128 - 0x80
      11'h51C: dout  = 8'b10000000; // 1308 : 128 - 0x80
      11'h51D: dout  = 8'b10000000; // 1309 : 128 - 0x80
      11'h51E: dout  = 8'b10000000; // 1310 : 128 - 0x80
      11'h51F: dout  = 8'b10000000; // 1311 : 128 - 0x80
      11'h520: dout  = 8'b00001000; // 1312 :   8 - 0x8 -- Background 0xa4
      11'h521: dout  = 8'b10001000; // 1313 : 136 - 0x88
      11'h522: dout  = 8'b10010001; // 1314 : 145 - 0x91
      11'h523: dout  = 8'b11010001; // 1315 : 209 - 0xd1
      11'h524: dout  = 8'b01010011; // 1316 :  83 - 0x53
      11'h525: dout  = 8'b01010011; // 1317 :  83 - 0x53
      11'h526: dout  = 8'b01110011; // 1318 : 115 - 0x73
      11'h527: dout  = 8'b00111111; // 1319 :  63 - 0x3f
      11'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Background 0xa5
      11'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout  = 8'b00000111; // 1322 :   7 - 0x7
      11'h52B: dout  = 8'b00001111; // 1323 :  15 - 0xf
      11'h52C: dout  = 8'b00001100; // 1324 :  12 - 0xc
      11'h52D: dout  = 8'b00011011; // 1325 :  27 - 0x1b
      11'h52E: dout  = 8'b00011011; // 1326 :  27 - 0x1b
      11'h52F: dout  = 8'b00011011; // 1327 :  27 - 0x1b
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Background 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b11100000; // 1330 : 224 - 0xe0
      11'h533: dout  = 8'b11110000; // 1331 : 240 - 0xf0
      11'h534: dout  = 8'b11110000; // 1332 : 240 - 0xf0
      11'h535: dout  = 8'b11111000; // 1333 : 248 - 0xf8
      11'h536: dout  = 8'b11111000; // 1334 : 248 - 0xf8
      11'h537: dout  = 8'b11111000; // 1335 : 248 - 0xf8
      11'h538: dout  = 8'b00011011; // 1336 :  27 - 0x1b -- Background 0xa7
      11'h539: dout  = 8'b00011011; // 1337 :  27 - 0x1b
      11'h53A: dout  = 8'b00011011; // 1338 :  27 - 0x1b
      11'h53B: dout  = 8'b00011011; // 1339 :  27 - 0x1b
      11'h53C: dout  = 8'b00011011; // 1340 :  27 - 0x1b
      11'h53D: dout  = 8'b00001111; // 1341 :  15 - 0xf
      11'h53E: dout  = 8'b00001111; // 1342 :  15 - 0xf
      11'h53F: dout  = 8'b00000111; // 1343 :   7 - 0x7
      11'h540: dout  = 8'b11111000; // 1344 : 248 - 0xf8 -- Background 0xa8
      11'h541: dout  = 8'b11111000; // 1345 : 248 - 0xf8
      11'h542: dout  = 8'b11111000; // 1346 : 248 - 0xf8
      11'h543: dout  = 8'b11111000; // 1347 : 248 - 0xf8
      11'h544: dout  = 8'b11111000; // 1348 : 248 - 0xf8
      11'h545: dout  = 8'b11110000; // 1349 : 240 - 0xf0
      11'h546: dout  = 8'b11110000; // 1350 : 240 - 0xf0
      11'h547: dout  = 8'b11100000; // 1351 : 224 - 0xe0
      11'h548: dout  = 8'b11110001; // 1352 : 241 - 0xf1 -- Background 0xa9
      11'h549: dout  = 8'b00010001; // 1353 :  17 - 0x11
      11'h54A: dout  = 8'b00010001; // 1354 :  17 - 0x11
      11'h54B: dout  = 8'b00011111; // 1355 :  31 - 0x1f
      11'h54C: dout  = 8'b00010000; // 1356 :  16 - 0x10
      11'h54D: dout  = 8'b00010000; // 1357 :  16 - 0x10
      11'h54E: dout  = 8'b00010000; // 1358 :  16 - 0x10
      11'h54F: dout  = 8'b11111111; // 1359 : 255 - 0xff
      11'h550: dout  = 8'b00011111; // 1360 :  31 - 0x1f -- Background 0xaa
      11'h551: dout  = 8'b00010000; // 1361 :  16 - 0x10
      11'h552: dout  = 8'b00010000; // 1362 :  16 - 0x10
      11'h553: dout  = 8'b11110000; // 1363 : 240 - 0xf0
      11'h554: dout  = 8'b00010000; // 1364 :  16 - 0x10
      11'h555: dout  = 8'b00010000; // 1365 :  16 - 0x10
      11'h556: dout  = 8'b00010000; // 1366 :  16 - 0x10
      11'h557: dout  = 8'b11111111; // 1367 : 255 - 0xff
      11'h558: dout  = 8'b01111111; // 1368 : 127 - 0x7f -- Background 0xab
      11'h559: dout  = 8'b10111111; // 1369 : 191 - 0xbf
      11'h55A: dout  = 8'b11011111; // 1370 : 223 - 0xdf
      11'h55B: dout  = 8'b11101111; // 1371 : 239 - 0xef
      11'h55C: dout  = 8'b11110000; // 1372 : 240 - 0xf0
      11'h55D: dout  = 8'b11110000; // 1373 : 240 - 0xf0
      11'h55E: dout  = 8'b11110000; // 1374 : 240 - 0xf0
      11'h55F: dout  = 8'b11110000; // 1375 : 240 - 0xf0
      11'h560: dout  = 8'b11110000; // 1376 : 240 - 0xf0 -- Background 0xac
      11'h561: dout  = 8'b11110000; // 1377 : 240 - 0xf0
      11'h562: dout  = 8'b11110000; // 1378 : 240 - 0xf0
      11'h563: dout  = 8'b11110000; // 1379 : 240 - 0xf0
      11'h564: dout  = 8'b11111111; // 1380 : 255 - 0xff
      11'h565: dout  = 8'b11111111; // 1381 : 255 - 0xff
      11'h566: dout  = 8'b11111111; // 1382 : 255 - 0xff
      11'h567: dout  = 8'b11111111; // 1383 : 255 - 0xff
      11'h568: dout  = 8'b11111111; // 1384 : 255 - 0xff -- Background 0xad
      11'h569: dout  = 8'b11111111; // 1385 : 255 - 0xff
      11'h56A: dout  = 8'b11111111; // 1386 : 255 - 0xff
      11'h56B: dout  = 8'b11111111; // 1387 : 255 - 0xff
      11'h56C: dout  = 8'b00001111; // 1388 :  15 - 0xf
      11'h56D: dout  = 8'b00001111; // 1389 :  15 - 0xf
      11'h56E: dout  = 8'b00001111; // 1390 :  15 - 0xf
      11'h56F: dout  = 8'b00001111; // 1391 :  15 - 0xf
      11'h570: dout  = 8'b00001111; // 1392 :  15 - 0xf -- Background 0xae
      11'h571: dout  = 8'b00001111; // 1393 :  15 - 0xf
      11'h572: dout  = 8'b00001111; // 1394 :  15 - 0xf
      11'h573: dout  = 8'b00001111; // 1395 :  15 - 0xf
      11'h574: dout  = 8'b11110111; // 1396 : 247 - 0xf7
      11'h575: dout  = 8'b11111011; // 1397 : 251 - 0xfb
      11'h576: dout  = 8'b11111101; // 1398 : 253 - 0xfd
      11'h577: dout  = 8'b11111110; // 1399 : 254 - 0xfe
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Background 0xaf
      11'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      11'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      11'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      11'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      11'h57E: dout  = 8'b00011000; // 1406 :  24 - 0x18
      11'h57F: dout  = 8'b00011000; // 1407 :  24 - 0x18
      11'h580: dout  = 8'b00011111; // 1408 :  31 - 0x1f -- Background 0xb0
      11'h581: dout  = 8'b00111111; // 1409 :  63 - 0x3f
      11'h582: dout  = 8'b01111111; // 1410 : 127 - 0x7f
      11'h583: dout  = 8'b01111111; // 1411 : 127 - 0x7f
      11'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      11'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      11'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      11'h587: dout  = 8'b11111111; // 1415 : 255 - 0xff
      11'h588: dout  = 8'b11111111; // 1416 : 255 - 0xff -- Background 0xb1
      11'h589: dout  = 8'b11111111; // 1417 : 255 - 0xff
      11'h58A: dout  = 8'b11111111; // 1418 : 255 - 0xff
      11'h58B: dout  = 8'b01111111; // 1419 : 127 - 0x7f
      11'h58C: dout  = 8'b01111111; // 1420 : 127 - 0x7f
      11'h58D: dout  = 8'b01111111; // 1421 : 127 - 0x7f
      11'h58E: dout  = 8'b00111111; // 1422 :  63 - 0x3f
      11'h58F: dout  = 8'b00011110; // 1423 :  30 - 0x1e
      11'h590: dout  = 8'b11111000; // 1424 : 248 - 0xf8 -- Background 0xb2
      11'h591: dout  = 8'b11111100; // 1425 : 252 - 0xfc
      11'h592: dout  = 8'b11111110; // 1426 : 254 - 0xfe
      11'h593: dout  = 8'b11111110; // 1427 : 254 - 0xfe
      11'h594: dout  = 8'b11111110; // 1428 : 254 - 0xfe
      11'h595: dout  = 8'b11111111; // 1429 : 255 - 0xff
      11'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      11'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      11'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff -- Background 0xb3
      11'h599: dout  = 8'b11111111; // 1433 : 255 - 0xff
      11'h59A: dout  = 8'b11111111; // 1434 : 255 - 0xff
      11'h59B: dout  = 8'b11111110; // 1435 : 254 - 0xfe
      11'h59C: dout  = 8'b11111110; // 1436 : 254 - 0xfe
      11'h59D: dout  = 8'b11111110; // 1437 : 254 - 0xfe
      11'h59E: dout  = 8'b11111100; // 1438 : 252 - 0xfc
      11'h59F: dout  = 8'b01111000; // 1439 : 120 - 0x78
      11'h5A0: dout  = 8'b01111111; // 1440 : 127 - 0x7f -- Background 0xb4
      11'h5A1: dout  = 8'b10000000; // 1441 : 128 - 0x80
      11'h5A2: dout  = 8'b10000000; // 1442 : 128 - 0x80
      11'h5A3: dout  = 8'b10000000; // 1443 : 128 - 0x80
      11'h5A4: dout  = 8'b10000000; // 1444 : 128 - 0x80
      11'h5A5: dout  = 8'b10000000; // 1445 : 128 - 0x80
      11'h5A6: dout  = 8'b10000000; // 1446 : 128 - 0x80
      11'h5A7: dout  = 8'b10000000; // 1447 : 128 - 0x80
      11'h5A8: dout  = 8'b11011110; // 1448 : 222 - 0xde -- Background 0xb5
      11'h5A9: dout  = 8'b01100001; // 1449 :  97 - 0x61
      11'h5AA: dout  = 8'b01100001; // 1450 :  97 - 0x61
      11'h5AB: dout  = 8'b01100001; // 1451 :  97 - 0x61
      11'h5AC: dout  = 8'b01110001; // 1452 : 113 - 0x71
      11'h5AD: dout  = 8'b01011110; // 1453 :  94 - 0x5e
      11'h5AE: dout  = 8'b01111111; // 1454 : 127 - 0x7f
      11'h5AF: dout  = 8'b01100001; // 1455 :  97 - 0x61
      11'h5B0: dout  = 8'b10000000; // 1456 : 128 - 0x80 -- Background 0xb6
      11'h5B1: dout  = 8'b10000000; // 1457 : 128 - 0x80
      11'h5B2: dout  = 8'b11000000; // 1458 : 192 - 0xc0
      11'h5B3: dout  = 8'b11110000; // 1459 : 240 - 0xf0
      11'h5B4: dout  = 8'b10111111; // 1460 : 191 - 0xbf
      11'h5B5: dout  = 8'b10001111; // 1461 : 143 - 0x8f
      11'h5B6: dout  = 8'b10000001; // 1462 : 129 - 0x81
      11'h5B7: dout  = 8'b01111110; // 1463 : 126 - 0x7e
      11'h5B8: dout  = 8'b01100001; // 1464 :  97 - 0x61 -- Background 0xb7
      11'h5B9: dout  = 8'b01100001; // 1465 :  97 - 0x61
      11'h5BA: dout  = 8'b11000001; // 1466 : 193 - 0xc1
      11'h5BB: dout  = 8'b11000001; // 1467 : 193 - 0xc1
      11'h5BC: dout  = 8'b10000001; // 1468 : 129 - 0x81
      11'h5BD: dout  = 8'b10000001; // 1469 : 129 - 0x81
      11'h5BE: dout  = 8'b10000011; // 1470 : 131 - 0x83
      11'h5BF: dout  = 8'b11111110; // 1471 : 254 - 0xfe
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Background 0xb8
      11'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      11'h5C2: dout  = 8'b00000011; // 1474 :   3 - 0x3
      11'h5C3: dout  = 8'b00001111; // 1475 :  15 - 0xf
      11'h5C4: dout  = 8'b00011111; // 1476 :  31 - 0x1f
      11'h5C5: dout  = 8'b00111111; // 1477 :  63 - 0x3f
      11'h5C6: dout  = 8'b01111111; // 1478 : 127 - 0x7f
      11'h5C7: dout  = 8'b01111111; // 1479 : 127 - 0x7f
      11'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- Background 0xb9
      11'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      11'h5CA: dout  = 8'b11000000; // 1482 : 192 - 0xc0
      11'h5CB: dout  = 8'b11110000; // 1483 : 240 - 0xf0
      11'h5CC: dout  = 8'b11111000; // 1484 : 248 - 0xf8
      11'h5CD: dout  = 8'b11111100; // 1485 : 252 - 0xfc
      11'h5CE: dout  = 8'b11111110; // 1486 : 254 - 0xfe
      11'h5CF: dout  = 8'b11111110; // 1487 : 254 - 0xfe
      11'h5D0: dout  = 8'b11111111; // 1488 : 255 - 0xff -- Background 0xba
      11'h5D1: dout  = 8'b11111111; // 1489 : 255 - 0xff
      11'h5D2: dout  = 8'b11111111; // 1490 : 255 - 0xff
      11'h5D3: dout  = 8'b11111111; // 1491 : 255 - 0xff
      11'h5D4: dout  = 8'b11111111; // 1492 : 255 - 0xff
      11'h5D5: dout  = 8'b11111111; // 1493 : 255 - 0xff
      11'h5D6: dout  = 8'b11111111; // 1494 : 255 - 0xff
      11'h5D7: dout  = 8'b11111111; // 1495 : 255 - 0xff
      11'h5D8: dout  = 8'b11111111; // 1496 : 255 - 0xff -- Background 0xbb
      11'h5D9: dout  = 8'b11111111; // 1497 : 255 - 0xff
      11'h5DA: dout  = 8'b11111111; // 1498 : 255 - 0xff
      11'h5DB: dout  = 8'b11111111; // 1499 : 255 - 0xff
      11'h5DC: dout  = 8'b11111111; // 1500 : 255 - 0xff
      11'h5DD: dout  = 8'b11111111; // 1501 : 255 - 0xff
      11'h5DE: dout  = 8'b11111111; // 1502 : 255 - 0xff
      11'h5DF: dout  = 8'b11111111; // 1503 : 255 - 0xff
      11'h5E0: dout  = 8'b01111111; // 1504 : 127 - 0x7f -- Background 0xbc
      11'h5E1: dout  = 8'b01111111; // 1505 : 127 - 0x7f
      11'h5E2: dout  = 8'b01111111; // 1506 : 127 - 0x7f
      11'h5E3: dout  = 8'b00111111; // 1507 :  63 - 0x3f
      11'h5E4: dout  = 8'b00111111; // 1508 :  63 - 0x3f
      11'h5E5: dout  = 8'b00011111; // 1509 :  31 - 0x1f
      11'h5E6: dout  = 8'b00001111; // 1510 :  15 - 0xf
      11'h5E7: dout  = 8'b00000111; // 1511 :   7 - 0x7
      11'h5E8: dout  = 8'b11111110; // 1512 : 254 - 0xfe -- Background 0xbd
      11'h5E9: dout  = 8'b11111110; // 1513 : 254 - 0xfe
      11'h5EA: dout  = 8'b11111110; // 1514 : 254 - 0xfe
      11'h5EB: dout  = 8'b11111100; // 1515 : 252 - 0xfc
      11'h5EC: dout  = 8'b11111100; // 1516 : 252 - 0xfc
      11'h5ED: dout  = 8'b11111000; // 1517 : 248 - 0xf8
      11'h5EE: dout  = 8'b11110000; // 1518 : 240 - 0xf0
      11'h5EF: dout  = 8'b11110000; // 1519 : 240 - 0xf0
      11'h5F0: dout  = 8'b00001111; // 1520 :  15 - 0xf -- Background 0xbe
      11'h5F1: dout  = 8'b00001111; // 1521 :  15 - 0xf
      11'h5F2: dout  = 8'b00001111; // 1522 :  15 - 0xf
      11'h5F3: dout  = 8'b00001111; // 1523 :  15 - 0xf
      11'h5F4: dout  = 8'b00001111; // 1524 :  15 - 0xf
      11'h5F5: dout  = 8'b00001111; // 1525 :  15 - 0xf
      11'h5F6: dout  = 8'b00000111; // 1526 :   7 - 0x7
      11'h5F7: dout  = 8'b00001111; // 1527 :  15 - 0xf
      11'h5F8: dout  = 8'b11110000; // 1528 : 240 - 0xf0 -- Background 0xbf
      11'h5F9: dout  = 8'b11110000; // 1529 : 240 - 0xf0
      11'h5FA: dout  = 8'b11110000; // 1530 : 240 - 0xf0
      11'h5FB: dout  = 8'b11110000; // 1531 : 240 - 0xf0
      11'h5FC: dout  = 8'b11110000; // 1532 : 240 - 0xf0
      11'h5FD: dout  = 8'b11110000; // 1533 : 240 - 0xf0
      11'h5FE: dout  = 8'b11100000; // 1534 : 224 - 0xe0
      11'h5FF: dout  = 8'b11110000; // 1535 : 240 - 0xf0
      11'h600: dout  = 8'b10000001; // 1536 : 129 - 0x81 -- Background 0xc0
      11'h601: dout  = 8'b11000001; // 1537 : 193 - 0xc1
      11'h602: dout  = 8'b10100011; // 1538 : 163 - 0xa3
      11'h603: dout  = 8'b10100011; // 1539 : 163 - 0xa3
      11'h604: dout  = 8'b10011101; // 1540 : 157 - 0x9d
      11'h605: dout  = 8'b10000001; // 1541 : 129 - 0x81
      11'h606: dout  = 8'b10000001; // 1542 : 129 - 0x81
      11'h607: dout  = 8'b10000001; // 1543 : 129 - 0x81
      11'h608: dout  = 8'b11100011; // 1544 : 227 - 0xe3 -- Background 0xc1
      11'h609: dout  = 8'b11110111; // 1545 : 247 - 0xf7
      11'h60A: dout  = 8'b11000001; // 1546 : 193 - 0xc1
      11'h60B: dout  = 8'b11000001; // 1547 : 193 - 0xc1
      11'h60C: dout  = 8'b11000001; // 1548 : 193 - 0xc1
      11'h60D: dout  = 8'b11000001; // 1549 : 193 - 0xc1
      11'h60E: dout  = 8'b11110111; // 1550 : 247 - 0xf7
      11'h60F: dout  = 8'b11100011; // 1551 : 227 - 0xe3
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Background 0xc2
      11'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout  = 8'b00000111; // 1554 :   7 - 0x7
      11'h613: dout  = 8'b00001111; // 1555 :  15 - 0xf
      11'h614: dout  = 8'b00001100; // 1556 :  12 - 0xc
      11'h615: dout  = 8'b00011011; // 1557 :  27 - 0x1b
      11'h616: dout  = 8'b00011011; // 1558 :  27 - 0x1b
      11'h617: dout  = 8'b00011011; // 1559 :  27 - 0x1b
      11'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- Background 0xc3
      11'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout  = 8'b11100000; // 1562 : 224 - 0xe0
      11'h61B: dout  = 8'b11110000; // 1563 : 240 - 0xf0
      11'h61C: dout  = 8'b11110000; // 1564 : 240 - 0xf0
      11'h61D: dout  = 8'b11111000; // 1565 : 248 - 0xf8
      11'h61E: dout  = 8'b11111000; // 1566 : 248 - 0xf8
      11'h61F: dout  = 8'b11111000; // 1567 : 248 - 0xf8
      11'h620: dout  = 8'b00011011; // 1568 :  27 - 0x1b -- Background 0xc4
      11'h621: dout  = 8'b00011011; // 1569 :  27 - 0x1b
      11'h622: dout  = 8'b00011011; // 1570 :  27 - 0x1b
      11'h623: dout  = 8'b00011011; // 1571 :  27 - 0x1b
      11'h624: dout  = 8'b00011011; // 1572 :  27 - 0x1b
      11'h625: dout  = 8'b00001111; // 1573 :  15 - 0xf
      11'h626: dout  = 8'b00001111; // 1574 :  15 - 0xf
      11'h627: dout  = 8'b00000111; // 1575 :   7 - 0x7
      11'h628: dout  = 8'b11111000; // 1576 : 248 - 0xf8 -- Background 0xc5
      11'h629: dout  = 8'b11111000; // 1577 : 248 - 0xf8
      11'h62A: dout  = 8'b11111000; // 1578 : 248 - 0xf8
      11'h62B: dout  = 8'b11111000; // 1579 : 248 - 0xf8
      11'h62C: dout  = 8'b11111000; // 1580 : 248 - 0xf8
      11'h62D: dout  = 8'b11110000; // 1581 : 240 - 0xf0
      11'h62E: dout  = 8'b11110000; // 1582 : 240 - 0xf0
      11'h62F: dout  = 8'b11100000; // 1583 : 224 - 0xe0
      11'h630: dout  = 8'b11100000; // 1584 : 224 - 0xe0 -- Background 0xc6
      11'h631: dout  = 8'b11111111; // 1585 : 255 - 0xff
      11'h632: dout  = 8'b11111111; // 1586 : 255 - 0xff
      11'h633: dout  = 8'b11111111; // 1587 : 255 - 0xff
      11'h634: dout  = 8'b11111111; // 1588 : 255 - 0xff
      11'h635: dout  = 8'b11111111; // 1589 : 255 - 0xff
      11'h636: dout  = 8'b11111111; // 1590 : 255 - 0xff
      11'h637: dout  = 8'b11111111; // 1591 : 255 - 0xff
      11'h638: dout  = 8'b00000111; // 1592 :   7 - 0x7 -- Background 0xc7
      11'h639: dout  = 8'b11111111; // 1593 : 255 - 0xff
      11'h63A: dout  = 8'b11111111; // 1594 : 255 - 0xff
      11'h63B: dout  = 8'b11111111; // 1595 : 255 - 0xff
      11'h63C: dout  = 8'b11111111; // 1596 : 255 - 0xff
      11'h63D: dout  = 8'b11111111; // 1597 : 255 - 0xff
      11'h63E: dout  = 8'b11111111; // 1598 : 255 - 0xff
      11'h63F: dout  = 8'b11111111; // 1599 : 255 - 0xff
      11'h640: dout  = 8'b11111111; // 1600 : 255 - 0xff -- Background 0xc8
      11'h641: dout  = 8'b11111111; // 1601 : 255 - 0xff
      11'h642: dout  = 8'b11111111; // 1602 : 255 - 0xff
      11'h643: dout  = 8'b11111111; // 1603 : 255 - 0xff
      11'h644: dout  = 8'b11111111; // 1604 : 255 - 0xff
      11'h645: dout  = 8'b11111110; // 1605 : 254 - 0xfe
      11'h646: dout  = 8'b11111111; // 1606 : 255 - 0xff
      11'h647: dout  = 8'b11101111; // 1607 : 239 - 0xef
      11'h648: dout  = 8'b11111111; // 1608 : 255 - 0xff -- Background 0xc9
      11'h649: dout  = 8'b11011111; // 1609 : 223 - 0xdf
      11'h64A: dout  = 8'b11101111; // 1610 : 239 - 0xef
      11'h64B: dout  = 8'b10101111; // 1611 : 175 - 0xaf
      11'h64C: dout  = 8'b10101111; // 1612 : 175 - 0xaf
      11'h64D: dout  = 8'b01101111; // 1613 : 111 - 0x6f
      11'h64E: dout  = 8'b11101111; // 1614 : 239 - 0xef
      11'h64F: dout  = 8'b11100111; // 1615 : 231 - 0xe7
      11'h650: dout  = 8'b00011111; // 1616 :  31 - 0x1f -- Background 0xca
      11'h651: dout  = 8'b00011111; // 1617 :  31 - 0x1f
      11'h652: dout  = 8'b00111111; // 1618 :  63 - 0x3f
      11'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      11'h654: dout  = 8'b01110000; // 1620 : 112 - 0x70
      11'h655: dout  = 8'b01100011; // 1621 :  99 - 0x63
      11'h656: dout  = 8'b11100111; // 1622 : 231 - 0xe7
      11'h657: dout  = 8'b11100101; // 1623 : 229 - 0xe5
      11'h658: dout  = 8'b11110000; // 1624 : 240 - 0xf0 -- Background 0xcb
      11'h659: dout  = 8'b11110000; // 1625 : 240 - 0xf0
      11'h65A: dout  = 8'b11111000; // 1626 : 248 - 0xf8
      11'h65B: dout  = 8'b11111000; // 1627 : 248 - 0xf8
      11'h65C: dout  = 8'b00001100; // 1628 :  12 - 0xc
      11'h65D: dout  = 8'b11000100; // 1629 : 196 - 0xc4
      11'h65E: dout  = 8'b11100100; // 1630 : 228 - 0xe4
      11'h65F: dout  = 8'b10100110; // 1631 : 166 - 0xa6
      11'h660: dout  = 8'b11101001; // 1632 : 233 - 0xe9 -- Background 0xcc
      11'h661: dout  = 8'b11101001; // 1633 : 233 - 0xe9
      11'h662: dout  = 8'b11101001; // 1634 : 233 - 0xe9
      11'h663: dout  = 8'b11101111; // 1635 : 239 - 0xef
      11'h664: dout  = 8'b11100010; // 1636 : 226 - 0xe2
      11'h665: dout  = 8'b11100011; // 1637 : 227 - 0xe3
      11'h666: dout  = 8'b11110000; // 1638 : 240 - 0xf0
      11'h667: dout  = 8'b11111111; // 1639 : 255 - 0xff
      11'h668: dout  = 8'b10010110; // 1640 : 150 - 0x96 -- Background 0xcd
      11'h669: dout  = 8'b10010110; // 1641 : 150 - 0x96
      11'h66A: dout  = 8'b10010110; // 1642 : 150 - 0x96
      11'h66B: dout  = 8'b11110110; // 1643 : 246 - 0xf6
      11'h66C: dout  = 8'b01000110; // 1644 :  70 - 0x46
      11'h66D: dout  = 8'b11000110; // 1645 : 198 - 0xc6
      11'h66E: dout  = 8'b00001110; // 1646 :  14 - 0xe
      11'h66F: dout  = 8'b11111110; // 1647 : 254 - 0xfe
      11'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Background 0xce
      11'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      11'h676: dout  = 8'b01111110; // 1654 : 126 - 0x7e
      11'h677: dout  = 8'b00111100; // 1655 :  60 - 0x3c
      11'h678: dout  = 8'b00111100; // 1656 :  60 - 0x3c -- Background 0xcf
      11'h679: dout  = 8'b01000010; // 1657 :  66 - 0x42
      11'h67A: dout  = 8'b10011001; // 1658 : 153 - 0x99
      11'h67B: dout  = 8'b10100001; // 1659 : 161 - 0xa1
      11'h67C: dout  = 8'b10100001; // 1660 : 161 - 0xa1
      11'h67D: dout  = 8'b10011001; // 1661 : 153 - 0x99
      11'h67E: dout  = 8'b01000010; // 1662 :  66 - 0x42
      11'h67F: dout  = 8'b00111100; // 1663 :  60 - 0x3c
      11'h680: dout  = 8'b00001111; // 1664 :  15 - 0xf -- Background 0xd0
      11'h681: dout  = 8'b00011111; // 1665 :  31 - 0x1f
      11'h682: dout  = 8'b00011111; // 1666 :  31 - 0x1f
      11'h683: dout  = 8'b00111111; // 1667 :  63 - 0x3f
      11'h684: dout  = 8'b00111111; // 1668 :  63 - 0x3f
      11'h685: dout  = 8'b01111111; // 1669 : 127 - 0x7f
      11'h686: dout  = 8'b01111111; // 1670 : 127 - 0x7f
      11'h687: dout  = 8'b01111111; // 1671 : 127 - 0x7f
      11'h688: dout  = 8'b11110000; // 1672 : 240 - 0xf0 -- Background 0xd1
      11'h689: dout  = 8'b11111000; // 1673 : 248 - 0xf8
      11'h68A: dout  = 8'b11111000; // 1674 : 248 - 0xf8
      11'h68B: dout  = 8'b11111100; // 1675 : 252 - 0xfc
      11'h68C: dout  = 8'b11111100; // 1676 : 252 - 0xfc
      11'h68D: dout  = 8'b11111110; // 1677 : 254 - 0xfe
      11'h68E: dout  = 8'b11111110; // 1678 : 254 - 0xfe
      11'h68F: dout  = 8'b11111110; // 1679 : 254 - 0xfe
      11'h690: dout  = 8'b01111111; // 1680 : 127 - 0x7f -- Background 0xd2
      11'h691: dout  = 8'b01111111; // 1681 : 127 - 0x7f
      11'h692: dout  = 8'b00111111; // 1682 :  63 - 0x3f
      11'h693: dout  = 8'b00111111; // 1683 :  63 - 0x3f
      11'h694: dout  = 8'b00111111; // 1684 :  63 - 0x3f
      11'h695: dout  = 8'b00111111; // 1685 :  63 - 0x3f
      11'h696: dout  = 8'b00011111; // 1686 :  31 - 0x1f
      11'h697: dout  = 8'b00011111; // 1687 :  31 - 0x1f
      11'h698: dout  = 8'b11111110; // 1688 : 254 - 0xfe -- Background 0xd3
      11'h699: dout  = 8'b11111111; // 1689 : 255 - 0xff
      11'h69A: dout  = 8'b11111111; // 1690 : 255 - 0xff
      11'h69B: dout  = 8'b11111111; // 1691 : 255 - 0xff
      11'h69C: dout  = 8'b11111100; // 1692 : 252 - 0xfc
      11'h69D: dout  = 8'b11111100; // 1693 : 252 - 0xfc
      11'h69E: dout  = 8'b11111110; // 1694 : 254 - 0xfe
      11'h69F: dout  = 8'b11111110; // 1695 : 254 - 0xfe
      11'h6A0: dout  = 8'b01111111; // 1696 : 127 - 0x7f -- Background 0xd4
      11'h6A1: dout  = 8'b01111111; // 1697 : 127 - 0x7f
      11'h6A2: dout  = 8'b01111111; // 1698 : 127 - 0x7f
      11'h6A3: dout  = 8'b00111111; // 1699 :  63 - 0x3f
      11'h6A4: dout  = 8'b00111111; // 1700 :  63 - 0x3f
      11'h6A5: dout  = 8'b00111111; // 1701 :  63 - 0x3f
      11'h6A6: dout  = 8'b00111111; // 1702 :  63 - 0x3f
      11'h6A7: dout  = 8'b00011111; // 1703 :  31 - 0x1f
      11'h6A8: dout  = 8'b11111110; // 1704 : 254 - 0xfe -- Background 0xd5
      11'h6A9: dout  = 8'b11111110; // 1705 : 254 - 0xfe
      11'h6AA: dout  = 8'b11111111; // 1706 : 255 - 0xff
      11'h6AB: dout  = 8'b11111111; // 1707 : 255 - 0xff
      11'h6AC: dout  = 8'b11111111; // 1708 : 255 - 0xff
      11'h6AD: dout  = 8'b11111111; // 1709 : 255 - 0xff
      11'h6AE: dout  = 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout  = 8'b11111110; // 1711 : 254 - 0xfe
      11'h6B0: dout  = 8'b00011111; // 1712 :  31 - 0x1f -- Background 0xd6
      11'h6B1: dout  = 8'b00001111; // 1713 :  15 - 0xf
      11'h6B2: dout  = 8'b00001111; // 1714 :  15 - 0xf
      11'h6B3: dout  = 8'b00000111; // 1715 :   7 - 0x7
      11'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      11'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      11'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      11'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      11'h6B8: dout  = 8'b11111110; // 1720 : 254 - 0xfe -- Background 0xd7
      11'h6B9: dout  = 8'b11111100; // 1721 : 252 - 0xfc
      11'h6BA: dout  = 8'b11111100; // 1722 : 252 - 0xfc
      11'h6BB: dout  = 8'b11111000; // 1723 : 248 - 0xf8
      11'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      11'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      11'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      11'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout  = 8'b01111110; // 1728 : 126 - 0x7e -- Background 0xd8
      11'h6C1: dout  = 8'b01111110; // 1729 : 126 - 0x7e
      11'h6C2: dout  = 8'b01111110; // 1730 : 126 - 0x7e
      11'h6C3: dout  = 8'b01111110; // 1731 : 126 - 0x7e
      11'h6C4: dout  = 8'b01111111; // 1732 : 127 - 0x7f
      11'h6C5: dout  = 8'b01111111; // 1733 : 127 - 0x7f
      11'h6C6: dout  = 8'b01111111; // 1734 : 127 - 0x7f
      11'h6C7: dout  = 8'b01111111; // 1735 : 127 - 0x7f
      11'h6C8: dout  = 8'b11111111; // 1736 : 255 - 0xff -- Background 0xd9
      11'h6C9: dout  = 8'b11111111; // 1737 : 255 - 0xff
      11'h6CA: dout  = 8'b11111111; // 1738 : 255 - 0xff
      11'h6CB: dout  = 8'b11111111; // 1739 : 255 - 0xff
      11'h6CC: dout  = 8'b11111111; // 1740 : 255 - 0xff
      11'h6CD: dout  = 8'b11111111; // 1741 : 255 - 0xff
      11'h6CE: dout  = 8'b11111111; // 1742 : 255 - 0xff
      11'h6CF: dout  = 8'b11111110; // 1743 : 254 - 0xfe
      11'h6D0: dout  = 8'b11111110; // 1744 : 254 - 0xfe -- Background 0xda
      11'h6D1: dout  = 8'b11111110; // 1745 : 254 - 0xfe
      11'h6D2: dout  = 8'b11111110; // 1746 : 254 - 0xfe
      11'h6D3: dout  = 8'b11111110; // 1747 : 254 - 0xfe
      11'h6D4: dout  = 8'b11111111; // 1748 : 255 - 0xff
      11'h6D5: dout  = 8'b11111111; // 1749 : 255 - 0xff
      11'h6D6: dout  = 8'b11111111; // 1750 : 255 - 0xff
      11'h6D7: dout  = 8'b11111111; // 1751 : 255 - 0xff
      11'h6D8: dout  = 8'b01111111; // 1752 : 127 - 0x7f -- Background 0xdb
      11'h6D9: dout  = 8'b01111111; // 1753 : 127 - 0x7f
      11'h6DA: dout  = 8'b01111111; // 1754 : 127 - 0x7f
      11'h6DB: dout  = 8'b01111111; // 1755 : 127 - 0x7f
      11'h6DC: dout  = 8'b01111111; // 1756 : 127 - 0x7f
      11'h6DD: dout  = 8'b01111111; // 1757 : 127 - 0x7f
      11'h6DE: dout  = 8'b01111111; // 1758 : 127 - 0x7f
      11'h6DF: dout  = 8'b01111111; // 1759 : 127 - 0x7f
      11'h6E0: dout  = 8'b11111111; // 1760 : 255 - 0xff -- Background 0xdc
      11'h6E1: dout  = 8'b11111111; // 1761 : 255 - 0xff
      11'h6E2: dout  = 8'b11111111; // 1762 : 255 - 0xff
      11'h6E3: dout  = 8'b11111111; // 1763 : 255 - 0xff
      11'h6E4: dout  = 8'b11111100; // 1764 : 252 - 0xfc
      11'h6E5: dout  = 8'b11111110; // 1765 : 254 - 0xfe
      11'h6E6: dout  = 8'b11111110; // 1766 : 254 - 0xfe
      11'h6E7: dout  = 8'b01111110; // 1767 : 126 - 0x7e
      11'h6E8: dout  = 8'b11111111; // 1768 : 255 - 0xff -- Background 0xdd
      11'h6E9: dout  = 8'b11111111; // 1769 : 255 - 0xff
      11'h6EA: dout  = 8'b11111111; // 1770 : 255 - 0xff
      11'h6EB: dout  = 8'b11111111; // 1771 : 255 - 0xff
      11'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      11'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      11'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      11'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout  = 8'b01111111; // 1776 : 127 - 0x7f -- Background 0xde
      11'h6F1: dout  = 8'b01111111; // 1777 : 127 - 0x7f
      11'h6F2: dout  = 8'b01111111; // 1778 : 127 - 0x7f
      11'h6F3: dout  = 8'b01111111; // 1779 : 127 - 0x7f
      11'h6F4: dout  = 8'b01111111; // 1780 : 127 - 0x7f
      11'h6F5: dout  = 8'b01111111; // 1781 : 127 - 0x7f
      11'h6F6: dout  = 8'b01111111; // 1782 : 127 - 0x7f
      11'h6F7: dout  = 8'b01111111; // 1783 : 127 - 0x7f
      11'h6F8: dout  = 8'b11111111; // 1784 : 255 - 0xff -- Background 0xdf
      11'h6F9: dout  = 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout  = 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout  = 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout  = 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout  = 8'b11111110; // 1791 : 254 - 0xfe
      11'h700: dout  = 8'b01111110; // 1792 : 126 - 0x7e -- Background 0xe0
      11'h701: dout  = 8'b01111110; // 1793 : 126 - 0x7e
      11'h702: dout  = 8'b01111111; // 1794 : 127 - 0x7f
      11'h703: dout  = 8'b01111111; // 1795 : 127 - 0x7f
      11'h704: dout  = 8'b01111111; // 1796 : 127 - 0x7f
      11'h705: dout  = 8'b01111111; // 1797 : 127 - 0x7f
      11'h706: dout  = 8'b01111111; // 1798 : 127 - 0x7f
      11'h707: dout  = 8'b01111111; // 1799 : 127 - 0x7f
      11'h708: dout  = 8'b00111111; // 1800 :  63 - 0x3f -- Background 0xe1
      11'h709: dout  = 8'b00111111; // 1801 :  63 - 0x3f
      11'h70A: dout  = 8'b00111111; // 1802 :  63 - 0x3f
      11'h70B: dout  = 8'b00111111; // 1803 :  63 - 0x3f
      11'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      11'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout  = 8'b01111110; // 1808 : 126 - 0x7e -- Background 0xe2
      11'h711: dout  = 8'b01111100; // 1809 : 124 - 0x7c
      11'h712: dout  = 8'b01111100; // 1810 : 124 - 0x7c
      11'h713: dout  = 8'b01111000; // 1811 : 120 - 0x78
      11'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      11'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout  = 8'b11111110; // 1816 : 254 - 0xfe -- Background 0xe3
      11'h719: dout  = 8'b11111110; // 1817 : 254 - 0xfe
      11'h71A: dout  = 8'b11111111; // 1818 : 255 - 0xff
      11'h71B: dout  = 8'b11111111; // 1819 : 255 - 0xff
      11'h71C: dout  = 8'b01111111; // 1820 : 127 - 0x7f
      11'h71D: dout  = 8'b01111111; // 1821 : 127 - 0x7f
      11'h71E: dout  = 8'b01111111; // 1822 : 127 - 0x7f
      11'h71F: dout  = 8'b01111111; // 1823 : 127 - 0x7f
      11'h720: dout  = 8'b01111111; // 1824 : 127 - 0x7f -- Background 0xe4
      11'h721: dout  = 8'b01111111; // 1825 : 127 - 0x7f
      11'h722: dout  = 8'b00111111; // 1826 :  63 - 0x3f
      11'h723: dout  = 8'b00111111; // 1827 :  63 - 0x3f
      11'h724: dout  = 8'b00111111; // 1828 :  63 - 0x3f
      11'h725: dout  = 8'b00111111; // 1829 :  63 - 0x3f
      11'h726: dout  = 8'b00011111; // 1830 :  31 - 0x1f
      11'h727: dout  = 8'b00011111; // 1831 :  31 - 0x1f
      11'h728: dout  = 8'b00111111; // 1832 :  63 - 0x3f -- Background 0xe5
      11'h729: dout  = 8'b10111111; // 1833 : 191 - 0xbf
      11'h72A: dout  = 8'b11111111; // 1834 : 255 - 0xff
      11'h72B: dout  = 8'b11111111; // 1835 : 255 - 0xff
      11'h72C: dout  = 8'b11111100; // 1836 : 252 - 0xfc
      11'h72D: dout  = 8'b11111100; // 1837 : 252 - 0xfc
      11'h72E: dout  = 8'b11111110; // 1838 : 254 - 0xfe
      11'h72F: dout  = 8'b11111110; // 1839 : 254 - 0xfe
      11'h730: dout  = 8'b01111111; // 1840 : 127 - 0x7f -- Background 0xe6
      11'h731: dout  = 8'b01111111; // 1841 : 127 - 0x7f
      11'h732: dout  = 8'b01111110; // 1842 : 126 - 0x7e
      11'h733: dout  = 8'b01111110; // 1843 : 126 - 0x7e
      11'h734: dout  = 8'b01111111; // 1844 : 127 - 0x7f
      11'h735: dout  = 8'b01111111; // 1845 : 127 - 0x7f
      11'h736: dout  = 8'b01111111; // 1846 : 127 - 0x7f
      11'h737: dout  = 8'b01111111; // 1847 : 127 - 0x7f
      11'h738: dout  = 8'b01111110; // 1848 : 126 - 0x7e -- Background 0xe7
      11'h739: dout  = 8'b01111110; // 1849 : 126 - 0x7e
      11'h73A: dout  = 8'b01111110; // 1850 : 126 - 0x7e
      11'h73B: dout  = 8'b01111110; // 1851 : 126 - 0x7e
      11'h73C: dout  = 8'b01111111; // 1852 : 127 - 0x7f
      11'h73D: dout  = 8'b01111111; // 1853 : 127 - 0x7f
      11'h73E: dout  = 8'b01111111; // 1854 : 127 - 0x7f
      11'h73F: dout  = 8'b01111111; // 1855 : 127 - 0x7f
      11'h740: dout  = 8'b10000001; // 1856 : 129 - 0x81 -- Background 0xe8
      11'h741: dout  = 8'b11000011; // 1857 : 195 - 0xc3
      11'h742: dout  = 8'b11000011; // 1858 : 195 - 0xc3
      11'h743: dout  = 8'b11100111; // 1859 : 231 - 0xe7
      11'h744: dout  = 8'b11100111; // 1860 : 231 - 0xe7
      11'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout  = 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout  = 8'b00001111; // 1864 :  15 - 0xf -- Background 0xe9
      11'h749: dout  = 8'b01000011; // 1865 :  67 - 0x43
      11'h74A: dout  = 8'b01011011; // 1866 :  91 - 0x5b
      11'h74B: dout  = 8'b01010011; // 1867 :  83 - 0x53
      11'h74C: dout  = 8'b00110001; // 1868 :  49 - 0x31
      11'h74D: dout  = 8'b00011001; // 1869 :  25 - 0x19
      11'h74E: dout  = 8'b00001111; // 1870 :  15 - 0xf
      11'h74F: dout  = 8'b00000111; // 1871 :   7 - 0x7
      11'h750: dout  = 8'b11000001; // 1872 : 193 - 0xc1 -- Background 0xea
      11'h751: dout  = 8'b11000011; // 1873 : 195 - 0xc3
      11'h752: dout  = 8'b11000110; // 1874 : 198 - 0xc6
      11'h753: dout  = 8'b10000100; // 1875 : 132 - 0x84
      11'h754: dout  = 8'b11111100; // 1876 : 252 - 0xfc
      11'h755: dout  = 8'b11111100; // 1877 : 252 - 0xfc
      11'h756: dout  = 8'b00001110; // 1878 :  14 - 0xe
      11'h757: dout  = 8'b00000010; // 1879 :   2 - 0x2
      11'h758: dout  = 8'b00010000; // 1880 :  16 - 0x10 -- Background 0xeb
      11'h759: dout  = 8'b00100000; // 1881 :  32 - 0x20
      11'h75A: dout  = 8'b00100010; // 1882 :  34 - 0x22
      11'h75B: dout  = 8'b10111010; // 1883 : 186 - 0xba
      11'h75C: dout  = 8'b11100110; // 1884 : 230 - 0xe6
      11'h75D: dout  = 8'b11100001; // 1885 : 225 - 0xe1
      11'h75E: dout  = 8'b11000000; // 1886 : 192 - 0xc0
      11'h75F: dout  = 8'b11000000; // 1887 : 192 - 0xc0
      11'h760: dout  = 8'b00100000; // 1888 :  32 - 0x20 -- Background 0xec
      11'h761: dout  = 8'b10100110; // 1889 : 166 - 0xa6
      11'h762: dout  = 8'b01010100; // 1890 :  84 - 0x54
      11'h763: dout  = 8'b00100110; // 1891 :  38 - 0x26
      11'h764: dout  = 8'b00100000; // 1892 :  32 - 0x20
      11'h765: dout  = 8'b11000110; // 1893 : 198 - 0xc6
      11'h766: dout  = 8'b01010100; // 1894 :  84 - 0x54
      11'h767: dout  = 8'b00100110; // 1895 :  38 - 0x26
      11'h768: dout  = 8'b00100000; // 1896 :  32 - 0x20 -- Background 0xed
      11'h769: dout  = 8'b10000101; // 1897 : 133 - 0x85
      11'h76A: dout  = 8'b00000001; // 1898 :   1 - 0x1
      11'h76B: dout  = 8'b01000100; // 1899 :  68 - 0x44
      11'h76C: dout  = 8'b00100000; // 1900 :  32 - 0x20
      11'h76D: dout  = 8'b10000110; // 1901 : 134 - 0x86
      11'h76E: dout  = 8'b01010100; // 1902 :  84 - 0x54
      11'h76F: dout  = 8'b01001000; // 1903 :  72 - 0x48
      11'h770: dout  = 8'b00100000; // 1904 :  32 - 0x20 -- Background 0xee
      11'h771: dout  = 8'b10111010; // 1905 : 186 - 0xba
      11'h772: dout  = 8'b11001001; // 1906 : 201 - 0xc9
      11'h773: dout  = 8'b01001010; // 1907 :  74 - 0x4a
      11'h774: dout  = 8'b00100000; // 1908 :  32 - 0x20
      11'h775: dout  = 8'b10100110; // 1909 : 166 - 0xa6
      11'h776: dout  = 8'b00001010; // 1910 :  10 - 0xa
      11'h777: dout  = 8'b11010000; // 1911 : 208 - 0xd0
      11'h778: dout  = 8'b11010001; // 1912 : 209 - 0xd1 -- Background 0xef
      11'h779: dout  = 8'b00100000; // 1913 :  32 - 0x20
      11'h77A: dout  = 8'b11000110; // 1914 : 198 - 0xc6
      11'h77B: dout  = 8'b00001010; // 1915 :  10 - 0xa
      11'h77C: dout  = 8'b11010010; // 1916 : 210 - 0xd2
      11'h77D: dout  = 8'b11010011; // 1917 : 211 - 0xd3
      11'h77E: dout  = 8'b11011011; // 1918 : 219 - 0xdb
      11'h77F: dout  = 8'b11011011; // 1919 : 219 - 0xdb
      11'h780: dout  = 8'b00001010; // 1920 :  10 - 0xa -- Background 0xf0
      11'h781: dout  = 8'b11010100; // 1921 : 212 - 0xd4
      11'h782: dout  = 8'b11010101; // 1922 : 213 - 0xd5
      11'h783: dout  = 8'b11010100; // 1923 : 212 - 0xd4
      11'h784: dout  = 8'b11011001; // 1924 : 217 - 0xd9
      11'h785: dout  = 8'b11011011; // 1925 : 219 - 0xdb
      11'h786: dout  = 8'b11100010; // 1926 : 226 - 0xe2
      11'h787: dout  = 8'b11010100; // 1927 : 212 - 0xd4
      11'h788: dout  = 8'b11010110; // 1928 : 214 - 0xd6 -- Background 0xf1
      11'h789: dout  = 8'b11010111; // 1929 : 215 - 0xd7
      11'h78A: dout  = 8'b11100001; // 1930 : 225 - 0xe1
      11'h78B: dout  = 8'b00100110; // 1931 :  38 - 0x26
      11'h78C: dout  = 8'b11010110; // 1932 : 214 - 0xd6
      11'h78D: dout  = 8'b11011101; // 1933 : 221 - 0xdd
      11'h78E: dout  = 8'b11100001; // 1934 : 225 - 0xe1
      11'h78F: dout  = 8'b11100001; // 1935 : 225 - 0xe1
      11'h790: dout  = 8'b11011110; // 1936 : 222 - 0xde -- Background 0xf2
      11'h791: dout  = 8'b11010001; // 1937 : 209 - 0xd1
      11'h792: dout  = 8'b11011000; // 1938 : 216 - 0xd8
      11'h793: dout  = 8'b11010000; // 1939 : 208 - 0xd0
      11'h794: dout  = 8'b11010001; // 1940 : 209 - 0xd1
      11'h795: dout  = 8'b00100110; // 1941 :  38 - 0x26
      11'h796: dout  = 8'b11011110; // 1942 : 222 - 0xde
      11'h797: dout  = 8'b11010001; // 1943 : 209 - 0xd1
      11'h798: dout  = 8'b01000110; // 1944 :  70 - 0x46 -- Background 0xf3
      11'h799: dout  = 8'b00010100; // 1945 :  20 - 0x14
      11'h79A: dout  = 8'b11011011; // 1946 : 219 - 0xdb
      11'h79B: dout  = 8'b01000010; // 1947 :  66 - 0x42
      11'h79C: dout  = 8'b01000010; // 1948 :  66 - 0x42
      11'h79D: dout  = 8'b11011011; // 1949 : 219 - 0xdb
      11'h79E: dout  = 8'b01000010; // 1950 :  66 - 0x42
      11'h79F: dout  = 8'b11011011; // 1951 : 219 - 0xdb
      11'h7A0: dout  = 8'b01000010; // 1952 :  66 - 0x42 -- Background 0xf4
      11'h7A1: dout  = 8'b11011011; // 1953 : 219 - 0xdb
      11'h7A2: dout  = 8'b01000010; // 1954 :  66 - 0x42
      11'h7A3: dout  = 8'b11011011; // 1955 : 219 - 0xdb
      11'h7A4: dout  = 8'b01000010; // 1956 :  66 - 0x42
      11'h7A5: dout  = 8'b00100110; // 1957 :  38 - 0x26
      11'h7A6: dout  = 8'b00100001; // 1958 :  33 - 0x21
      11'h7A7: dout  = 8'b01100110; // 1959 : 102 - 0x66
      11'h7A8: dout  = 8'b11011011; // 1960 : 219 - 0xdb -- Background 0xf5
      11'h7A9: dout  = 8'b00100110; // 1961 :  38 - 0x26
      11'h7AA: dout  = 8'b11011011; // 1962 : 219 - 0xdb
      11'h7AB: dout  = 8'b11011111; // 1963 : 223 - 0xdf
      11'h7AC: dout  = 8'b11011011; // 1964 : 219 - 0xdb
      11'h7AD: dout  = 8'b11011111; // 1965 : 223 - 0xdf
      11'h7AE: dout  = 8'b11011011; // 1966 : 219 - 0xdb
      11'h7AF: dout  = 8'b11011011; // 1967 : 219 - 0xdb
      11'h7B0: dout  = 8'b11011011; // 1968 : 219 - 0xdb -- Background 0xf6
      11'h7B1: dout  = 8'b11011110; // 1969 : 222 - 0xde
      11'h7B2: dout  = 8'b01000011; // 1970 :  67 - 0x43
      11'h7B3: dout  = 8'b11011011; // 1971 : 219 - 0xdb
      11'h7B4: dout  = 8'b11100000; // 1972 : 224 - 0xe0
      11'h7B5: dout  = 8'b11011011; // 1973 : 219 - 0xdb
      11'h7B6: dout  = 8'b11011011; // 1974 : 219 - 0xdb
      11'h7B7: dout  = 8'b11011011; // 1975 : 219 - 0xdb
      11'h7B8: dout  = 8'b11100011; // 1976 : 227 - 0xe3 -- Background 0xf7
      11'h7B9: dout  = 8'b00100110; // 1977 :  38 - 0x26
      11'h7BA: dout  = 8'b00100001; // 1978 :  33 - 0x21
      11'h7BB: dout  = 8'b10100110; // 1979 : 166 - 0xa6
      11'h7BC: dout  = 8'b00010100; // 1980 :  20 - 0x14
      11'h7BD: dout  = 8'b11011011; // 1981 : 219 - 0xdb
      11'h7BE: dout  = 8'b11011011; // 1982 : 219 - 0xdb
      11'h7BF: dout  = 8'b11011011; // 1983 : 219 - 0xdb
      11'h7C0: dout  = 8'b11011011; // 1984 : 219 - 0xdb -- Background 0xf8
      11'h7C1: dout  = 8'b11011001; // 1985 : 217 - 0xd9
      11'h7C2: dout  = 8'b11011011; // 1986 : 219 - 0xdb
      11'h7C3: dout  = 8'b11011011; // 1987 : 219 - 0xdb
      11'h7C4: dout  = 8'b11010100; // 1988 : 212 - 0xd4
      11'h7C5: dout  = 8'b11011001; // 1989 : 217 - 0xd9
      11'h7C6: dout  = 8'b11010100; // 1990 : 212 - 0xd4
      11'h7C7: dout  = 8'b11011001; // 1991 : 217 - 0xd9
      11'h7C8: dout  = 8'b10010101; // 1992 : 149 - 0x95 -- Background 0xf9
      11'h7C9: dout  = 8'b10010101; // 1993 : 149 - 0x95
      11'h7CA: dout  = 8'b10010101; // 1994 : 149 - 0x95
      11'h7CB: dout  = 8'b10010101; // 1995 : 149 - 0x95
      11'h7CC: dout  = 8'b10010101; // 1996 : 149 - 0x95
      11'h7CD: dout  = 8'b10010111; // 1997 : 151 - 0x97
      11'h7CE: dout  = 8'b10011000; // 1998 : 152 - 0x98
      11'h7CF: dout  = 8'b01111000; // 1999 : 120 - 0x78
      11'h7D0: dout  = 8'b10010101; // 2000 : 149 - 0x95 -- Background 0xfa
      11'h7D1: dout  = 8'b01111010; // 2001 : 122 - 0x7a
      11'h7D2: dout  = 8'b00100001; // 2002 :  33 - 0x21
      11'h7D3: dout  = 8'b11101101; // 2003 : 237 - 0xed
      11'h7D4: dout  = 8'b00001110; // 2004 :  14 - 0xe
      11'h7D5: dout  = 8'b11001111; // 2005 : 207 - 0xcf
      11'h7D6: dout  = 8'b00000001; // 2006 :   1 - 0x1
      11'h7D7: dout  = 8'b00001001; // 2007 :   9 - 0x9
      11'h7D8: dout  = 8'b00010111; // 2008 :  23 - 0x17 -- Background 0xfb
      11'h7D9: dout  = 8'b00001101; // 2009 :  13 - 0xd
      11'h7DA: dout  = 8'b00011000; // 2010 :  24 - 0x18
      11'h7DB: dout  = 8'b00100010; // 2011 :  34 - 0x22
      11'h7DC: dout  = 8'b01001011; // 2012 :  75 - 0x4b
      11'h7DD: dout  = 8'b00001101; // 2013 :  13 - 0xd
      11'h7DE: dout  = 8'b00000001; // 2014 :   1 - 0x1
      11'h7DF: dout  = 8'b00100100; // 2015 :  36 - 0x24
      11'h7E0: dout  = 8'b00001010; // 2016 :  10 - 0xa -- Background 0xfc
      11'h7E1: dout  = 8'b00010110; // 2017 :  22 - 0x16
      11'h7E2: dout  = 8'b00001110; // 2018 :  14 - 0xe
      11'h7E3: dout  = 8'b00100010; // 2019 :  34 - 0x22
      11'h7E4: dout  = 8'b10001011; // 2020 : 139 - 0x8b
      11'h7E5: dout  = 8'b00001101; // 2021 :  13 - 0xd
      11'h7E6: dout  = 8'b00000010; // 2022 :   2 - 0x2
      11'h7E7: dout  = 8'b00100100; // 2023 :  36 - 0x24
      11'h7E8: dout  = 8'b00001010; // 2024 :  10 - 0xa -- Background 0xfd
      11'h7E9: dout  = 8'b00010110; // 2025 :  22 - 0x16
      11'h7EA: dout  = 8'b00001110; // 2026 :  14 - 0xe
      11'h7EB: dout  = 8'b00100010; // 2027 :  34 - 0x22
      11'h7EC: dout  = 8'b11101100; // 2028 : 236 - 0xec
      11'h7ED: dout  = 8'b00000100; // 2029 :   4 - 0x4
      11'h7EE: dout  = 8'b00011101; // 2030 :  29 - 0x1d
      11'h7EF: dout  = 8'b00011000; // 2031 :  24 - 0x18
      11'h7F0: dout  = 8'b01010110; // 2032 :  86 - 0x56 -- Background 0xfe
      11'h7F1: dout  = 8'b01010101; // 2033 :  85 - 0x55
      11'h7F2: dout  = 8'b00100011; // 2034 :  35 - 0x23
      11'h7F3: dout  = 8'b11100010; // 2035 : 226 - 0xe2
      11'h7F4: dout  = 8'b00000100; // 2036 :   4 - 0x4
      11'h7F5: dout  = 8'b10011001; // 2037 : 153 - 0x99
      11'h7F6: dout  = 8'b10101010; // 2038 : 170 - 0xaa
      11'h7F7: dout  = 8'b10101010; // 2039 : 170 - 0xaa
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Background 0xff
      11'h7F9: dout  = 8'b11111111; // 2041 : 255 - 0xff
      11'h7FA: dout  = 8'b11111111; // 2042 : 255 - 0xff
      11'h7FB: dout  = 8'b11111111; // 2043 : 255 - 0xff
      11'h7FC: dout  = 8'b11111111; // 2044 : 255 - 0xff
      11'h7FD: dout  = 8'b11111111; // 2045 : 255 - 0xff
      11'h7FE: dout  = 8'b11111111; // 2046 : 255 - 0xff
      11'h7FF: dout  = 8'b11111111; // 2047 : 255 - 0xff
    endcase
  end

endmodule
