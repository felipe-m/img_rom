//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_DONKEYKONG_color0
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      12'h2: dout <= 8'b00000111; //    2 :   7 - 0x7
      12'h3: dout <= 8'b00000111; //    3 :   7 - 0x7
      12'h4: dout <= 8'b00001001; //    4 :   9 - 0x9
      12'h5: dout <= 8'b00001001; //    5 :   9 - 0x9
      12'h6: dout <= 8'b00011100; //    6 :  28 - 0x1c
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00001111; //    8 :  15 - 0xf -- Sprite 0x1
      12'h9: dout <= 8'b00001111; //    9 :  15 - 0xf
      12'hA: dout <= 8'b00001111; //   10 :  15 - 0xf
      12'hB: dout <= 8'b11111111; //   11 : 255 - 0xff
      12'hC: dout <= 8'b11111111; //   12 : 255 - 0xff
      12'hD: dout <= 8'b11111100; //   13 : 252 - 0xfc
      12'hE: dout <= 8'b10000001; //   14 : 129 - 0x81
      12'hF: dout <= 8'b00000001; //   15 :   1 - 0x1
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      12'h11: dout <= 8'b11000000; //   17 : 192 - 0xc0
      12'h12: dout <= 8'b11111000; //   18 : 248 - 0xf8
      12'h13: dout <= 8'b10000000; //   19 : 128 - 0x80
      12'h14: dout <= 8'b00100000; //   20 :  32 - 0x20
      12'h15: dout <= 8'b10010000; //   21 : 144 - 0x90
      12'h16: dout <= 8'b00111100; //   22 :  60 - 0x3c
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b11000000; //   24 : 192 - 0xc0 -- Sprite 0x3
      12'h19: dout <= 8'b11000000; //   25 : 192 - 0xc0
      12'h1A: dout <= 8'b11000000; //   26 : 192 - 0xc0
      12'h1B: dout <= 8'b11110000; //   27 : 240 - 0xf0
      12'h1C: dout <= 8'b11110000; //   28 : 240 - 0xf0
      12'h1D: dout <= 8'b11100000; //   29 : 224 - 0xe0
      12'h1E: dout <= 8'b11000000; //   30 : 192 - 0xc0
      12'h1F: dout <= 8'b11100000; //   31 : 224 - 0xe0
      12'h20: dout <= 8'b00000111; //   32 :   7 - 0x7 -- Sprite 0x4
      12'h21: dout <= 8'b00001111; //   33 :  15 - 0xf
      12'h22: dout <= 8'b00001111; //   34 :  15 - 0xf
      12'h23: dout <= 8'b00010010; //   35 :  18 - 0x12
      12'h24: dout <= 8'b00010011; //   36 :  19 - 0x13
      12'h25: dout <= 8'b00111000; //   37 :  56 - 0x38
      12'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout <= 8'b00001111; //   39 :  15 - 0xf
      12'h28: dout <= 8'b00011111; //   40 :  31 - 0x1f -- Sprite 0x5
      12'h29: dout <= 8'b00011111; //   41 :  31 - 0x1f
      12'h2A: dout <= 8'b00011111; //   42 :  31 - 0x1f
      12'h2B: dout <= 8'b00011000; //   43 :  24 - 0x18
      12'h2C: dout <= 8'b00011001; //   44 :  25 - 0x19
      12'h2D: dout <= 8'b00011110; //   45 :  30 - 0x1e
      12'h2E: dout <= 8'b00011100; //   46 :  28 - 0x1c
      12'h2F: dout <= 8'b00011110; //   47 :  30 - 0x1e
      12'h30: dout <= 8'b10000000; //   48 : 128 - 0x80 -- Sprite 0x6
      12'h31: dout <= 8'b11110000; //   49 : 240 - 0xf0
      12'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout <= 8'b01000000; //   51 :  64 - 0x40
      12'h34: dout <= 8'b00100000; //   52 :  32 - 0x20
      12'h35: dout <= 8'b01111000; //   53 : 120 - 0x78
      12'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      12'h37: dout <= 8'b11000000; //   55 : 192 - 0xc0
      12'h38: dout <= 8'b11100000; //   56 : 224 - 0xe0 -- Sprite 0x7
      12'h39: dout <= 8'b01100000; //   57 :  96 - 0x60
      12'h3A: dout <= 8'b11110000; //   58 : 240 - 0xf0
      12'h3B: dout <= 8'b11110000; //   59 : 240 - 0xf0
      12'h3C: dout <= 8'b11110000; //   60 : 240 - 0xf0
      12'h3D: dout <= 8'b11100000; //   61 : 224 - 0xe0
      12'h3E: dout <= 8'b11100000; //   62 : 224 - 0xe0
      12'h3F: dout <= 8'b11110000; //   63 : 240 - 0xf0
      12'h40: dout <= 8'b00000111; //   64 :   7 - 0x7 -- Sprite 0x8
      12'h41: dout <= 8'b00001111; //   65 :  15 - 0xf
      12'h42: dout <= 8'b00001111; //   66 :  15 - 0xf
      12'h43: dout <= 8'b00010010; //   67 :  18 - 0x12
      12'h44: dout <= 8'b00010011; //   68 :  19 - 0x13
      12'h45: dout <= 8'b00111000; //   69 :  56 - 0x38
      12'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout <= 8'b00111111; //   71 :  63 - 0x3f
      12'h48: dout <= 8'b00111111; //   72 :  63 - 0x3f -- Sprite 0x9
      12'h49: dout <= 8'b00001110; //   73 :  14 - 0xe
      12'h4A: dout <= 8'b00001111; //   74 :  15 - 0xf
      12'h4B: dout <= 8'b00011111; //   75 :  31 - 0x1f
      12'h4C: dout <= 8'b00111111; //   76 :  63 - 0x3f
      12'h4D: dout <= 8'b01111100; //   77 : 124 - 0x7c
      12'h4E: dout <= 8'b01110000; //   78 : 112 - 0x70
      12'h4F: dout <= 8'b00111000; //   79 :  56 - 0x38
      12'h50: dout <= 8'b10000000; //   80 : 128 - 0x80 -- Sprite 0xa
      12'h51: dout <= 8'b11110000; //   81 : 240 - 0xf0
      12'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      12'h53: dout <= 8'b01000000; //   83 :  64 - 0x40
      12'h54: dout <= 8'b00100000; //   84 :  32 - 0x20
      12'h55: dout <= 8'b01111000; //   85 : 120 - 0x78
      12'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout <= 8'b11000000; //   87 : 192 - 0xc0
      12'h58: dout <= 8'b11110000; //   88 : 240 - 0xf0 -- Sprite 0xb
      12'h59: dout <= 8'b11111000; //   89 : 248 - 0xf8
      12'h5A: dout <= 8'b11100100; //   90 : 228 - 0xe4
      12'h5B: dout <= 8'b11111100; //   91 : 252 - 0xfc
      12'h5C: dout <= 8'b11111100; //   92 : 252 - 0xfc
      12'h5D: dout <= 8'b01111100; //   93 : 124 - 0x7c
      12'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      12'h61: dout <= 8'b00000010; //   97 :   2 - 0x2
      12'h62: dout <= 8'b00000110; //   98 :   6 - 0x6
      12'h63: dout <= 8'b00000111; //   99 :   7 - 0x7
      12'h64: dout <= 8'b00001001; //  100 :   9 - 0x9
      12'h65: dout <= 8'b00001001; //  101 :   9 - 0x9
      12'h66: dout <= 8'b00011101; //  102 :  29 - 0x1d
      12'h67: dout <= 8'b00000011; //  103 :   3 - 0x3
      12'h68: dout <= 8'b00001111; //  104 :  15 - 0xf -- Sprite 0xd
      12'h69: dout <= 8'b00001111; //  105 :  15 - 0xf
      12'h6A: dout <= 8'b00001111; //  106 :  15 - 0xf
      12'h6B: dout <= 8'b11111111; //  107 : 255 - 0xff
      12'h6C: dout <= 8'b11111111; //  108 : 255 - 0xff
      12'h6D: dout <= 8'b11111100; //  109 : 252 - 0xfc
      12'h6E: dout <= 8'b10000001; //  110 : 129 - 0x81
      12'h6F: dout <= 8'b00000001; //  111 :   1 - 0x1
      12'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      12'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      12'h72: dout <= 8'b00111000; //  114 :  56 - 0x38
      12'h73: dout <= 8'b11000000; //  115 : 192 - 0xc0
      12'h74: dout <= 8'b11100000; //  116 : 224 - 0xe0
      12'h75: dout <= 8'b11010000; //  117 : 208 - 0xd0
      12'h76: dout <= 8'b11111100; //  118 : 252 - 0xfc
      12'h77: dout <= 8'b11000000; //  119 : 192 - 0xc0
      12'h78: dout <= 8'b11100000; //  120 : 224 - 0xe0 -- Sprite 0xf
      12'h79: dout <= 8'b11100000; //  121 : 224 - 0xe0
      12'h7A: dout <= 8'b10110000; //  122 : 176 - 0xb0
      12'h7B: dout <= 8'b11110000; //  123 : 240 - 0xf0
      12'h7C: dout <= 8'b11110000; //  124 : 240 - 0xf0
      12'h7D: dout <= 8'b11100000; //  125 : 224 - 0xe0
      12'h7E: dout <= 8'b11000000; //  126 : 192 - 0xc0
      12'h7F: dout <= 8'b11100000; //  127 : 224 - 0xe0
      12'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout <= 8'b00000011; //  129 :   3 - 0x3
      12'h82: dout <= 8'b00000111; //  130 :   7 - 0x7
      12'h83: dout <= 8'b00000111; //  131 :   7 - 0x7
      12'h84: dout <= 8'b00001001; //  132 :   9 - 0x9
      12'h85: dout <= 8'b00001001; //  133 :   9 - 0x9
      12'h86: dout <= 8'b00011100; //  134 :  28 - 0x1c
      12'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout <= 8'b00001111; //  136 :  15 - 0xf -- Sprite 0x11
      12'h89: dout <= 8'b00001111; //  137 :  15 - 0xf
      12'h8A: dout <= 8'b00001111; //  138 :  15 - 0xf
      12'h8B: dout <= 8'b11111111; //  139 : 255 - 0xff
      12'h8C: dout <= 8'b11111111; //  140 : 255 - 0xff
      12'h8D: dout <= 8'b11111100; //  141 : 252 - 0xfc
      12'h8E: dout <= 8'b10000001; //  142 : 129 - 0x81
      12'h8F: dout <= 8'b00000001; //  143 :   1 - 0x1
      12'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      12'h91: dout <= 8'b11000000; //  145 : 192 - 0xc0
      12'h92: dout <= 8'b11111000; //  146 : 248 - 0xf8
      12'h93: dout <= 8'b10000000; //  147 : 128 - 0x80
      12'h94: dout <= 8'b00100000; //  148 :  32 - 0x20
      12'h95: dout <= 8'b10010000; //  149 : 144 - 0x90
      12'h96: dout <= 8'b00111100; //  150 :  60 - 0x3c
      12'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout <= 8'b11100000; //  152 : 224 - 0xe0 -- Sprite 0x13
      12'h99: dout <= 8'b11110000; //  153 : 240 - 0xf0
      12'h9A: dout <= 8'b11110000; //  154 : 240 - 0xf0
      12'h9B: dout <= 8'b11110000; //  155 : 240 - 0xf0
      12'h9C: dout <= 8'b11110000; //  156 : 240 - 0xf0
      12'h9D: dout <= 8'b11100000; //  157 : 224 - 0xe0
      12'h9E: dout <= 8'b11000000; //  158 : 192 - 0xc0
      12'h9F: dout <= 8'b11100000; //  159 : 224 - 0xe0
      12'hA0: dout <= 8'b00000100; //  160 :   4 - 0x4 -- Sprite 0x14
      12'hA1: dout <= 8'b00001100; //  161 :  12 - 0xc
      12'hA2: dout <= 8'b00001100; //  162 :  12 - 0xc
      12'hA3: dout <= 8'b00010011; //  163 :  19 - 0x13
      12'hA4: dout <= 8'b00010011; //  164 :  19 - 0x13
      12'hA5: dout <= 8'b00111011; //  165 :  59 - 0x3b
      12'hA6: dout <= 8'b00000111; //  166 :   7 - 0x7
      12'hA7: dout <= 8'b00001111; //  167 :  15 - 0xf
      12'hA8: dout <= 8'b00001111; //  168 :  15 - 0xf -- Sprite 0x15
      12'hA9: dout <= 8'b00001111; //  169 :  15 - 0xf
      12'hAA: dout <= 8'b00001111; //  170 :  15 - 0xf
      12'hAB: dout <= 8'b00011111; //  171 :  31 - 0x1f
      12'hAC: dout <= 8'b00011111; //  172 :  31 - 0x1f
      12'hAD: dout <= 8'b00011110; //  173 :  30 - 0x1e
      12'hAE: dout <= 8'b00011100; //  174 :  28 - 0x1c
      12'hAF: dout <= 8'b00011110; //  175 :  30 - 0x1e
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      12'hB1: dout <= 8'b01110000; //  177 : 112 - 0x70
      12'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      12'hB3: dout <= 8'b11000000; //  179 : 192 - 0xc0
      12'hB4: dout <= 8'b10100000; //  180 : 160 - 0xa0
      12'hB5: dout <= 8'b11111000; //  181 : 248 - 0xf8
      12'hB6: dout <= 8'b10000000; //  182 : 128 - 0x80
      12'hB7: dout <= 8'b11000000; //  183 : 192 - 0xc0
      12'hB8: dout <= 8'b11100000; //  184 : 224 - 0xe0 -- Sprite 0x17
      12'hB9: dout <= 8'b01100000; //  185 :  96 - 0x60
      12'hBA: dout <= 8'b11110000; //  186 : 240 - 0xf0
      12'hBB: dout <= 8'b11110000; //  187 : 240 - 0xf0
      12'hBC: dout <= 8'b11110000; //  188 : 240 - 0xf0
      12'hBD: dout <= 8'b11100000; //  189 : 224 - 0xe0
      12'hBE: dout <= 8'b11100000; //  190 : 224 - 0xe0
      12'hBF: dout <= 8'b11110000; //  191 : 240 - 0xf0
      12'hC0: dout <= 8'b00000111; //  192 :   7 - 0x7 -- Sprite 0x18
      12'hC1: dout <= 8'b00001111; //  193 :  15 - 0xf
      12'hC2: dout <= 8'b00001111; //  194 :  15 - 0xf
      12'hC3: dout <= 8'b00010010; //  195 :  18 - 0x12
      12'hC4: dout <= 8'b00010011; //  196 :  19 - 0x13
      12'hC5: dout <= 8'b00111000; //  197 :  56 - 0x38
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00001111; //  199 :  15 - 0xf
      12'hC8: dout <= 8'b00011111; //  200 :  31 - 0x1f -- Sprite 0x19
      12'hC9: dout <= 8'b00011111; //  201 :  31 - 0x1f
      12'hCA: dout <= 8'b00011111; //  202 :  31 - 0x1f
      12'hCB: dout <= 8'b00011111; //  203 :  31 - 0x1f
      12'hCC: dout <= 8'b00011111; //  204 :  31 - 0x1f
      12'hCD: dout <= 8'b00011110; //  205 :  30 - 0x1e
      12'hCE: dout <= 8'b00011100; //  206 :  28 - 0x1c
      12'hCF: dout <= 8'b00011110; //  207 :  30 - 0x1e
      12'hD0: dout <= 8'b10000000; //  208 : 128 - 0x80 -- Sprite 0x1a
      12'hD1: dout <= 8'b11110000; //  209 : 240 - 0xf0
      12'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      12'hD3: dout <= 8'b01000000; //  211 :  64 - 0x40
      12'hD4: dout <= 8'b00100000; //  212 :  32 - 0x20
      12'hD5: dout <= 8'b01111000; //  213 : 120 - 0x78
      12'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout <= 8'b11000000; //  215 : 192 - 0xc0
      12'hD8: dout <= 8'b11111000; //  216 : 248 - 0xf8 -- Sprite 0x1b
      12'hD9: dout <= 8'b11111000; //  217 : 248 - 0xf8
      12'hDA: dout <= 8'b11110000; //  218 : 240 - 0xf0
      12'hDB: dout <= 8'b11110000; //  219 : 240 - 0xf0
      12'hDC: dout <= 8'b11110000; //  220 : 240 - 0xf0
      12'hDD: dout <= 8'b11100000; //  221 : 224 - 0xe0
      12'hDE: dout <= 8'b11100000; //  222 : 224 - 0xe0
      12'hDF: dout <= 8'b11110000; //  223 : 240 - 0xf0
      12'hE0: dout <= 8'b00000100; //  224 :   4 - 0x4 -- Sprite 0x1c
      12'hE1: dout <= 8'b00001100; //  225 :  12 - 0xc
      12'hE2: dout <= 8'b00001100; //  226 :  12 - 0xc
      12'hE3: dout <= 8'b00010011; //  227 :  19 - 0x13
      12'hE4: dout <= 8'b00010011; //  228 :  19 - 0x13
      12'hE5: dout <= 8'b00111111; //  229 :  63 - 0x3f
      12'hE6: dout <= 8'b00000111; //  230 :   7 - 0x7
      12'hE7: dout <= 8'b00001111; //  231 :  15 - 0xf
      12'hE8: dout <= 8'b00001111; //  232 :  15 - 0xf -- Sprite 0x1d
      12'hE9: dout <= 8'b00001111; //  233 :  15 - 0xf
      12'hEA: dout <= 8'b00001111; //  234 :  15 - 0xf
      12'hEB: dout <= 8'b00011111; //  235 :  31 - 0x1f
      12'hEC: dout <= 8'b00111111; //  236 :  63 - 0x3f
      12'hED: dout <= 8'b01111100; //  237 : 124 - 0x7c
      12'hEE: dout <= 8'b01110000; //  238 : 112 - 0x70
      12'hEF: dout <= 8'b00111000; //  239 :  56 - 0x38
      12'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x1e
      12'hF1: dout <= 8'b01110000; //  241 : 112 - 0x70
      12'hF2: dout <= 8'b00000000; //  242 :   0 - 0x0
      12'hF3: dout <= 8'b11000000; //  243 : 192 - 0xc0
      12'hF4: dout <= 8'b10100000; //  244 : 160 - 0xa0
      12'hF5: dout <= 8'b11111000; //  245 : 248 - 0xf8
      12'hF6: dout <= 8'b10000000; //  246 : 128 - 0x80
      12'hF7: dout <= 8'b11000000; //  247 : 192 - 0xc0
      12'hF8: dout <= 8'b11000000; //  248 : 192 - 0xc0 -- Sprite 0x1f
      12'hF9: dout <= 8'b01100000; //  249 :  96 - 0x60
      12'hFA: dout <= 8'b11100100; //  250 : 228 - 0xe4
      12'hFB: dout <= 8'b11111100; //  251 : 252 - 0xfc
      12'hFC: dout <= 8'b11111100; //  252 : 252 - 0xfc
      12'hFD: dout <= 8'b01111100; //  253 : 124 - 0x7c
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x20
      12'h101: dout <= 8'b00001111; //  257 :  15 - 0xf
      12'h102: dout <= 8'b00001111; //  258 :  15 - 0xf
      12'h103: dout <= 8'b00010010; //  259 :  18 - 0x12
      12'h104: dout <= 8'b00010011; //  260 :  19 - 0x13
      12'h105: dout <= 8'b00111000; //  261 :  56 - 0x38
      12'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout <= 8'b00000111; //  263 :   7 - 0x7
      12'h108: dout <= 8'b00001111; //  264 :  15 - 0xf -- Sprite 0x21
      12'h109: dout <= 8'b00001111; //  265 :  15 - 0xf
      12'h10A: dout <= 8'b00001111; //  266 :  15 - 0xf
      12'h10B: dout <= 8'b00011111; //  267 :  31 - 0x1f
      12'h10C: dout <= 8'b00111111; //  268 :  63 - 0x3f
      12'h10D: dout <= 8'b01111100; //  269 : 124 - 0x7c
      12'h10E: dout <= 8'b01110000; //  270 : 112 - 0x70
      12'h10F: dout <= 8'b00111000; //  271 :  56 - 0x38
      12'h110: dout <= 8'b10000000; //  272 : 128 - 0x80 -- Sprite 0x22
      12'h111: dout <= 8'b11110000; //  273 : 240 - 0xf0
      12'h112: dout <= 8'b00000000; //  274 :   0 - 0x0
      12'h113: dout <= 8'b01000000; //  275 :  64 - 0x40
      12'h114: dout <= 8'b00100000; //  276 :  32 - 0x20
      12'h115: dout <= 8'b01111000; //  277 : 120 - 0x78
      12'h116: dout <= 8'b00000000; //  278 :   0 - 0x0
      12'h117: dout <= 8'b11000000; //  279 : 192 - 0xc0
      12'h118: dout <= 8'b11111000; //  280 : 248 - 0xf8 -- Sprite 0x23
      12'h119: dout <= 8'b11111000; //  281 : 248 - 0xf8
      12'h11A: dout <= 8'b11100000; //  282 : 224 - 0xe0
      12'h11B: dout <= 8'b11111100; //  283 : 252 - 0xfc
      12'h11C: dout <= 8'b11111100; //  284 : 252 - 0xfc
      12'h11D: dout <= 8'b01111100; //  285 : 124 - 0x7c
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      12'h121: dout <= 8'b00000111; //  289 :   7 - 0x7
      12'h122: dout <= 8'b00000111; //  290 :   7 - 0x7
      12'h123: dout <= 8'b00001111; //  291 :  15 - 0xf
      12'h124: dout <= 8'b00001111; //  292 :  15 - 0xf
      12'h125: dout <= 8'b00111000; //  293 :  56 - 0x38
      12'h126: dout <= 8'b01111111; //  294 : 127 - 0x7f
      12'h127: dout <= 8'b01111111; //  295 : 127 - 0x7f
      12'h128: dout <= 8'b00011111; //  296 :  31 - 0x1f -- Sprite 0x25
      12'h129: dout <= 8'b00011111; //  297 :  31 - 0x1f
      12'h12A: dout <= 8'b00011111; //  298 :  31 - 0x1f
      12'h12B: dout <= 8'b00011111; //  299 :  31 - 0x1f
      12'h12C: dout <= 8'b00001111; //  300 :  15 - 0xf
      12'h12D: dout <= 8'b00001111; //  301 :  15 - 0xf
      12'h12E: dout <= 8'b00001111; //  302 :  15 - 0xf
      12'h12F: dout <= 8'b00000111; //  303 :   7 - 0x7
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout <= 8'b11100000; //  305 : 224 - 0xe0
      12'h132: dout <= 8'b11111000; //  306 : 248 - 0xf8
      12'h133: dout <= 8'b11111100; //  307 : 252 - 0xfc
      12'h134: dout <= 8'b11111100; //  308 : 252 - 0xfc
      12'h135: dout <= 8'b00011100; //  309 :  28 - 0x1c
      12'h136: dout <= 8'b11111000; //  310 : 248 - 0xf8
      12'h137: dout <= 8'b11111000; //  311 : 248 - 0xf8
      12'h138: dout <= 8'b11111000; //  312 : 248 - 0xf8 -- Sprite 0x27
      12'h139: dout <= 8'b11111100; //  313 : 252 - 0xfc
      12'h13A: dout <= 8'b11111100; //  314 : 252 - 0xfc
      12'h13B: dout <= 8'b11111000; //  315 : 248 - 0xf8
      12'h13C: dout <= 8'b01111000; //  316 : 120 - 0x78
      12'h13D: dout <= 8'b10000000; //  317 : 128 - 0x80
      12'h13E: dout <= 8'b11000000; //  318 : 192 - 0xc0
      12'h13F: dout <= 8'b11000000; //  319 : 192 - 0xc0
      12'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout <= 8'b00000011; //  321 :   3 - 0x3
      12'h142: dout <= 8'b00000111; //  322 :   7 - 0x7
      12'h143: dout <= 8'b00000111; //  323 :   7 - 0x7
      12'h144: dout <= 8'b00001001; //  324 :   9 - 0x9
      12'h145: dout <= 8'b00001001; //  325 :   9 - 0x9
      12'h146: dout <= 8'b00011100; //  326 :  28 - 0x1c
      12'h147: dout <= 8'b00000000; //  327 :   0 - 0x0
      12'h148: dout <= 8'b00011111; //  328 :  31 - 0x1f -- Sprite 0x29
      12'h149: dout <= 8'b00001111; //  329 :  15 - 0xf
      12'h14A: dout <= 8'b00000111; //  330 :   7 - 0x7
      12'h14B: dout <= 8'b00110111; //  331 :  55 - 0x37
      12'h14C: dout <= 8'b01111111; //  332 : 127 - 0x7f
      12'h14D: dout <= 8'b11011111; //  333 : 223 - 0xdf
      12'h14E: dout <= 8'b00001111; //  334 :  15 - 0xf
      12'h14F: dout <= 8'b00000110; //  335 :   6 - 0x6
      12'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x2a
      12'h151: dout <= 8'b11000000; //  337 : 192 - 0xc0
      12'h152: dout <= 8'b11111000; //  338 : 248 - 0xf8
      12'h153: dout <= 8'b10000000; //  339 : 128 - 0x80
      12'h154: dout <= 8'b00100000; //  340 :  32 - 0x20
      12'h155: dout <= 8'b10010000; //  341 : 144 - 0x90
      12'h156: dout <= 8'b00111100; //  342 :  60 - 0x3c
      12'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout <= 8'b11100100; //  344 : 228 - 0xe4 -- Sprite 0x2b
      12'h159: dout <= 8'b11111110; //  345 : 254 - 0xfe
      12'h15A: dout <= 8'b01110000; //  346 : 112 - 0x70
      12'h15B: dout <= 8'b11110001; //  347 : 241 - 0xf1
      12'h15C: dout <= 8'b11111111; //  348 : 255 - 0xff
      12'h15D: dout <= 8'b11111111; //  349 : 255 - 0xff
      12'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00000111; //  352 :   7 - 0x7 -- Sprite 0x2c
      12'h161: dout <= 8'b00001111; //  353 :  15 - 0xf
      12'h162: dout <= 8'b00001111; //  354 :  15 - 0xf
      12'h163: dout <= 8'b00010010; //  355 :  18 - 0x12
      12'h164: dout <= 8'b00010011; //  356 :  19 - 0x13
      12'h165: dout <= 8'b00111000; //  357 :  56 - 0x38
      12'h166: dout <= 8'b01110000; //  358 : 112 - 0x70
      12'h167: dout <= 8'b11111111; //  359 : 255 - 0xff
      12'h168: dout <= 8'b11011111; //  360 : 223 - 0xdf -- Sprite 0x2d
      12'h169: dout <= 8'b00011110; //  361 :  30 - 0x1e
      12'h16A: dout <= 8'b00011111; //  362 :  31 - 0x1f
      12'h16B: dout <= 8'b00011111; //  363 :  31 - 0x1f
      12'h16C: dout <= 8'b00011111; //  364 :  31 - 0x1f
      12'h16D: dout <= 8'b00001111; //  365 :  15 - 0xf
      12'h16E: dout <= 8'b00000111; //  366 :   7 - 0x7
      12'h16F: dout <= 8'b00000001; //  367 :   1 - 0x1
      12'h170: dout <= 8'b10000000; //  368 : 128 - 0x80 -- Sprite 0x2e
      12'h171: dout <= 8'b11110000; //  369 : 240 - 0xf0
      12'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout <= 8'b01000000; //  371 :  64 - 0x40
      12'h174: dout <= 8'b00100000; //  372 :  32 - 0x20
      12'h175: dout <= 8'b01111000; //  373 : 120 - 0x78
      12'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout <= 8'b11111100; //  375 : 252 - 0xfc
      12'h178: dout <= 8'b11110000; //  376 : 240 - 0xf0 -- Sprite 0x2f
      12'h179: dout <= 8'b11100000; //  377 : 224 - 0xe0
      12'h17A: dout <= 8'b11100000; //  378 : 224 - 0xe0
      12'h17B: dout <= 8'b11110000; //  379 : 240 - 0xf0
      12'h17C: dout <= 8'b11111010; //  380 : 250 - 0xfa
      12'h17D: dout <= 8'b11111110; //  381 : 254 - 0xfe
      12'h17E: dout <= 8'b11111100; //  382 : 252 - 0xfc
      12'h17F: dout <= 8'b11011000; //  383 : 216 - 0xd8
      12'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x30
      12'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      12'h182: dout <= 8'b00000111; //  386 :   7 - 0x7
      12'h183: dout <= 8'b00001000; //  387 :   8 - 0x8
      12'h184: dout <= 8'b00010000; //  388 :  16 - 0x10
      12'h185: dout <= 8'b00100000; //  389 :  32 - 0x20
      12'h186: dout <= 8'b01000000; //  390 :  64 - 0x40
      12'h187: dout <= 8'b01000000; //  391 :  64 - 0x40
      12'h188: dout <= 8'b01000000; //  392 :  64 - 0x40 -- Sprite 0x31
      12'h189: dout <= 8'b01000000; //  393 :  64 - 0x40
      12'h18A: dout <= 8'b00100000; //  394 :  32 - 0x20
      12'h18B: dout <= 8'b00010000; //  395 :  16 - 0x10
      12'h18C: dout <= 8'b00001000; //  396 :   8 - 0x8
      12'h18D: dout <= 8'b00000111; //  397 :   7 - 0x7
      12'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      12'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      12'h192: dout <= 8'b11100000; //  402 : 224 - 0xe0
      12'h193: dout <= 8'b00010000; //  403 :  16 - 0x10
      12'h194: dout <= 8'b00001000; //  404 :   8 - 0x8
      12'h195: dout <= 8'b00000100; //  405 :   4 - 0x4
      12'h196: dout <= 8'b00000010; //  406 :   2 - 0x2
      12'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      12'h198: dout <= 8'b00000010; //  408 :   2 - 0x2 -- Sprite 0x33
      12'h199: dout <= 8'b00000010; //  409 :   2 - 0x2
      12'h19A: dout <= 8'b00000100; //  410 :   4 - 0x4
      12'h19B: dout <= 8'b00001000; //  411 :   8 - 0x8
      12'h19C: dout <= 8'b00010000; //  412 :  16 - 0x10
      12'h19D: dout <= 8'b11100000; //  413 : 224 - 0xe0
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      12'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      12'h1A2: dout <= 8'b00000000; //  418 :   0 - 0x0
      12'h1A3: dout <= 8'b00000000; //  419 :   0 - 0x0
      12'h1A4: dout <= 8'b00000011; //  420 :   3 - 0x3
      12'h1A5: dout <= 8'b00000100; //  421 :   4 - 0x4
      12'h1A6: dout <= 8'b00001000; //  422 :   8 - 0x8
      12'h1A7: dout <= 8'b00010000; //  423 :  16 - 0x10
      12'h1A8: dout <= 8'b00010000; //  424 :  16 - 0x10 -- Sprite 0x35
      12'h1A9: dout <= 8'b00001000; //  425 :   8 - 0x8
      12'h1AA: dout <= 8'b00000100; //  426 :   4 - 0x4
      12'h1AB: dout <= 8'b00000011; //  427 :   3 - 0x3
      12'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      12'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      12'h1B3: dout <= 8'b00000000; //  435 :   0 - 0x0
      12'h1B4: dout <= 8'b11000000; //  436 : 192 - 0xc0
      12'h1B5: dout <= 8'b00100000; //  437 :  32 - 0x20
      12'h1B6: dout <= 8'b00010000; //  438 :  16 - 0x10
      12'h1B7: dout <= 8'b00001000; //  439 :   8 - 0x8
      12'h1B8: dout <= 8'b00001000; //  440 :   8 - 0x8 -- Sprite 0x37
      12'h1B9: dout <= 8'b00010000; //  441 :  16 - 0x10
      12'h1BA: dout <= 8'b00100000; //  442 :  32 - 0x20
      12'h1BB: dout <= 8'b11000000; //  443 : 192 - 0xc0
      12'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      12'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout <= 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout <= 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout <= 8'b00000000; //  452 :   0 - 0x0
      12'h1C5: dout <= 8'b00000000; //  453 :   0 - 0x0
      12'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      12'h1C7: dout <= 8'b00000001; //  455 :   1 - 0x1
      12'h1C8: dout <= 8'b00000010; //  456 :   2 - 0x2 -- Sprite 0x39
      12'h1C9: dout <= 8'b00000001; //  457 :   1 - 0x1
      12'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout <= 8'b00000000; //  467 :   0 - 0x0
      12'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      12'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      12'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b10000000; //  472 : 128 - 0x80 -- Sprite 0x3b
      12'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout <= 8'b00000001; //  483 :   1 - 0x1
      12'h1E4: dout <= 8'b00100001; //  484 :  33 - 0x21
      12'h1E5: dout <= 8'b00010000; //  485 :  16 - 0x10
      12'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b01100000; //  488 :  96 - 0x60 -- Sprite 0x3d
      12'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout <= 8'b00010000; //  491 :  16 - 0x10
      12'h1EC: dout <= 8'b00100001; //  492 :  33 - 0x21
      12'h1ED: dout <= 8'b00000001; //  493 :   1 - 0x1
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      12'h1F3: dout <= 8'b00000000; //  499 :   0 - 0x0
      12'h1F4: dout <= 8'b00001000; //  500 :   8 - 0x8
      12'h1F5: dout <= 8'b00010000; //  501 :  16 - 0x10
      12'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b00001100; //  504 :  12 - 0xc -- Sprite 0x3f
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout <= 8'b00010000; //  507 :  16 - 0x10
      12'h1FC: dout <= 8'b00001000; //  508 :   8 - 0x8
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000100; //  512 :   4 - 0x4 -- Sprite 0x40
      12'h201: dout <= 8'b00000010; //  513 :   2 - 0x2
      12'h202: dout <= 8'b00000001; //  514 :   1 - 0x1
      12'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      12'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000001; //  526 :   1 - 0x1
      12'h20F: dout <= 8'b00000011; //  527 :   3 - 0x3
      12'h210: dout <= 8'b00000111; //  528 :   7 - 0x7 -- Sprite 0x42
      12'h211: dout <= 8'b00000111; //  529 :   7 - 0x7
      12'h212: dout <= 8'b00000111; //  530 :   7 - 0x7
      12'h213: dout <= 8'b00000011; //  531 :   3 - 0x3
      12'h214: dout <= 8'b00000001; //  532 :   1 - 0x1
      12'h215: dout <= 8'b00000000; //  533 :   0 - 0x0
      12'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      12'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      12'h221: dout <= 8'b01000010; //  545 :  66 - 0x42
      12'h222: dout <= 8'b00111001; //  546 :  57 - 0x39
      12'h223: dout <= 8'b11111111; //  547 : 255 - 0xff
      12'h224: dout <= 8'b11111111; //  548 : 255 - 0xff
      12'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      12'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      12'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      12'h228: dout <= 8'b01111111; //  552 : 127 - 0x7f -- Sprite 0x45
      12'h229: dout <= 8'b00111111; //  553 :  63 - 0x3f
      12'h22A: dout <= 8'b00011111; //  554 :  31 - 0x1f
      12'h22B: dout <= 8'b00001111; //  555 :  15 - 0xf
      12'h22C: dout <= 8'b00011111; //  556 :  31 - 0x1f
      12'h22D: dout <= 8'b11111111; //  557 : 255 - 0xff
      12'h22E: dout <= 8'b11111111; //  558 : 255 - 0xff
      12'h22F: dout <= 8'b11111111; //  559 : 255 - 0xff
      12'h230: dout <= 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x46
      12'h231: dout <= 8'b11110111; //  561 : 247 - 0xf7
      12'h232: dout <= 8'b11101111; //  562 : 239 - 0xef
      12'h233: dout <= 8'b11111111; //  563 : 255 - 0xff
      12'h234: dout <= 8'b11111111; //  564 : 255 - 0xff
      12'h235: dout <= 8'b11111110; //  565 : 254 - 0xfe
      12'h236: dout <= 8'b01111110; //  566 : 126 - 0x7e
      12'h237: dout <= 8'b00111110; //  567 :  62 - 0x3e
      12'h238: dout <= 8'b00000111; //  568 :   7 - 0x7 -- Sprite 0x47
      12'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      12'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout <= 8'b11000000; //  579 : 192 - 0xc0
      12'h244: dout <= 8'b11100000; //  580 : 224 - 0xe0
      12'h245: dout <= 8'b11110000; //  581 : 240 - 0xf0
      12'h246: dout <= 8'b11011011; //  582 : 219 - 0xdb
      12'h247: dout <= 8'b11110110; //  583 : 246 - 0xf6
      12'h248: dout <= 8'b11001011; //  584 : 203 - 0xcb -- Sprite 0x49
      12'h249: dout <= 8'b11100000; //  585 : 224 - 0xe0
      12'h24A: dout <= 8'b11000100; //  586 : 196 - 0xc4
      12'h24B: dout <= 8'b00000010; //  587 :   2 - 0x2
      12'h24C: dout <= 8'b11010001; //  588 : 209 - 0xd1
      12'h24D: dout <= 8'b11100001; //  589 : 225 - 0xe1
      12'h24E: dout <= 8'b11010001; //  590 : 209 - 0xd1
      12'h24F: dout <= 8'b10000011; //  591 : 131 - 0x83
      12'h250: dout <= 8'b00001111; //  592 :  15 - 0xf -- Sprite 0x4a
      12'h251: dout <= 8'b11111111; //  593 : 255 - 0xff
      12'h252: dout <= 8'b11100000; //  594 : 224 - 0xe0
      12'h253: dout <= 8'b10001111; //  595 : 143 - 0x8f
      12'h254: dout <= 8'b01101110; //  596 : 110 - 0x6e
      12'h255: dout <= 8'b01000100; //  597 :  68 - 0x44
      12'h256: dout <= 8'b11101110; //  598 : 238 - 0xee
      12'h257: dout <= 8'b01100000; //  599 :  96 - 0x60
      12'h258: dout <= 8'b10000011; //  600 : 131 - 0x83 -- Sprite 0x4b
      12'h259: dout <= 8'b11100000; //  601 : 224 - 0xe0
      12'h25A: dout <= 8'b11100100; //  602 : 228 - 0xe4
      12'h25B: dout <= 8'b11000110; //  603 : 198 - 0xc6
      12'h25C: dout <= 8'b01100001; //  604 :  97 - 0x61
      12'h25D: dout <= 8'b00110011; //  605 :  51 - 0x33
      12'h25E: dout <= 8'b00011111; //  606 :  31 - 0x1f
      12'h25F: dout <= 8'b00001111; //  607 :  15 - 0xf
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      12'h261: dout <= 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout <= 8'b00000000; //  610 :   0 - 0x0
      12'h263: dout <= 8'b00000011; //  611 :   3 - 0x3
      12'h264: dout <= 8'b00000111; //  612 :   7 - 0x7
      12'h265: dout <= 8'b00001111; //  613 :  15 - 0xf
      12'h266: dout <= 8'b01011011; //  614 :  91 - 0x5b
      12'h267: dout <= 8'b10100111; //  615 : 167 - 0xa7
      12'h268: dout <= 8'b01110011; //  616 : 115 - 0x73 -- Sprite 0x4d
      12'h269: dout <= 8'b00000111; //  617 :   7 - 0x7
      12'h26A: dout <= 8'b00100111; //  618 :  39 - 0x27
      12'h26B: dout <= 8'b01000000; //  619 :  64 - 0x40
      12'h26C: dout <= 8'b10001011; //  620 : 139 - 0x8b
      12'h26D: dout <= 8'b10000111; //  621 : 135 - 0x87
      12'h26E: dout <= 8'b10001011; //  622 : 139 - 0x8b
      12'h26F: dout <= 8'b11000001; //  623 : 193 - 0xc1
      12'h270: dout <= 8'b11110000; //  624 : 240 - 0xf0 -- Sprite 0x4e
      12'h271: dout <= 8'b11111111; //  625 : 255 - 0xff
      12'h272: dout <= 8'b00001111; //  626 :  15 - 0xf
      12'h273: dout <= 8'b11100001; //  627 : 225 - 0xe1
      12'h274: dout <= 8'b11101100; //  628 : 236 - 0xec
      12'h275: dout <= 8'b01000100; //  629 :  68 - 0x44
      12'h276: dout <= 8'b11101110; //  630 : 238 - 0xee
      12'h277: dout <= 8'b00001100; //  631 :  12 - 0xc
      12'h278: dout <= 8'b10000000; //  632 : 128 - 0x80 -- Sprite 0x4f
      12'h279: dout <= 8'b00001110; //  633 :  14 - 0xe
      12'h27A: dout <= 8'b01001110; //  634 :  78 - 0x4e
      12'h27B: dout <= 8'b11000110; //  635 : 198 - 0xc6
      12'h27C: dout <= 8'b00001100; //  636 :  12 - 0xc
      12'h27D: dout <= 8'b10011000; //  637 : 152 - 0x98
      12'h27E: dout <= 8'b11110000; //  638 : 240 - 0xf0
      12'h27F: dout <= 8'b11100000; //  639 : 224 - 0xe0
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout <= 8'b01000010; //  641 :  66 - 0x42
      12'h282: dout <= 8'b10011100; //  642 : 156 - 0x9c
      12'h283: dout <= 8'b11111111; //  643 : 255 - 0xff
      12'h284: dout <= 8'b11111111; //  644 : 255 - 0xff
      12'h285: dout <= 8'b11111111; //  645 : 255 - 0xff
      12'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      12'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      12'h288: dout <= 8'b11111110; //  648 : 254 - 0xfe -- Sprite 0x51
      12'h289: dout <= 8'b11111100; //  649 : 252 - 0xfc
      12'h28A: dout <= 8'b11111000; //  650 : 248 - 0xf8
      12'h28B: dout <= 8'b11110000; //  651 : 240 - 0xf0
      12'h28C: dout <= 8'b11111000; //  652 : 248 - 0xf8
      12'h28D: dout <= 8'b11111111; //  653 : 255 - 0xff
      12'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      12'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      12'h290: dout <= 8'b00011111; //  656 :  31 - 0x1f -- Sprite 0x52
      12'h291: dout <= 8'b11101111; //  657 : 239 - 0xef
      12'h292: dout <= 8'b11110111; //  658 : 247 - 0xf7
      12'h293: dout <= 8'b11111111; //  659 : 255 - 0xff
      12'h294: dout <= 8'b11111111; //  660 : 255 - 0xff
      12'h295: dout <= 8'b11111110; //  661 : 254 - 0xfe
      12'h296: dout <= 8'b01111100; //  662 : 124 - 0x7c
      12'h297: dout <= 8'b01110000; //  663 : 112 - 0x70
      12'h298: dout <= 8'b11100000; //  664 : 224 - 0xe0 -- Sprite 0x53
      12'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout <= 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout <= 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout <= 8'b00100000; //  672 :  32 - 0x20 -- Sprite 0x54
      12'h2A1: dout <= 8'b01000000; //  673 :  64 - 0x40
      12'h2A2: dout <= 8'b10000000; //  674 : 128 - 0x80
      12'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      12'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      12'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      12'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      12'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout <= 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout <= 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout <= 8'b10000000; //  686 : 128 - 0x80
      12'h2AF: dout <= 8'b11000000; //  687 : 192 - 0xc0
      12'h2B0: dout <= 8'b11100000; //  688 : 224 - 0xe0 -- Sprite 0x56
      12'h2B1: dout <= 8'b11100000; //  689 : 224 - 0xe0
      12'h2B2: dout <= 8'b11100000; //  690 : 224 - 0xe0
      12'h2B3: dout <= 8'b11000000; //  691 : 192 - 0xc0
      12'h2B4: dout <= 8'b10000000; //  692 : 128 - 0x80
      12'h2B5: dout <= 8'b00000000; //  693 :   0 - 0x0
      12'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      12'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      12'h2C1: dout <= 8'b11111111; //  705 : 255 - 0xff
      12'h2C2: dout <= 8'b11111111; //  706 : 255 - 0xff
      12'h2C3: dout <= 8'b11111111; //  707 : 255 - 0xff
      12'h2C4: dout <= 8'b11111111; //  708 : 255 - 0xff
      12'h2C5: dout <= 8'b11111111; //  709 : 255 - 0xff
      12'h2C6: dout <= 8'b11111111; //  710 : 255 - 0xff
      12'h2C7: dout <= 8'b11111111; //  711 : 255 - 0xff
      12'h2C8: dout <= 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      12'h2C9: dout <= 8'b11111111; //  713 : 255 - 0xff
      12'h2CA: dout <= 8'b11111111; //  714 : 255 - 0xff
      12'h2CB: dout <= 8'b11111111; //  715 : 255 - 0xff
      12'h2CC: dout <= 8'b11111111; //  716 : 255 - 0xff
      12'h2CD: dout <= 8'b11111111; //  717 : 255 - 0xff
      12'h2CE: dout <= 8'b11111111; //  718 : 255 - 0xff
      12'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      12'h2D0: dout <= 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      12'h2D1: dout <= 8'b11111111; //  721 : 255 - 0xff
      12'h2D2: dout <= 8'b11111111; //  722 : 255 - 0xff
      12'h2D3: dout <= 8'b11111111; //  723 : 255 - 0xff
      12'h2D4: dout <= 8'b11111111; //  724 : 255 - 0xff
      12'h2D5: dout <= 8'b11111111; //  725 : 255 - 0xff
      12'h2D6: dout <= 8'b11111111; //  726 : 255 - 0xff
      12'h2D7: dout <= 8'b11111111; //  727 : 255 - 0xff
      12'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      12'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      12'h2DA: dout <= 8'b11111111; //  730 : 255 - 0xff
      12'h2DB: dout <= 8'b11111111; //  731 : 255 - 0xff
      12'h2DC: dout <= 8'b11111111; //  732 : 255 - 0xff
      12'h2DD: dout <= 8'b11111111; //  733 : 255 - 0xff
      12'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      12'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout <= 8'b11111111; //  736 : 255 - 0xff -- Sprite 0x5c
      12'h2E1: dout <= 8'b11111111; //  737 : 255 - 0xff
      12'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      12'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      12'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      12'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      12'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      12'h2E7: dout <= 8'b11111111; //  743 : 255 - 0xff
      12'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      12'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      12'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      12'h2EB: dout <= 8'b11111111; //  747 : 255 - 0xff
      12'h2EC: dout <= 8'b11111111; //  748 : 255 - 0xff
      12'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      12'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      12'h2EF: dout <= 8'b11111111; //  751 : 255 - 0xff
      12'h2F0: dout <= 8'b11111111; //  752 : 255 - 0xff -- Sprite 0x5e
      12'h2F1: dout <= 8'b11111111; //  753 : 255 - 0xff
      12'h2F2: dout <= 8'b11111111; //  754 : 255 - 0xff
      12'h2F3: dout <= 8'b11111111; //  755 : 255 - 0xff
      12'h2F4: dout <= 8'b11111111; //  756 : 255 - 0xff
      12'h2F5: dout <= 8'b11111111; //  757 : 255 - 0xff
      12'h2F6: dout <= 8'b11111111; //  758 : 255 - 0xff
      12'h2F7: dout <= 8'b11111111; //  759 : 255 - 0xff
      12'h2F8: dout <= 8'b11111111; //  760 : 255 - 0xff -- Sprite 0x5f
      12'h2F9: dout <= 8'b11111111; //  761 : 255 - 0xff
      12'h2FA: dout <= 8'b11111111; //  762 : 255 - 0xff
      12'h2FB: dout <= 8'b11111111; //  763 : 255 - 0xff
      12'h2FC: dout <= 8'b11111111; //  764 : 255 - 0xff
      12'h2FD: dout <= 8'b11111111; //  765 : 255 - 0xff
      12'h2FE: dout <= 8'b11111111; //  766 : 255 - 0xff
      12'h2FF: dout <= 8'b11111111; //  767 : 255 - 0xff
      12'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b00011111; //  770 :  31 - 0x1f
      12'h303: dout <= 8'b00111111; //  771 :  63 - 0x3f
      12'h304: dout <= 8'b00111111; //  772 :  63 - 0x3f
      12'h305: dout <= 8'b01111111; //  773 : 127 - 0x7f
      12'h306: dout <= 8'b01111111; //  774 : 127 - 0x7f
      12'h307: dout <= 8'b01111111; //  775 : 127 - 0x7f
      12'h308: dout <= 8'b01111111; //  776 : 127 - 0x7f -- Sprite 0x61
      12'h309: dout <= 8'b00111110; //  777 :  62 - 0x3e
      12'h30A: dout <= 8'b00011111; //  778 :  31 - 0x1f
      12'h30B: dout <= 8'b00011111; //  779 :  31 - 0x1f
      12'h30C: dout <= 8'b00001111; //  780 :  15 - 0xf
      12'h30D: dout <= 8'b00001111; //  781 :  15 - 0xf
      12'h30E: dout <= 8'b00001111; //  782 :  15 - 0xf
      12'h30F: dout <= 8'b00000111; //  783 :   7 - 0x7
      12'h310: dout <= 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      12'h311: dout <= 8'b01100000; //  785 :  96 - 0x60
      12'h312: dout <= 8'b11110000; //  786 : 240 - 0xf0
      12'h313: dout <= 8'b11111000; //  787 : 248 - 0xf8
      12'h314: dout <= 8'b11111000; //  788 : 248 - 0xf8
      12'h315: dout <= 8'b11111000; //  789 : 248 - 0xf8
      12'h316: dout <= 8'b11111100; //  790 : 252 - 0xfc
      12'h317: dout <= 8'b11111100; //  791 : 252 - 0xfc
      12'h318: dout <= 8'b11111000; //  792 : 248 - 0xf8 -- Sprite 0x63
      12'h319: dout <= 8'b11110000; //  793 : 240 - 0xf0
      12'h31A: dout <= 8'b11110000; //  794 : 240 - 0xf0
      12'h31B: dout <= 8'b11100000; //  795 : 224 - 0xe0
      12'h31C: dout <= 8'b10000000; //  796 : 128 - 0x80
      12'h31D: dout <= 8'b10000000; //  797 : 128 - 0x80
      12'h31E: dout <= 8'b11000000; //  798 : 192 - 0xc0
      12'h31F: dout <= 8'b11000000; //  799 : 192 - 0xc0
      12'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      12'h321: dout <= 8'b00011111; //  801 :  31 - 0x1f
      12'h322: dout <= 8'b00111111; //  802 :  63 - 0x3f
      12'h323: dout <= 8'b01111111; //  803 : 127 - 0x7f
      12'h324: dout <= 8'b11111111; //  804 : 255 - 0xff
      12'h325: dout <= 8'b11111111; //  805 : 255 - 0xff
      12'h326: dout <= 8'b00111110; //  806 :  62 - 0x3e
      12'h327: dout <= 8'b00001111; //  807 :  15 - 0xf
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b00000001; //  811 :   1 - 0x1
      12'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      12'h331: dout <= 8'b11100000; //  817 : 224 - 0xe0
      12'h332: dout <= 8'b11110000; //  818 : 240 - 0xf0
      12'h333: dout <= 8'b11111100; //  819 : 252 - 0xfc
      12'h334: dout <= 8'b11111110; //  820 : 254 - 0xfe
      12'h335: dout <= 8'b11111110; //  821 : 254 - 0xfe
      12'h336: dout <= 8'b11111111; //  822 : 255 - 0xff
      12'h337: dout <= 8'b11111100; //  823 : 252 - 0xfc
      12'h338: dout <= 8'b01111100; //  824 : 124 - 0x7c -- Sprite 0x67
      12'h339: dout <= 8'b11111100; //  825 : 252 - 0xfc
      12'h33A: dout <= 8'b11111000; //  826 : 248 - 0xf8
      12'h33B: dout <= 8'b11110000; //  827 : 240 - 0xf0
      12'h33C: dout <= 8'b11100000; //  828 : 224 - 0xe0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout <= 8'b00000111; //  833 :   7 - 0x7
      12'h342: dout <= 8'b00000111; //  834 :   7 - 0x7
      12'h343: dout <= 8'b00001111; //  835 :  15 - 0xf
      12'h344: dout <= 8'b00001111; //  836 :  15 - 0xf
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00011111; //  838 :  31 - 0x1f
      12'h347: dout <= 8'b00111111; //  839 :  63 - 0x3f
      12'h348: dout <= 8'b01111111; //  840 : 127 - 0x7f -- Sprite 0x69
      12'h349: dout <= 8'b01111111; //  841 : 127 - 0x7f
      12'h34A: dout <= 8'b00011111; //  842 :  31 - 0x1f
      12'h34B: dout <= 8'b00011111; //  843 :  31 - 0x1f
      12'h34C: dout <= 8'b00011111; //  844 :  31 - 0x1f
      12'h34D: dout <= 8'b00011110; //  845 :  30 - 0x1e
      12'h34E: dout <= 8'b00001111; //  846 :  15 - 0xf
      12'h34F: dout <= 8'b00011111; //  847 :  31 - 0x1f
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout <= 8'b11100000; //  849 : 224 - 0xe0
      12'h352: dout <= 8'b11100000; //  850 : 224 - 0xe0
      12'h353: dout <= 8'b11110000; //  851 : 240 - 0xf0
      12'h354: dout <= 8'b11110000; //  852 : 240 - 0xf0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b11111000; //  854 : 248 - 0xf8
      12'h357: dout <= 8'b11111100; //  855 : 252 - 0xfc
      12'h358: dout <= 8'b11111110; //  856 : 254 - 0xfe -- Sprite 0x6b
      12'h359: dout <= 8'b11111110; //  857 : 254 - 0xfe
      12'h35A: dout <= 8'b11111000; //  858 : 248 - 0xf8
      12'h35B: dout <= 8'b11111000; //  859 : 248 - 0xf8
      12'h35C: dout <= 8'b11111000; //  860 : 248 - 0xf8
      12'h35D: dout <= 8'b01111000; //  861 : 120 - 0x78
      12'h35E: dout <= 8'b11110000; //  862 : 240 - 0xf0
      12'h35F: dout <= 8'b11111000; //  863 : 248 - 0xf8
      12'h360: dout <= 8'b00000011; //  864 :   3 - 0x3 -- Sprite 0x6c
      12'h361: dout <= 8'b00000111; //  865 :   7 - 0x7
      12'h362: dout <= 8'b00000101; //  866 :   5 - 0x5
      12'h363: dout <= 8'b00001000; //  867 :   8 - 0x8
      12'h364: dout <= 8'b00011011; //  868 :  27 - 0x1b
      12'h365: dout <= 8'b00011001; //  869 :  25 - 0x19
      12'h366: dout <= 8'b00000101; //  870 :   5 - 0x5
      12'h367: dout <= 8'b00111111; //  871 :  63 - 0x3f
      12'h368: dout <= 8'b00111111; //  872 :  63 - 0x3f -- Sprite 0x6d
      12'h369: dout <= 8'b00001111; //  873 :  15 - 0xf
      12'h36A: dout <= 8'b00000101; //  874 :   5 - 0x5
      12'h36B: dout <= 8'b00110111; //  875 :  55 - 0x37
      12'h36C: dout <= 8'b00111111; //  876 :  63 - 0x3f
      12'h36D: dout <= 8'b00111111; //  877 :  63 - 0x3f
      12'h36E: dout <= 8'b00111110; //  878 :  62 - 0x3e
      12'h36F: dout <= 8'b00011100; //  879 :  28 - 0x1c
      12'h370: dout <= 8'b11100000; //  880 : 224 - 0xe0 -- Sprite 0x6e
      12'h371: dout <= 8'b11110000; //  881 : 240 - 0xf0
      12'h372: dout <= 8'b01010000; //  882 :  80 - 0x50
      12'h373: dout <= 8'b00001000; //  883 :   8 - 0x8
      12'h374: dout <= 8'b01101100; //  884 : 108 - 0x6c
      12'h375: dout <= 8'b11001100; //  885 : 204 - 0xcc
      12'h376: dout <= 8'b11010000; //  886 : 208 - 0xd0
      12'h377: dout <= 8'b11111110; //  887 : 254 - 0xfe
      12'h378: dout <= 8'b11111110; //  888 : 254 - 0xfe -- Sprite 0x6f
      12'h379: dout <= 8'b11111000; //  889 : 248 - 0xf8
      12'h37A: dout <= 8'b11010000; //  890 : 208 - 0xd0
      12'h37B: dout <= 8'b11111011; //  891 : 251 - 0xfb
      12'h37C: dout <= 8'b11111111; //  892 : 255 - 0xff
      12'h37D: dout <= 8'b11111111; //  893 : 255 - 0xff
      12'h37E: dout <= 8'b00111110; //  894 :  62 - 0x3e
      12'h37F: dout <= 8'b00001100; //  895 :  12 - 0xc
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      12'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout <= 8'b01111001; //  898 : 121 - 0x79
      12'h383: dout <= 8'b11111001; //  899 : 249 - 0xf9
      12'h384: dout <= 8'b11110011; //  900 : 243 - 0xf3
      12'h385: dout <= 8'b11111111; //  901 : 255 - 0xff
      12'h386: dout <= 8'b01111011; //  902 : 123 - 0x7b
      12'h387: dout <= 8'b00111111; //  903 :  63 - 0x3f
      12'h388: dout <= 8'b00111111; //  904 :  63 - 0x3f -- Sprite 0x71
      12'h389: dout <= 8'b00111111; //  905 :  63 - 0x3f
      12'h38A: dout <= 8'b01111011; //  906 : 123 - 0x7b
      12'h38B: dout <= 8'b01111111; //  907 : 127 - 0x7f
      12'h38C: dout <= 8'b11111011; //  908 : 251 - 0xfb
      12'h38D: dout <= 8'b11110001; //  909 : 241 - 0xf1
      12'h38E: dout <= 8'b01111001; //  910 : 121 - 0x79
      12'h38F: dout <= 8'b00111000; //  911 :  56 - 0x38
      12'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      12'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout <= 8'b10000000; //  914 : 128 - 0x80
      12'h393: dout <= 8'b10110000; //  915 : 176 - 0xb0
      12'h394: dout <= 8'b10111000; //  916 : 184 - 0xb8
      12'h395: dout <= 8'b11000110; //  917 : 198 - 0xc6
      12'h396: dout <= 8'b10010011; //  918 : 147 - 0x93
      12'h397: dout <= 8'b11110111; //  919 : 247 - 0xf7
      12'h398: dout <= 8'b11100011; //  920 : 227 - 0xe3 -- Sprite 0x73
      12'h399: dout <= 8'b11110111; //  921 : 247 - 0xf7
      12'h39A: dout <= 8'b10010011; //  922 : 147 - 0x93
      12'h39B: dout <= 8'b11000110; //  923 : 198 - 0xc6
      12'h39C: dout <= 8'b10111000; //  924 : 184 - 0xb8
      12'h39D: dout <= 8'b10110000; //  925 : 176 - 0xb0
      12'h39E: dout <= 8'b10000000; //  926 : 128 - 0x80
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00110000; //  928 :  48 - 0x30 -- Sprite 0x74
      12'h3A1: dout <= 8'b01111100; //  929 : 124 - 0x7c
      12'h3A2: dout <= 8'b11111111; //  930 : 255 - 0xff
      12'h3A3: dout <= 8'b11111111; //  931 : 255 - 0xff
      12'h3A4: dout <= 8'b11011111; //  932 : 223 - 0xdf
      12'h3A5: dout <= 8'b00001011; //  933 :  11 - 0xb
      12'h3A6: dout <= 8'b00011111; //  934 :  31 - 0x1f
      12'h3A7: dout <= 8'b01111111; //  935 : 127 - 0x7f
      12'h3A8: dout <= 8'b01111111; //  936 : 127 - 0x7f -- Sprite 0x75
      12'h3A9: dout <= 8'b00001011; //  937 :  11 - 0xb
      12'h3AA: dout <= 8'b00110011; //  938 :  51 - 0x33
      12'h3AB: dout <= 8'b00110110; //  939 :  54 - 0x36
      12'h3AC: dout <= 8'b00010000; //  940 :  16 - 0x10
      12'h3AD: dout <= 8'b00001010; //  941 :  10 - 0xa
      12'h3AE: dout <= 8'b00001111; //  942 :  15 - 0xf
      12'h3AF: dout <= 8'b00000111; //  943 :   7 - 0x7
      12'h3B0: dout <= 8'b00111000; //  944 :  56 - 0x38 -- Sprite 0x76
      12'h3B1: dout <= 8'b01111100; //  945 : 124 - 0x7c
      12'h3B2: dout <= 8'b11111100; //  946 : 252 - 0xfc
      12'h3B3: dout <= 8'b11111100; //  947 : 252 - 0xfc
      12'h3B4: dout <= 8'b11101100; //  948 : 236 - 0xec
      12'h3B5: dout <= 8'b10100000; //  949 : 160 - 0xa0
      12'h3B6: dout <= 8'b11110000; //  950 : 240 - 0xf0
      12'h3B7: dout <= 8'b11111100; //  951 : 252 - 0xfc
      12'h3B8: dout <= 8'b11111100; //  952 : 252 - 0xfc -- Sprite 0x77
      12'h3B9: dout <= 8'b10100000; //  953 : 160 - 0xa0
      12'h3BA: dout <= 8'b10011000; //  954 : 152 - 0x98
      12'h3BB: dout <= 8'b11011000; //  955 : 216 - 0xd8
      12'h3BC: dout <= 8'b00010000; //  956 :  16 - 0x10
      12'h3BD: dout <= 8'b10100000; //  957 : 160 - 0xa0
      12'h3BE: dout <= 8'b11100000; //  958 : 224 - 0xe0
      12'h3BF: dout <= 8'b11000000; //  959 : 192 - 0xc0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout <= 8'b00000001; //  961 :   1 - 0x1
      12'h3C2: dout <= 8'b00001101; //  962 :  13 - 0xd
      12'h3C3: dout <= 8'b00011101; //  963 :  29 - 0x1d
      12'h3C4: dout <= 8'b01100011; //  964 :  99 - 0x63
      12'h3C5: dout <= 8'b11001001; //  965 : 201 - 0xc9
      12'h3C6: dout <= 8'b11101111; //  966 : 239 - 0xef
      12'h3C7: dout <= 8'b11000111; //  967 : 199 - 0xc7
      12'h3C8: dout <= 8'b11101111; //  968 : 239 - 0xef -- Sprite 0x79
      12'h3C9: dout <= 8'b11001001; //  969 : 201 - 0xc9
      12'h3CA: dout <= 8'b01100011; //  970 :  99 - 0x63
      12'h3CB: dout <= 8'b00011101; //  971 :  29 - 0x1d
      12'h3CC: dout <= 8'b00001101; //  972 :  13 - 0xd
      12'h3CD: dout <= 8'b00000001; //  973 :   1 - 0x1
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00011100; //  976 :  28 - 0x1c -- Sprite 0x7a
      12'h3D1: dout <= 8'b10011110; //  977 : 158 - 0x9e
      12'h3D2: dout <= 8'b10001111; //  978 : 143 - 0x8f
      12'h3D3: dout <= 8'b11011111; //  979 : 223 - 0xdf
      12'h3D4: dout <= 8'b11111110; //  980 : 254 - 0xfe
      12'h3D5: dout <= 8'b11011110; //  981 : 222 - 0xde
      12'h3D6: dout <= 8'b11111100; //  982 : 252 - 0xfc
      12'h3D7: dout <= 8'b11111100; //  983 : 252 - 0xfc
      12'h3D8: dout <= 8'b11111100; //  984 : 252 - 0xfc -- Sprite 0x7b
      12'h3D9: dout <= 8'b11011110; //  985 : 222 - 0xde
      12'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      12'h3DB: dout <= 8'b11001111; //  987 : 207 - 0xcf
      12'h3DC: dout <= 8'b10011111; //  988 : 159 - 0x9f
      12'h3DD: dout <= 8'b10011110; //  989 : 158 - 0x9e
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout <= 8'b00011110; //  996 :  30 - 0x1e
      12'h3E5: dout <= 8'b00111111; //  997 :  63 - 0x3f
      12'h3E6: dout <= 8'b01111101; //  998 : 125 - 0x7d
      12'h3E7: dout <= 8'b01111000; //  999 : 120 - 0x78
      12'h3E8: dout <= 8'b01111100; // 1000 : 124 - 0x7c -- Sprite 0x7d
      12'h3E9: dout <= 8'b11111011; // 1001 : 251 - 0xfb
      12'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      12'h3EC: dout <= 8'b01011111; // 1004 :  95 - 0x5f
      12'h3ED: dout <= 8'b00011111; // 1005 :  31 - 0x1f
      12'h3EE: dout <= 8'b00011111; // 1006 :  31 - 0x1f
      12'h3EF: dout <= 8'b00011111; // 1007 :  31 - 0x1f
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout <= 8'b10000000; // 1013 : 128 - 0x80
      12'h3F6: dout <= 8'b10000000; // 1014 : 128 - 0x80
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      12'h3F9: dout <= 8'b00100001; // 1017 :  33 - 0x21
      12'h3FA: dout <= 8'b10100010; // 1018 : 162 - 0xa2
      12'h3FB: dout <= 8'b10100011; // 1019 : 163 - 0xa3
      12'h3FC: dout <= 8'b10110011; // 1020 : 179 - 0xb3
      12'h3FD: dout <= 8'b10001111; // 1021 : 143 - 0x8f
      12'h3FE: dout <= 8'b00100111; // 1022 :  39 - 0x27
      12'h3FF: dout <= 8'b11111110; // 1023 : 254 - 0xfe
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      12'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000011; // 1028 :   3 - 0x3
      12'h405: dout <= 8'b00001111; // 1029 :  15 - 0xf
      12'h406: dout <= 8'b00011111; // 1030 :  31 - 0x1f
      12'h407: dout <= 8'b00011111; // 1031 :  31 - 0x1f
      12'h408: dout <= 8'b00011111; // 1032 :  31 - 0x1f -- Sprite 0x81
      12'h409: dout <= 8'b00011111; // 1033 :  31 - 0x1f
      12'h40A: dout <= 8'b00001111; // 1034 :  15 - 0xf
      12'h40B: dout <= 8'b00000011; // 1035 :   3 - 0x3
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      12'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout <= 8'b11000000; // 1044 : 192 - 0xc0
      12'h415: dout <= 8'b11110000; // 1045 : 240 - 0xf0
      12'h416: dout <= 8'b11111000; // 1046 : 248 - 0xf8
      12'h417: dout <= 8'b11111000; // 1047 : 248 - 0xf8
      12'h418: dout <= 8'b11111000; // 1048 : 248 - 0xf8 -- Sprite 0x83
      12'h419: dout <= 8'b11111000; // 1049 : 248 - 0xf8
      12'h41A: dout <= 8'b11110000; // 1050 : 240 - 0xf0
      12'h41B: dout <= 8'b11000000; // 1051 : 192 - 0xc0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      12'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      12'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      12'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout <= 8'b00000011; // 1060 :   3 - 0x3
      12'h425: dout <= 8'b00001111; // 1061 :  15 - 0xf
      12'h426: dout <= 8'b00011111; // 1062 :  31 - 0x1f
      12'h427: dout <= 8'b00011111; // 1063 :  31 - 0x1f
      12'h428: dout <= 8'b00011111; // 1064 :  31 - 0x1f -- Sprite 0x85
      12'h429: dout <= 8'b00011111; // 1065 :  31 - 0x1f
      12'h42A: dout <= 8'b00001111; // 1066 :  15 - 0xf
      12'h42B: dout <= 8'b00000011; // 1067 :   3 - 0x3
      12'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b11000000; // 1076 : 192 - 0xc0
      12'h435: dout <= 8'b11110000; // 1077 : 240 - 0xf0
      12'h436: dout <= 8'b11111000; // 1078 : 248 - 0xf8
      12'h437: dout <= 8'b11111000; // 1079 : 248 - 0xf8
      12'h438: dout <= 8'b11111000; // 1080 : 248 - 0xf8 -- Sprite 0x87
      12'h439: dout <= 8'b11111000; // 1081 : 248 - 0xf8
      12'h43A: dout <= 8'b11110000; // 1082 : 240 - 0xf0
      12'h43B: dout <= 8'b11000000; // 1083 : 192 - 0xc0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      12'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      12'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      12'h443: dout <= 8'b00000000; // 1091 :   0 - 0x0
      12'h444: dout <= 8'b00000011; // 1092 :   3 - 0x3
      12'h445: dout <= 8'b00001111; // 1093 :  15 - 0xf
      12'h446: dout <= 8'b00011111; // 1094 :  31 - 0x1f
      12'h447: dout <= 8'b00011111; // 1095 :  31 - 0x1f
      12'h448: dout <= 8'b00011111; // 1096 :  31 - 0x1f -- Sprite 0x89
      12'h449: dout <= 8'b00011111; // 1097 :  31 - 0x1f
      12'h44A: dout <= 8'b00001111; // 1098 :  15 - 0xf
      12'h44B: dout <= 8'b00000011; // 1099 :   3 - 0x3
      12'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      12'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      12'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      12'h453: dout <= 8'b00000000; // 1107 :   0 - 0x0
      12'h454: dout <= 8'b11000000; // 1108 : 192 - 0xc0
      12'h455: dout <= 8'b11110000; // 1109 : 240 - 0xf0
      12'h456: dout <= 8'b11111000; // 1110 : 248 - 0xf8
      12'h457: dout <= 8'b11111000; // 1111 : 248 - 0xf8
      12'h458: dout <= 8'b11111000; // 1112 : 248 - 0xf8 -- Sprite 0x8b
      12'h459: dout <= 8'b11111000; // 1113 : 248 - 0xf8
      12'h45A: dout <= 8'b11110000; // 1114 : 240 - 0xf0
      12'h45B: dout <= 8'b11000000; // 1115 : 192 - 0xc0
      12'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      12'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      12'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      12'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      12'h464: dout <= 8'b00000011; // 1124 :   3 - 0x3
      12'h465: dout <= 8'b00001111; // 1125 :  15 - 0xf
      12'h466: dout <= 8'b00011111; // 1126 :  31 - 0x1f
      12'h467: dout <= 8'b00011111; // 1127 :  31 - 0x1f
      12'h468: dout <= 8'b00011111; // 1128 :  31 - 0x1f -- Sprite 0x8d
      12'h469: dout <= 8'b00011111; // 1129 :  31 - 0x1f
      12'h46A: dout <= 8'b00001111; // 1130 :  15 - 0xf
      12'h46B: dout <= 8'b00000011; // 1131 :   3 - 0x3
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      12'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      12'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout <= 8'b11000000; // 1140 : 192 - 0xc0
      12'h475: dout <= 8'b11110000; // 1141 : 240 - 0xf0
      12'h476: dout <= 8'b11111000; // 1142 : 248 - 0xf8
      12'h477: dout <= 8'b11111000; // 1143 : 248 - 0xf8
      12'h478: dout <= 8'b11111000; // 1144 : 248 - 0xf8 -- Sprite 0x8f
      12'h479: dout <= 8'b11111000; // 1145 : 248 - 0xf8
      12'h47A: dout <= 8'b11110000; // 1146 : 240 - 0xf0
      12'h47B: dout <= 8'b11000000; // 1147 : 192 - 0xc0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b00001111; // 1155 :  15 - 0xf
      12'h484: dout <= 8'b00110000; // 1156 :  48 - 0x30
      12'h485: dout <= 8'b01100000; // 1157 :  96 - 0x60
      12'h486: dout <= 8'b00111111; // 1158 :  63 - 0x3f
      12'h487: dout <= 8'b01111111; // 1159 : 127 - 0x7f
      12'h488: dout <= 8'b01111111; // 1160 : 127 - 0x7f -- Sprite 0x91
      12'h489: dout <= 8'b00111111; // 1161 :  63 - 0x3f
      12'h48A: dout <= 8'b01100000; // 1162 :  96 - 0x60
      12'h48B: dout <= 8'b00110000; // 1163 :  48 - 0x30
      12'h48C: dout <= 8'b00001111; // 1164 :  15 - 0xf
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      12'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      12'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout <= 8'b11111000; // 1171 : 248 - 0xf8
      12'h494: dout <= 8'b00000110; // 1172 :   6 - 0x6
      12'h495: dout <= 8'b00000011; // 1173 :   3 - 0x3
      12'h496: dout <= 8'b11111110; // 1174 : 254 - 0xfe
      12'h497: dout <= 8'b11111111; // 1175 : 255 - 0xff
      12'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- Sprite 0x93
      12'h499: dout <= 8'b11111110; // 1177 : 254 - 0xfe
      12'h49A: dout <= 8'b00000011; // 1178 :   3 - 0x3
      12'h49B: dout <= 8'b00000110; // 1179 :   6 - 0x6
      12'h49C: dout <= 8'b11111000; // 1180 : 248 - 0xf8
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      12'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout <= 8'b00101111; // 1188 :  47 - 0x2f
      12'h4A5: dout <= 8'b00111111; // 1189 :  63 - 0x3f
      12'h4A6: dout <= 8'b01100000; // 1190 :  96 - 0x60
      12'h4A7: dout <= 8'b00100000; // 1191 :  32 - 0x20
      12'h4A8: dout <= 8'b00100000; // 1192 :  32 - 0x20 -- Sprite 0x95
      12'h4A9: dout <= 8'b01100000; // 1193 :  96 - 0x60
      12'h4AA: dout <= 8'b00111111; // 1194 :  63 - 0x3f
      12'h4AB: dout <= 8'b00101111; // 1195 :  47 - 0x2f
      12'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      12'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout <= 8'b11111010; // 1204 : 250 - 0xfa
      12'h4B5: dout <= 8'b11111110; // 1205 : 254 - 0xfe
      12'h4B6: dout <= 8'b00000011; // 1206 :   3 - 0x3
      12'h4B7: dout <= 8'b00000010; // 1207 :   2 - 0x2
      12'h4B8: dout <= 8'b00000010; // 1208 :   2 - 0x2 -- Sprite 0x97
      12'h4B9: dout <= 8'b00000011; // 1209 :   3 - 0x3
      12'h4BA: dout <= 8'b11111110; // 1210 : 254 - 0xfe
      12'h4BB: dout <= 8'b11111010; // 1211 : 250 - 0xfa
      12'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      12'h4C1: dout <= 8'b01000100; // 1217 :  68 - 0x44
      12'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout <= 8'b01000001; // 1219 :  65 - 0x41
      12'h4C4: dout <= 8'b00100000; // 1220 :  32 - 0x20
      12'h4C5: dout <= 8'b01001011; // 1221 :  75 - 0x4b
      12'h4C6: dout <= 8'b00100111; // 1222 :  39 - 0x27
      12'h4C7: dout <= 8'b00011111; // 1223 :  31 - 0x1f
      12'h4C8: dout <= 8'b00001111; // 1224 :  15 - 0xf -- Sprite 0x99
      12'h4C9: dout <= 8'b00011110; // 1225 :  30 - 0x1e
      12'h4CA: dout <= 8'b00011111; // 1226 :  31 - 0x1f
      12'h4CB: dout <= 8'b00011111; // 1227 :  31 - 0x1f
      12'h4CC: dout <= 8'b00011111; // 1228 :  31 - 0x1f
      12'h4CD: dout <= 8'b00001111; // 1229 :  15 - 0xf
      12'h4CE: dout <= 8'b00001111; // 1230 :  15 - 0xf
      12'h4CF: dout <= 8'b00000011; // 1231 :   3 - 0x3
      12'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout <= 8'b00100000; // 1233 :  32 - 0x20
      12'h4D2: dout <= 8'b01010000; // 1234 :  80 - 0x50
      12'h4D3: dout <= 8'b00100000; // 1235 :  32 - 0x20
      12'h4D4: dout <= 8'b01100000; // 1236 :  96 - 0x60
      12'h4D5: dout <= 8'b01001000; // 1237 :  72 - 0x48
      12'h4D6: dout <= 8'b11100000; // 1238 : 224 - 0xe0
      12'h4D7: dout <= 8'b11110000; // 1239 : 240 - 0xf0
      12'h4D8: dout <= 8'b11111000; // 1240 : 248 - 0xf8 -- Sprite 0x9b
      12'h4D9: dout <= 8'b01111000; // 1241 : 120 - 0x78
      12'h4DA: dout <= 8'b00111100; // 1242 :  60 - 0x3c
      12'h4DB: dout <= 8'b00111100; // 1243 :  60 - 0x3c
      12'h4DC: dout <= 8'b00111100; // 1244 :  60 - 0x3c
      12'h4DD: dout <= 8'b11111100; // 1245 : 252 - 0xfc
      12'h4DE: dout <= 8'b11111000; // 1246 : 248 - 0xf8
      12'h4DF: dout <= 8'b11100000; // 1247 : 224 - 0xe0
      12'h4E0: dout <= 8'b00010000; // 1248 :  16 - 0x10 -- Sprite 0x9c
      12'h4E1: dout <= 8'b00000001; // 1249 :   1 - 0x1
      12'h4E2: dout <= 8'b00101010; // 1250 :  42 - 0x2a
      12'h4E3: dout <= 8'b00001100; // 1251 :  12 - 0xc
      12'h4E4: dout <= 8'b10100110; // 1252 : 166 - 0xa6
      12'h4E5: dout <= 8'b00010111; // 1253 :  23 - 0x17
      12'h4E6: dout <= 8'b00011111; // 1254 :  31 - 0x1f
      12'h4E7: dout <= 8'b00011111; // 1255 :  31 - 0x1f
      12'h4E8: dout <= 8'b01011110; // 1256 :  94 - 0x5e -- Sprite 0x9d
      12'h4E9: dout <= 8'b00111100; // 1257 :  60 - 0x3c
      12'h4EA: dout <= 8'b00111101; // 1258 :  61 - 0x3d
      12'h4EB: dout <= 8'b00111101; // 1259 :  61 - 0x3d
      12'h4EC: dout <= 8'b00111110; // 1260 :  62 - 0x3e
      12'h4ED: dout <= 8'b00011111; // 1261 :  31 - 0x1f
      12'h4EE: dout <= 8'b00001111; // 1262 :  15 - 0xf
      12'h4EF: dout <= 8'b00000111; // 1263 :   7 - 0x7
      12'h4F0: dout <= 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      12'h4F1: dout <= 8'b00000000; // 1265 :   0 - 0x0
      12'h4F2: dout <= 8'b10000000; // 1266 : 128 - 0x80
      12'h4F3: dout <= 8'b11001000; // 1267 : 200 - 0xc8
      12'h4F4: dout <= 8'b01100000; // 1268 :  96 - 0x60
      12'h4F5: dout <= 8'b11100000; // 1269 : 224 - 0xe0
      12'h4F6: dout <= 8'b11110100; // 1270 : 244 - 0xf4
      12'h4F7: dout <= 8'b11111000; // 1271 : 248 - 0xf8
      12'h4F8: dout <= 8'b01111100; // 1272 : 124 - 0x7c -- Sprite 0x9f
      12'h4F9: dout <= 8'b00011100; // 1273 :  28 - 0x1c
      12'h4FA: dout <= 8'b00101110; // 1274 :  46 - 0x2e
      12'h4FB: dout <= 8'b00101110; // 1275 :  46 - 0x2e
      12'h4FC: dout <= 8'b00011110; // 1276 :  30 - 0x1e
      12'h4FD: dout <= 8'b11111100; // 1277 : 252 - 0xfc
      12'h4FE: dout <= 8'b11111000; // 1278 : 248 - 0xf8
      12'h4FF: dout <= 8'b11100000; // 1279 : 224 - 0xe0
      12'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0xa0
      12'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      12'h502: dout <= 8'b00111000; // 1282 :  56 - 0x38
      12'h503: dout <= 8'b01101100; // 1283 : 108 - 0x6c
      12'h504: dout <= 8'b11000110; // 1284 : 198 - 0xc6
      12'h505: dout <= 8'b10000011; // 1285 : 131 - 0x83
      12'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      12'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      12'h508: dout <= 8'b11111111; // 1288 : 255 - 0xff -- Sprite 0xa1
      12'h509: dout <= 8'b11111111; // 1289 : 255 - 0xff
      12'h50A: dout <= 8'b00111000; // 1290 :  56 - 0x38
      12'h50B: dout <= 8'b01101100; // 1291 : 108 - 0x6c
      12'h50C: dout <= 8'b11000110; // 1292 : 198 - 0xc6
      12'h50D: dout <= 8'b10000011; // 1293 : 131 - 0x83
      12'h50E: dout <= 8'b11111111; // 1294 : 255 - 0xff
      12'h50F: dout <= 8'b11111111; // 1295 : 255 - 0xff
      12'h510: dout <= 8'b10010010; // 1296 : 146 - 0x92 -- Sprite 0xa2
      12'h511: dout <= 8'b01010100; // 1297 :  84 - 0x54
      12'h512: dout <= 8'b00111000; // 1298 :  56 - 0x38
      12'h513: dout <= 8'b11111110; // 1299 : 254 - 0xfe
      12'h514: dout <= 8'b00111000; // 1300 :  56 - 0x38
      12'h515: dout <= 8'b01010100; // 1301 :  84 - 0x54
      12'h516: dout <= 8'b10010010; // 1302 : 146 - 0x92
      12'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout <= 8'b11111111; // 1304 : 255 - 0xff -- Sprite 0xa3
      12'h519: dout <= 8'b11111111; // 1305 : 255 - 0xff
      12'h51A: dout <= 8'b11111111; // 1306 : 255 - 0xff
      12'h51B: dout <= 8'b11111111; // 1307 : 255 - 0xff
      12'h51C: dout <= 8'b11111111; // 1308 : 255 - 0xff
      12'h51D: dout <= 8'b11111111; // 1309 : 255 - 0xff
      12'h51E: dout <= 8'b11111111; // 1310 : 255 - 0xff
      12'h51F: dout <= 8'b11111111; // 1311 : 255 - 0xff
      12'h520: dout <= 8'b11111111; // 1312 : 255 - 0xff -- Sprite 0xa4
      12'h521: dout <= 8'b11111111; // 1313 : 255 - 0xff
      12'h522: dout <= 8'b11111111; // 1314 : 255 - 0xff
      12'h523: dout <= 8'b11111111; // 1315 : 255 - 0xff
      12'h524: dout <= 8'b11111111; // 1316 : 255 - 0xff
      12'h525: dout <= 8'b11111111; // 1317 : 255 - 0xff
      12'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      12'h527: dout <= 8'b11111111; // 1319 : 255 - 0xff
      12'h528: dout <= 8'b11111111; // 1320 : 255 - 0xff -- Sprite 0xa5
      12'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      12'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      12'h52B: dout <= 8'b11111111; // 1323 : 255 - 0xff
      12'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      12'h52D: dout <= 8'b11111111; // 1325 : 255 - 0xff
      12'h52E: dout <= 8'b11111111; // 1326 : 255 - 0xff
      12'h52F: dout <= 8'b11111111; // 1327 : 255 - 0xff
      12'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0xa6
      12'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      12'h532: dout <= 8'b11111111; // 1330 : 255 - 0xff
      12'h533: dout <= 8'b11111111; // 1331 : 255 - 0xff
      12'h534: dout <= 8'b11111111; // 1332 : 255 - 0xff
      12'h535: dout <= 8'b11111111; // 1333 : 255 - 0xff
      12'h536: dout <= 8'b11111111; // 1334 : 255 - 0xff
      12'h537: dout <= 8'b11111111; // 1335 : 255 - 0xff
      12'h538: dout <= 8'b11111111; // 1336 : 255 - 0xff -- Sprite 0xa7
      12'h539: dout <= 8'b11111111; // 1337 : 255 - 0xff
      12'h53A: dout <= 8'b11111111; // 1338 : 255 - 0xff
      12'h53B: dout <= 8'b11111111; // 1339 : 255 - 0xff
      12'h53C: dout <= 8'b11111111; // 1340 : 255 - 0xff
      12'h53D: dout <= 8'b11111111; // 1341 : 255 - 0xff
      12'h53E: dout <= 8'b11111111; // 1342 : 255 - 0xff
      12'h53F: dout <= 8'b11111111; // 1343 : 255 - 0xff
      12'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      12'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout <= 8'b00100011; // 1349 :  35 - 0x23
      12'h546: dout <= 8'b10010111; // 1350 : 151 - 0x97
      12'h547: dout <= 8'b00101111; // 1351 :  47 - 0x2f
      12'h548: dout <= 8'b01101110; // 1352 : 110 - 0x6e -- Sprite 0xa9
      12'h549: dout <= 8'b11101111; // 1353 : 239 - 0xef
      12'h54A: dout <= 8'b11110111; // 1354 : 247 - 0xf7
      12'h54B: dout <= 8'b11111111; // 1355 : 255 - 0xff
      12'h54C: dout <= 8'b01111111; // 1356 : 127 - 0x7f
      12'h54D: dout <= 8'b00111111; // 1357 :  63 - 0x3f
      12'h54E: dout <= 8'b01011111; // 1358 :  95 - 0x5f
      12'h54F: dout <= 8'b00001111; // 1359 :  15 - 0xf
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout <= 8'b11111000; // 1364 : 248 - 0xf8
      12'h555: dout <= 8'b11111100; // 1365 : 252 - 0xfc
      12'h556: dout <= 8'b11111110; // 1366 : 254 - 0xfe
      12'h557: dout <= 8'b01011110; // 1367 :  94 - 0x5e
      12'h558: dout <= 8'b01011110; // 1368 :  94 - 0x5e -- Sprite 0xab
      12'h559: dout <= 8'b00001100; // 1369 :  12 - 0xc
      12'h55A: dout <= 8'b10011110; // 1370 : 158 - 0x9e
      12'h55B: dout <= 8'b11111110; // 1371 : 254 - 0xfe
      12'h55C: dout <= 8'b11111110; // 1372 : 254 - 0xfe
      12'h55D: dout <= 8'b11111110; // 1373 : 254 - 0xfe
      12'h55E: dout <= 8'b11111000; // 1374 : 248 - 0xf8
      12'h55F: dout <= 8'b11000000; // 1375 : 192 - 0xc0
      12'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout <= 8'b00000011; // 1381 :   3 - 0x3
      12'h566: dout <= 8'b00000111; // 1382 :   7 - 0x7
      12'h567: dout <= 8'b00101111; // 1383 :  47 - 0x2f
      12'h568: dout <= 8'b01001110; // 1384 :  78 - 0x4e -- Sprite 0xad
      12'h569: dout <= 8'b01101110; // 1385 : 110 - 0x6e
      12'h56A: dout <= 8'b11111110; // 1386 : 254 - 0xfe
      12'h56B: dout <= 8'b01111111; // 1387 : 127 - 0x7f
      12'h56C: dout <= 8'b00111111; // 1388 :  63 - 0x3f
      12'h56D: dout <= 8'b00011111; // 1389 :  31 - 0x1f
      12'h56E: dout <= 8'b00001111; // 1390 :  15 - 0xf
      12'h56F: dout <= 8'b00000011; // 1391 :   3 - 0x3
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b11111000; // 1396 : 248 - 0xf8
      12'h575: dout <= 8'b11111100; // 1397 : 252 - 0xfc
      12'h576: dout <= 8'b11111110; // 1398 : 254 - 0xfe
      12'h577: dout <= 8'b01010110; // 1399 :  86 - 0x56
      12'h578: dout <= 8'b01010110; // 1400 :  86 - 0x56 -- Sprite 0xaf
      12'h579: dout <= 8'b00001100; // 1401 :  12 - 0xc
      12'h57A: dout <= 8'b00001110; // 1402 :  14 - 0xe
      12'h57B: dout <= 8'b00011111; // 1403 :  31 - 0x1f
      12'h57C: dout <= 8'b11111111; // 1404 : 255 - 0xff
      12'h57D: dout <= 8'b11111111; // 1405 : 255 - 0xff
      12'h57E: dout <= 8'b11111110; // 1406 : 254 - 0xfe
      12'h57F: dout <= 8'b11111000; // 1407 : 248 - 0xf8
      12'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0xb0
      12'h581: dout <= 8'b11111111; // 1409 : 255 - 0xff
      12'h582: dout <= 8'b11111111; // 1410 : 255 - 0xff
      12'h583: dout <= 8'b11111111; // 1411 : 255 - 0xff
      12'h584: dout <= 8'b11111111; // 1412 : 255 - 0xff
      12'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout <= 8'b11111111; // 1414 : 255 - 0xff
      12'h587: dout <= 8'b11111111; // 1415 : 255 - 0xff
      12'h588: dout <= 8'b11111111; // 1416 : 255 - 0xff -- Sprite 0xb1
      12'h589: dout <= 8'b11111111; // 1417 : 255 - 0xff
      12'h58A: dout <= 8'b11111111; // 1418 : 255 - 0xff
      12'h58B: dout <= 8'b11111111; // 1419 : 255 - 0xff
      12'h58C: dout <= 8'b11111111; // 1420 : 255 - 0xff
      12'h58D: dout <= 8'b11111111; // 1421 : 255 - 0xff
      12'h58E: dout <= 8'b11111111; // 1422 : 255 - 0xff
      12'h58F: dout <= 8'b11111111; // 1423 : 255 - 0xff
      12'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0xb2
      12'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      12'h592: dout <= 8'b11111111; // 1426 : 255 - 0xff
      12'h593: dout <= 8'b11111111; // 1427 : 255 - 0xff
      12'h594: dout <= 8'b11111111; // 1428 : 255 - 0xff
      12'h595: dout <= 8'b11111111; // 1429 : 255 - 0xff
      12'h596: dout <= 8'b11111111; // 1430 : 255 - 0xff
      12'h597: dout <= 8'b11111111; // 1431 : 255 - 0xff
      12'h598: dout <= 8'b11111111; // 1432 : 255 - 0xff -- Sprite 0xb3
      12'h599: dout <= 8'b11111111; // 1433 : 255 - 0xff
      12'h59A: dout <= 8'b11111111; // 1434 : 255 - 0xff
      12'h59B: dout <= 8'b11111111; // 1435 : 255 - 0xff
      12'h59C: dout <= 8'b11111111; // 1436 : 255 - 0xff
      12'h59D: dout <= 8'b11111111; // 1437 : 255 - 0xff
      12'h59E: dout <= 8'b11111111; // 1438 : 255 - 0xff
      12'h59F: dout <= 8'b11111111; // 1439 : 255 - 0xff
      12'h5A0: dout <= 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0xb4
      12'h5A1: dout <= 8'b11111111; // 1441 : 255 - 0xff
      12'h5A2: dout <= 8'b11111111; // 1442 : 255 - 0xff
      12'h5A3: dout <= 8'b11111111; // 1443 : 255 - 0xff
      12'h5A4: dout <= 8'b11111111; // 1444 : 255 - 0xff
      12'h5A5: dout <= 8'b11111111; // 1445 : 255 - 0xff
      12'h5A6: dout <= 8'b11111111; // 1446 : 255 - 0xff
      12'h5A7: dout <= 8'b11111111; // 1447 : 255 - 0xff
      12'h5A8: dout <= 8'b11111111; // 1448 : 255 - 0xff -- Sprite 0xb5
      12'h5A9: dout <= 8'b11111111; // 1449 : 255 - 0xff
      12'h5AA: dout <= 8'b11111111; // 1450 : 255 - 0xff
      12'h5AB: dout <= 8'b11111111; // 1451 : 255 - 0xff
      12'h5AC: dout <= 8'b11111111; // 1452 : 255 - 0xff
      12'h5AD: dout <= 8'b11111111; // 1453 : 255 - 0xff
      12'h5AE: dout <= 8'b11111111; // 1454 : 255 - 0xff
      12'h5AF: dout <= 8'b11111111; // 1455 : 255 - 0xff
      12'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0xb6
      12'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      12'h5B2: dout <= 8'b11111111; // 1458 : 255 - 0xff
      12'h5B3: dout <= 8'b11111111; // 1459 : 255 - 0xff
      12'h5B4: dout <= 8'b11111111; // 1460 : 255 - 0xff
      12'h5B5: dout <= 8'b11111111; // 1461 : 255 - 0xff
      12'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      12'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      12'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- Sprite 0xb7
      12'h5B9: dout <= 8'b11111111; // 1465 : 255 - 0xff
      12'h5BA: dout <= 8'b11111111; // 1466 : 255 - 0xff
      12'h5BB: dout <= 8'b11111111; // 1467 : 255 - 0xff
      12'h5BC: dout <= 8'b11111111; // 1468 : 255 - 0xff
      12'h5BD: dout <= 8'b11111111; // 1469 : 255 - 0xff
      12'h5BE: dout <= 8'b11111111; // 1470 : 255 - 0xff
      12'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      12'h5C1: dout <= 8'b00000111; // 1473 :   7 - 0x7
      12'h5C2: dout <= 8'b00001000; // 1474 :   8 - 0x8
      12'h5C3: dout <= 8'b00010000; // 1475 :  16 - 0x10
      12'h5C4: dout <= 8'b00010000; // 1476 :  16 - 0x10
      12'h5C5: dout <= 8'b00100000; // 1477 :  32 - 0x20
      12'h5C6: dout <= 8'b00100000; // 1478 :  32 - 0x20
      12'h5C7: dout <= 8'b00100000; // 1479 :  32 - 0x20
      12'h5C8: dout <= 8'b00011111; // 1480 :  31 - 0x1f -- Sprite 0xb9
      12'h5C9: dout <= 8'b00101111; // 1481 :  47 - 0x2f
      12'h5CA: dout <= 8'b00110111; // 1482 :  55 - 0x37
      12'h5CB: dout <= 8'b00111010; // 1483 :  58 - 0x3a
      12'h5CC: dout <= 8'b00111101; // 1484 :  61 - 0x3d
      12'h5CD: dout <= 8'b00111110; // 1485 :  62 - 0x3e
      12'h5CE: dout <= 8'b00111111; // 1486 :  63 - 0x3f
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      12'h5D1: dout <= 8'b00000101; // 1489 :   5 - 0x5
      12'h5D2: dout <= 8'b00011001; // 1490 :  25 - 0x19
      12'h5D3: dout <= 8'b00110011; // 1491 :  51 - 0x33
      12'h5D4: dout <= 8'b01100011; // 1492 :  99 - 0x63
      12'h5D5: dout <= 8'b11000111; // 1493 : 199 - 0xc7
      12'h5D6: dout <= 8'b11000111; // 1494 : 199 - 0xc7
      12'h5D7: dout <= 8'b11000100; // 1495 : 196 - 0xc4
      12'h5D8: dout <= 8'b10000000; // 1496 : 128 - 0x80 -- Sprite 0xbb
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b00000011; // 1501 :   3 - 0x3
      12'h5DE: dout <= 8'b00000011; // 1502 :   3 - 0x3
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      12'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      12'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      12'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout <= 8'b00000000; // 1508 :   0 - 0x0
      12'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      12'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b00001111; // 1514 :  15 - 0xf
      12'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout <= 8'b10000000; // 1516 : 128 - 0x80
      12'h5ED: dout <= 8'b01100011; // 1517 :  99 - 0x63
      12'h5EE: dout <= 8'b00011110; // 1518 :  30 - 0x1e
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000001; // 1520 :   1 - 0x1 -- Sprite 0xbe
      12'h5F1: dout <= 8'b00000011; // 1521 :   3 - 0x3
      12'h5F2: dout <= 8'b00011001; // 1522 :  25 - 0x19
      12'h5F3: dout <= 8'b00111100; // 1523 :  60 - 0x3c
      12'h5F4: dout <= 8'b00011001; // 1524 :  25 - 0x19
      12'h5F5: dout <= 8'b00100011; // 1525 :  35 - 0x23
      12'h5F6: dout <= 8'b01010001; // 1526 :  81 - 0x51
      12'h5F7: dout <= 8'b00100000; // 1527 :  32 - 0x20
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout <= 8'b00111111; // 1537 :  63 - 0x3f
      12'h602: dout <= 8'b00011111; // 1538 :  31 - 0x1f
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000001; // 1540 :   1 - 0x1
      12'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout <= 8'b00000001; // 1542 :   1 - 0x1
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00010001; // 1544 :  17 - 0x11 -- Sprite 0xc1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000001; // 1546 :   1 - 0x1
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000001; // 1548 :   1 - 0x1
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00011111; // 1550 :  31 - 0x1f
      12'h60F: dout <= 8'b00111111; // 1551 :  63 - 0x3f
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout <= 8'b11111100; // 1553 : 252 - 0xfc
      12'h612: dout <= 8'b11111000; // 1554 : 248 - 0xf8
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b10000000; // 1556 : 128 - 0x80
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b10000000; // 1558 : 128 - 0x80
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b10001000; // 1560 : 136 - 0x88 -- Sprite 0xc3
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b10000000; // 1562 : 128 - 0x80
      12'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout <= 8'b10000000; // 1564 : 128 - 0x80
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b11111000; // 1566 : 248 - 0xf8
      12'h61F: dout <= 8'b11111100; // 1567 : 252 - 0xfc
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout <= 8'b00111111; // 1573 :  63 - 0x3f
      12'h626: dout <= 8'b00011111; // 1574 :  31 - 0x1f
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b00000001; // 1576 :   1 - 0x1 -- Sprite 0xc5
      12'h629: dout <= 8'b00000001; // 1577 :   1 - 0x1
      12'h62A: dout <= 8'b01000001; // 1578 :  65 - 0x41
      12'h62B: dout <= 8'b00000001; // 1579 :   1 - 0x1
      12'h62C: dout <= 8'b00000001; // 1580 :   1 - 0x1
      12'h62D: dout <= 8'b00000000; // 1581 :   0 - 0x0
      12'h62E: dout <= 8'b00011111; // 1582 :  31 - 0x1f
      12'h62F: dout <= 8'b00111111; // 1583 :  63 - 0x3f
      12'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      12'h631: dout <= 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout <= 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout <= 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout <= 8'b11111100; // 1589 : 252 - 0xfc
      12'h636: dout <= 8'b11111000; // 1590 : 248 - 0xf8
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b10000000; // 1592 : 128 - 0x80 -- Sprite 0xc7
      12'h639: dout <= 8'b10000000; // 1593 : 128 - 0x80
      12'h63A: dout <= 8'b10000010; // 1594 : 130 - 0x82
      12'h63B: dout <= 8'b10000000; // 1595 : 128 - 0x80
      12'h63C: dout <= 8'b10000000; // 1596 : 128 - 0x80
      12'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout <= 8'b11111000; // 1598 : 248 - 0xf8
      12'h63F: dout <= 8'b11111100; // 1599 : 252 - 0xfc
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00011110; // 1603 :  30 - 0x1e
      12'h644: dout <= 8'b00111111; // 1604 :  63 - 0x3f
      12'h645: dout <= 8'b00111111; // 1605 :  63 - 0x3f
      12'h646: dout <= 8'b00111111; // 1606 :  63 - 0x3f
      12'h647: dout <= 8'b00111111; // 1607 :  63 - 0x3f
      12'h648: dout <= 8'b00011111; // 1608 :  31 - 0x1f -- Sprite 0xc9
      12'h649: dout <= 8'b00001111; // 1609 :  15 - 0xf
      12'h64A: dout <= 8'b00000111; // 1610 :   7 - 0x7
      12'h64B: dout <= 8'b00000011; // 1611 :   3 - 0x3
      12'h64C: dout <= 8'b00000001; // 1612 :   1 - 0x1
      12'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00111100; // 1619 :  60 - 0x3c
      12'h654: dout <= 8'b01111110; // 1620 : 126 - 0x7e
      12'h655: dout <= 8'b11111110; // 1621 : 254 - 0xfe
      12'h656: dout <= 8'b11111110; // 1622 : 254 - 0xfe
      12'h657: dout <= 8'b11111110; // 1623 : 254 - 0xfe
      12'h658: dout <= 8'b11111100; // 1624 : 252 - 0xfc -- Sprite 0xcb
      12'h659: dout <= 8'b11111000; // 1625 : 248 - 0xf8
      12'h65A: dout <= 8'b11110000; // 1626 : 240 - 0xf0
      12'h65B: dout <= 8'b11100000; // 1627 : 224 - 0xe0
      12'h65C: dout <= 8'b11000000; // 1628 : 192 - 0xc0
      12'h65D: dout <= 8'b10000000; // 1629 : 128 - 0x80
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b11111111; // 1632 : 255 - 0xff -- Sprite 0xcc
      12'h661: dout <= 8'b11111111; // 1633 : 255 - 0xff
      12'h662: dout <= 8'b11111111; // 1634 : 255 - 0xff
      12'h663: dout <= 8'b11111111; // 1635 : 255 - 0xff
      12'h664: dout <= 8'b11111111; // 1636 : 255 - 0xff
      12'h665: dout <= 8'b11111111; // 1637 : 255 - 0xff
      12'h666: dout <= 8'b11111111; // 1638 : 255 - 0xff
      12'h667: dout <= 8'b11111111; // 1639 : 255 - 0xff
      12'h668: dout <= 8'b11111111; // 1640 : 255 - 0xff -- Sprite 0xcd
      12'h669: dout <= 8'b11111111; // 1641 : 255 - 0xff
      12'h66A: dout <= 8'b11111111; // 1642 : 255 - 0xff
      12'h66B: dout <= 8'b11111111; // 1643 : 255 - 0xff
      12'h66C: dout <= 8'b11111111; // 1644 : 255 - 0xff
      12'h66D: dout <= 8'b11111111; // 1645 : 255 - 0xff
      12'h66E: dout <= 8'b11111111; // 1646 : 255 - 0xff
      12'h66F: dout <= 8'b11111111; // 1647 : 255 - 0xff
      12'h670: dout <= 8'b11111111; // 1648 : 255 - 0xff -- Sprite 0xce
      12'h671: dout <= 8'b11111111; // 1649 : 255 - 0xff
      12'h672: dout <= 8'b11111111; // 1650 : 255 - 0xff
      12'h673: dout <= 8'b11111111; // 1651 : 255 - 0xff
      12'h674: dout <= 8'b11111111; // 1652 : 255 - 0xff
      12'h675: dout <= 8'b11111111; // 1653 : 255 - 0xff
      12'h676: dout <= 8'b11111111; // 1654 : 255 - 0xff
      12'h677: dout <= 8'b11111111; // 1655 : 255 - 0xff
      12'h678: dout <= 8'b11111111; // 1656 : 255 - 0xff -- Sprite 0xcf
      12'h679: dout <= 8'b11111111; // 1657 : 255 - 0xff
      12'h67A: dout <= 8'b11111111; // 1658 : 255 - 0xff
      12'h67B: dout <= 8'b11111111; // 1659 : 255 - 0xff
      12'h67C: dout <= 8'b11111111; // 1660 : 255 - 0xff
      12'h67D: dout <= 8'b11111111; // 1661 : 255 - 0xff
      12'h67E: dout <= 8'b11111111; // 1662 : 255 - 0xff
      12'h67F: dout <= 8'b11111111; // 1663 : 255 - 0xff
      12'h680: dout <= 8'b00001000; // 1664 :   8 - 0x8 -- Sprite 0xd0
      12'h681: dout <= 8'b00011001; // 1665 :  25 - 0x19
      12'h682: dout <= 8'b00001001; // 1666 :   9 - 0x9
      12'h683: dout <= 8'b00001001; // 1667 :   9 - 0x9
      12'h684: dout <= 8'b00001001; // 1668 :   9 - 0x9
      12'h685: dout <= 8'b00001001; // 1669 :   9 - 0x9
      12'h686: dout <= 8'b00011100; // 1670 :  28 - 0x1c
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00111000; // 1672 :  56 - 0x38 -- Sprite 0xd1
      12'h689: dout <= 8'b00000101; // 1673 :   5 - 0x5
      12'h68A: dout <= 8'b00000101; // 1674 :   5 - 0x5
      12'h68B: dout <= 8'b00011001; // 1675 :  25 - 0x19
      12'h68C: dout <= 8'b00000101; // 1676 :   5 - 0x5
      12'h68D: dout <= 8'b00000101; // 1677 :   5 - 0x5
      12'h68E: dout <= 8'b00111000; // 1678 :  56 - 0x38
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b00111100; // 1680 :  60 - 0x3c -- Sprite 0xd2
      12'h691: dout <= 8'b00100001; // 1681 :  33 - 0x21
      12'h692: dout <= 8'b00100001; // 1682 :  33 - 0x21
      12'h693: dout <= 8'b00111101; // 1683 :  61 - 0x3d
      12'h694: dout <= 8'b00000101; // 1684 :   5 - 0x5
      12'h695: dout <= 8'b00000101; // 1685 :   5 - 0x5
      12'h696: dout <= 8'b00111000; // 1686 :  56 - 0x38
      12'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout <= 8'b00011000; // 1688 :  24 - 0x18 -- Sprite 0xd3
      12'h699: dout <= 8'b00100101; // 1689 :  37 - 0x25
      12'h69A: dout <= 8'b00100101; // 1690 :  37 - 0x25
      12'h69B: dout <= 8'b00011001; // 1691 :  25 - 0x19
      12'h69C: dout <= 8'b00100101; // 1692 :  37 - 0x25
      12'h69D: dout <= 8'b00100101; // 1693 :  37 - 0x25
      12'h69E: dout <= 8'b00011000; // 1694 :  24 - 0x18
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b11000110; // 1696 : 198 - 0xc6 -- Sprite 0xd4
      12'h6A1: dout <= 8'b00101001; // 1697 :  41 - 0x29
      12'h6A2: dout <= 8'b00101001; // 1698 :  41 - 0x29
      12'h6A3: dout <= 8'b00101001; // 1699 :  41 - 0x29
      12'h6A4: dout <= 8'b00101001; // 1700 :  41 - 0x29
      12'h6A5: dout <= 8'b00101001; // 1701 :  41 - 0x29
      12'h6A6: dout <= 8'b11000110; // 1702 : 198 - 0xc6
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      12'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout <= 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout <= 8'b00111100; // 1716 :  60 - 0x3c
      12'h6B5: dout <= 8'b10110110; // 1717 : 182 - 0xb6
      12'h6B6: dout <= 8'b01111100; // 1718 : 124 - 0x7c
      12'h6B7: dout <= 8'b11111000; // 1719 : 248 - 0xf8
      12'h6B8: dout <= 8'b00000011; // 1720 :   3 - 0x3 -- Sprite 0xd7
      12'h6B9: dout <= 8'b00000011; // 1721 :   3 - 0x3
      12'h6BA: dout <= 8'b00000011; // 1722 :   3 - 0x3
      12'h6BB: dout <= 8'b00000111; // 1723 :   7 - 0x7
      12'h6BC: dout <= 8'b00001100; // 1724 :  12 - 0xc
      12'h6BD: dout <= 8'b00011011; // 1725 :  27 - 0x1b
      12'h6BE: dout <= 8'b01110111; // 1726 : 119 - 0x77
      12'h6BF: dout <= 8'b00000111; // 1727 :   7 - 0x7
      12'h6C0: dout <= 8'b00001111; // 1728 :  15 - 0xf -- Sprite 0xd8
      12'h6C1: dout <= 8'b00001111; // 1729 :  15 - 0xf
      12'h6C2: dout <= 8'b00011111; // 1730 :  31 - 0x1f
      12'h6C3: dout <= 8'b00111111; // 1731 :  63 - 0x3f
      12'h6C4: dout <= 8'b01111111; // 1732 : 127 - 0x7f
      12'h6C5: dout <= 8'b00111111; // 1733 :  63 - 0x3f
      12'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout <= 8'b11100000; // 1736 : 224 - 0xe0 -- Sprite 0xd9
      12'h6C9: dout <= 8'b11110000; // 1737 : 240 - 0xf0
      12'h6CA: dout <= 8'b11110000; // 1738 : 240 - 0xf0
      12'h6CB: dout <= 8'b11110000; // 1739 : 240 - 0xf0
      12'h6CC: dout <= 8'b00011000; // 1740 :  24 - 0x18
      12'h6CD: dout <= 8'b11111100; // 1741 : 252 - 0xfc
      12'h6CE: dout <= 8'b11111100; // 1742 : 252 - 0xfc
      12'h6CF: dout <= 8'b11111100; // 1743 : 252 - 0xfc
      12'h6D0: dout <= 8'b11111000; // 1744 : 248 - 0xf8 -- Sprite 0xda
      12'h6D1: dout <= 8'b11111100; // 1745 : 252 - 0xfc
      12'h6D2: dout <= 8'b11111111; // 1746 : 255 - 0xff
      12'h6D3: dout <= 8'b11111111; // 1747 : 255 - 0xff
      12'h6D4: dout <= 8'b11111110; // 1748 : 254 - 0xfe
      12'h6D5: dout <= 8'b11110000; // 1749 : 240 - 0xf0
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000011; // 1752 :   3 - 0x3 -- Sprite 0xdb
      12'h6D9: dout <= 8'b00000011; // 1753 :   3 - 0x3
      12'h6DA: dout <= 8'b00000011; // 1754 :   3 - 0x3
      12'h6DB: dout <= 8'b00000011; // 1755 :   3 - 0x3
      12'h6DC: dout <= 8'b00000001; // 1756 :   1 - 0x1
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000111; // 1758 :   7 - 0x7
      12'h6DF: dout <= 8'b00011111; // 1759 :  31 - 0x1f
      12'h6E0: dout <= 8'b11111111; // 1760 : 255 - 0xff -- Sprite 0xdc
      12'h6E1: dout <= 8'b11111111; // 1761 : 255 - 0xff
      12'h6E2: dout <= 8'b01111111; // 1762 : 127 - 0x7f
      12'h6E3: dout <= 8'b00111111; // 1763 :  63 - 0x3f
      12'h6E4: dout <= 8'b00001111; // 1764 :  15 - 0xf
      12'h6E5: dout <= 8'b00000011; // 1765 :   3 - 0x3
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b11100000; // 1768 : 224 - 0xe0 -- Sprite 0xdd
      12'h6E9: dout <= 8'b11110000; // 1769 : 240 - 0xf0
      12'h6EA: dout <= 8'b11110000; // 1770 : 240 - 0xf0
      12'h6EB: dout <= 8'b11100000; // 1771 : 224 - 0xe0
      12'h6EC: dout <= 8'b11111110; // 1772 : 254 - 0xfe
      12'h6ED: dout <= 8'b00111100; // 1773 :  60 - 0x3c
      12'h6EE: dout <= 8'b11110000; // 1774 : 240 - 0xf0
      12'h6EF: dout <= 8'b11111100; // 1775 : 252 - 0xfc
      12'h6F0: dout <= 8'b11111100; // 1776 : 252 - 0xfc -- Sprite 0xde
      12'h6F1: dout <= 8'b11111000; // 1777 : 248 - 0xf8
      12'h6F2: dout <= 8'b11111000; // 1778 : 248 - 0xf8
      12'h6F3: dout <= 8'b11111000; // 1779 : 248 - 0xf8
      12'h6F4: dout <= 8'b11111000; // 1780 : 248 - 0xf8
      12'h6F5: dout <= 8'b11111000; // 1781 : 248 - 0xf8
      12'h6F6: dout <= 8'b11111000; // 1782 : 248 - 0xf8
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b11111111; // 1784 : 255 - 0xff -- Sprite 0xdf
      12'h6F9: dout <= 8'b11111111; // 1785 : 255 - 0xff
      12'h6FA: dout <= 8'b11111111; // 1786 : 255 - 0xff
      12'h6FB: dout <= 8'b11111111; // 1787 : 255 - 0xff
      12'h6FC: dout <= 8'b11111111; // 1788 : 255 - 0xff
      12'h6FD: dout <= 8'b11111111; // 1789 : 255 - 0xff
      12'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      12'h6FF: dout <= 8'b11111111; // 1791 : 255 - 0xff
      12'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0xe0
      12'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      12'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      12'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      12'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      12'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      12'h70A: dout <= 8'b11111111; // 1802 : 255 - 0xff
      12'h70B: dout <= 8'b11111111; // 1803 : 255 - 0xff
      12'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      12'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      12'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      12'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      12'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0xe2
      12'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      12'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      12'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      12'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      12'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      12'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      12'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      12'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      12'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      12'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      12'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      12'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      12'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0xe4
      12'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      12'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      12'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      12'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      12'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      12'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      12'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      12'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      12'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      12'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      12'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      12'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      12'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0xe6
      12'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      12'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      12'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      12'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      12'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout <= 8'b11111111; // 1850 : 255 - 0xff
      12'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      12'h73C: dout <= 8'b11111111; // 1852 : 255 - 0xff
      12'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      12'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      12'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      12'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      12'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      12'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      12'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      12'h748: dout <= 8'b11111111; // 1864 : 255 - 0xff -- Sprite 0xe9
      12'h749: dout <= 8'b11111111; // 1865 : 255 - 0xff
      12'h74A: dout <= 8'b11111111; // 1866 : 255 - 0xff
      12'h74B: dout <= 8'b11111111; // 1867 : 255 - 0xff
      12'h74C: dout <= 8'b11111111; // 1868 : 255 - 0xff
      12'h74D: dout <= 8'b11111111; // 1869 : 255 - 0xff
      12'h74E: dout <= 8'b11111111; // 1870 : 255 - 0xff
      12'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      12'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      12'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      12'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      12'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      12'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff -- Sprite 0xeb
      12'h759: dout <= 8'b11111111; // 1881 : 255 - 0xff
      12'h75A: dout <= 8'b11111111; // 1882 : 255 - 0xff
      12'h75B: dout <= 8'b11111111; // 1883 : 255 - 0xff
      12'h75C: dout <= 8'b11111111; // 1884 : 255 - 0xff
      12'h75D: dout <= 8'b11111111; // 1885 : 255 - 0xff
      12'h75E: dout <= 8'b11111111; // 1886 : 255 - 0xff
      12'h75F: dout <= 8'b11111111; // 1887 : 255 - 0xff
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b00000001; // 1889 :   1 - 0x1
      12'h762: dout <= 8'b00000011; // 1890 :   3 - 0x3
      12'h763: dout <= 8'b00110011; // 1891 :  51 - 0x33
      12'h764: dout <= 8'b00011001; // 1892 :  25 - 0x19
      12'h765: dout <= 8'b00001111; // 1893 :  15 - 0xf
      12'h766: dout <= 8'b00111111; // 1894 :  63 - 0x3f
      12'h767: dout <= 8'b00011111; // 1895 :  31 - 0x1f
      12'h768: dout <= 8'b00101011; // 1896 :  43 - 0x2b -- Sprite 0xed
      12'h769: dout <= 8'b00000111; // 1897 :   7 - 0x7
      12'h76A: dout <= 8'b00000101; // 1898 :   5 - 0x5
      12'h76B: dout <= 8'b00001101; // 1899 :  13 - 0xd
      12'h76C: dout <= 8'b00001011; // 1900 :  11 - 0xb
      12'h76D: dout <= 8'b00011011; // 1901 :  27 - 0x1b
      12'h76E: dout <= 8'b00011011; // 1902 :  27 - 0x1b
      12'h76F: dout <= 8'b00111011; // 1903 :  59 - 0x3b
      12'h770: dout <= 8'b00001001; // 1904 :   9 - 0x9 -- Sprite 0xee
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000111; // 1906 :   7 - 0x7
      12'h773: dout <= 8'b00000111; // 1907 :   7 - 0x7
      12'h774: dout <= 8'b00001111; // 1908 :  15 - 0xf
      12'h775: dout <= 8'b00001101; // 1909 :  13 - 0xd
      12'h776: dout <= 8'b00000001; // 1910 :   1 - 0x1
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b11111000; // 1912 : 248 - 0xf8 -- Sprite 0xef
      12'h779: dout <= 8'b11111100; // 1913 : 252 - 0xfc
      12'h77A: dout <= 8'b11111000; // 1914 : 248 - 0xf8
      12'h77B: dout <= 8'b11101100; // 1915 : 236 - 0xec
      12'h77C: dout <= 8'b11111000; // 1916 : 248 - 0xf8
      12'h77D: dout <= 8'b11110000; // 1917 : 240 - 0xf0
      12'h77E: dout <= 8'b11000000; // 1918 : 192 - 0xc0
      12'h77F: dout <= 8'b11000000; // 1919 : 192 - 0xc0
      12'h780: dout <= 8'b11110000; // 1920 : 240 - 0xf0 -- Sprite 0xf0
      12'h781: dout <= 8'b11111000; // 1921 : 248 - 0xf8
      12'h782: dout <= 8'b11111000; // 1922 : 248 - 0xf8
      12'h783: dout <= 8'b11101000; // 1923 : 232 - 0xe8
      12'h784: dout <= 8'b11001100; // 1924 : 204 - 0xcc
      12'h785: dout <= 8'b11100110; // 1925 : 230 - 0xe6
      12'h786: dout <= 8'b11111011; // 1926 : 251 - 0xfb
      12'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      12'h789: dout <= 8'b11111110; // 1929 : 254 - 0xfe
      12'h78A: dout <= 8'b11111110; // 1930 : 254 - 0xfe
      12'h78B: dout <= 8'b11111110; // 1931 : 254 - 0xfe
      12'h78C: dout <= 8'b11111110; // 1932 : 254 - 0xfe
      12'h78D: dout <= 8'b10001111; // 1933 : 143 - 0x8f
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000001; // 1936 :   1 - 0x1 -- Sprite 0xf2
      12'h791: dout <= 8'b00001111; // 1937 :  15 - 0xf
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000100; // 1940 :   4 - 0x4
      12'h795: dout <= 8'b00011110; // 1941 :  30 - 0x1e
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000011; // 1943 :   3 - 0x3
      12'h798: dout <= 8'b00000111; // 1944 :   7 - 0x7 -- Sprite 0xf3
      12'h799: dout <= 8'b00001111; // 1945 :  15 - 0xf
      12'h79A: dout <= 8'b00011111; // 1946 :  31 - 0x1f
      12'h79B: dout <= 8'b00001111; // 1947 :  15 - 0xf
      12'h79C: dout <= 8'b00000111; // 1948 :   7 - 0x7
      12'h79D: dout <= 8'b00001111; // 1949 :  15 - 0xf
      12'h79E: dout <= 8'b00001111; // 1950 :  15 - 0xf
      12'h79F: dout <= 8'b00000011; // 1951 :   3 - 0x3
      12'h7A0: dout <= 8'b11100000; // 1952 : 224 - 0xe0 -- Sprite 0xf4
      12'h7A1: dout <= 8'b11110000; // 1953 : 240 - 0xf0
      12'h7A2: dout <= 8'b11110000; // 1954 : 240 - 0xf0
      12'h7A3: dout <= 8'b01001000; // 1955 :  72 - 0x48
      12'h7A4: dout <= 8'b11001000; // 1956 : 200 - 0xc8
      12'h7A5: dout <= 8'b10011100; // 1957 : 156 - 0x9c
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b11110000; // 1959 : 240 - 0xf0
      12'h7A8: dout <= 8'b11111000; // 1960 : 248 - 0xf8 -- Sprite 0xf5
      12'h7A9: dout <= 8'b11111100; // 1961 : 252 - 0xfc
      12'h7AA: dout <= 8'b11111100; // 1962 : 252 - 0xfc
      12'h7AB: dout <= 8'b11111000; // 1963 : 248 - 0xf8
      12'h7AC: dout <= 8'b11111000; // 1964 : 248 - 0xf8
      12'h7AD: dout <= 8'b01111000; // 1965 : 120 - 0x78
      12'h7AE: dout <= 8'b01110000; // 1966 : 112 - 0x70
      12'h7AF: dout <= 8'b01100000; // 1967 :  96 - 0x60
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b01111100; // 1970 : 124 - 0x7c
      12'h7B3: dout <= 8'b10001010; // 1971 : 138 - 0x8a
      12'h7B4: dout <= 8'b11111110; // 1972 : 254 - 0xfe
      12'h7B5: dout <= 8'b11111110; // 1973 : 254 - 0xfe
      12'h7B6: dout <= 8'b11111110; // 1974 : 254 - 0xfe
      12'h7B7: dout <= 8'b11111110; // 1975 : 254 - 0xfe
      12'h7B8: dout <= 8'b11111110; // 1976 : 254 - 0xfe -- Sprite 0xf7
      12'h7B9: dout <= 8'b01111100; // 1977 : 124 - 0x7c
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000111; // 1984 :   7 - 0x7 -- Sprite 0xf8
      12'h7C1: dout <= 8'b00001011; // 1985 :  11 - 0xb
      12'h7C2: dout <= 8'b00001111; // 1986 :  15 - 0xf
      12'h7C3: dout <= 8'b00001011; // 1987 :  11 - 0xb
      12'h7C4: dout <= 8'b00001011; // 1988 :  11 - 0xb
      12'h7C5: dout <= 8'b00001011; // 1989 :  11 - 0xb
      12'h7C6: dout <= 8'b00001011; // 1990 :  11 - 0xb
      12'h7C7: dout <= 8'b00000111; // 1991 :   7 - 0x7
      12'h7C8: dout <= 8'b11000000; // 1992 : 192 - 0xc0 -- Sprite 0xf9
      12'h7C9: dout <= 8'b11100000; // 1993 : 224 - 0xe0
      12'h7CA: dout <= 8'b11100000; // 1994 : 224 - 0xe0
      12'h7CB: dout <= 8'b11100000; // 1995 : 224 - 0xe0
      12'h7CC: dout <= 8'b11100000; // 1996 : 224 - 0xe0
      12'h7CD: dout <= 8'b11100000; // 1997 : 224 - 0xe0
      12'h7CE: dout <= 8'b11100000; // 1998 : 224 - 0xe0
      12'h7CF: dout <= 8'b11000000; // 1999 : 192 - 0xc0
      12'h7D0: dout <= 8'b00000011; // 2000 :   3 - 0x3 -- Sprite 0xfa
      12'h7D1: dout <= 8'b00000111; // 2001 :   7 - 0x7
      12'h7D2: dout <= 8'b00000111; // 2002 :   7 - 0x7
      12'h7D3: dout <= 8'b00000111; // 2003 :   7 - 0x7
      12'h7D4: dout <= 8'b00000111; // 2004 :   7 - 0x7
      12'h7D5: dout <= 8'b00000111; // 2005 :   7 - 0x7
      12'h7D6: dout <= 8'b00000111; // 2006 :   7 - 0x7
      12'h7D7: dout <= 8'b00000011; // 2007 :   3 - 0x3
      12'h7D8: dout <= 8'b11100000; // 2008 : 224 - 0xe0 -- Sprite 0xfb
      12'h7D9: dout <= 8'b11010000; // 2009 : 208 - 0xd0
      12'h7DA: dout <= 8'b11010000; // 2010 : 208 - 0xd0
      12'h7DB: dout <= 8'b11010000; // 2011 : 208 - 0xd0
      12'h7DC: dout <= 8'b11010000; // 2012 : 208 - 0xd0
      12'h7DD: dout <= 8'b11110000; // 2013 : 240 - 0xf0
      12'h7DE: dout <= 8'b11010000; // 2014 : 208 - 0xd0
      12'h7DF: dout <= 8'b11100000; // 2015 : 224 - 0xe0
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout <= 8'b00000001; // 2017 :   1 - 0x1
      12'h7E2: dout <= 8'b00010011; // 2018 :  19 - 0x13
      12'h7E3: dout <= 8'b00110111; // 2019 :  55 - 0x37
      12'h7E4: dout <= 8'b00111011; // 2020 :  59 - 0x3b
      12'h7E5: dout <= 8'b01110100; // 2021 : 116 - 0x74
      12'h7E6: dout <= 8'b01111010; // 2022 : 122 - 0x7a
      12'h7E7: dout <= 8'b00111110; // 2023 :  62 - 0x3e
      12'h7E8: dout <= 8'b11011000; // 2024 : 216 - 0xd8 -- Sprite 0xfd
      12'h7E9: dout <= 8'b10011000; // 2025 : 152 - 0x98
      12'h7EA: dout <= 8'b10101000; // 2026 : 168 - 0xa8
      12'h7EB: dout <= 8'b11011000; // 2027 : 216 - 0xd8
      12'h7EC: dout <= 8'b11011010; // 2028 : 218 - 0xda
      12'h7ED: dout <= 8'b01110100; // 2029 : 116 - 0x74
      12'h7EE: dout <= 8'b00101000; // 2030 :  40 - 0x28
      12'h7EF: dout <= 8'b11001000; // 2031 : 200 - 0xc8
      12'h7F0: dout <= 8'b00001000; // 2032 :   8 - 0x8 -- Sprite 0xfe
      12'h7F1: dout <= 8'b01011001; // 2033 :  89 - 0x59
      12'h7F2: dout <= 8'b00110000; // 2034 :  48 - 0x30
      12'h7F3: dout <= 8'b01110001; // 2035 : 113 - 0x71
      12'h7F4: dout <= 8'b01111001; // 2036 : 121 - 0x79
      12'h7F5: dout <= 8'b00101011; // 2037 :  43 - 0x2b
      12'h7F6: dout <= 8'b00110110; // 2038 :  54 - 0x36
      12'h7F7: dout <= 8'b00010110; // 2039 :  22 - 0x16
      12'h7F8: dout <= 8'b11000110; // 2040 : 198 - 0xc6 -- Sprite 0xff
      12'h7F9: dout <= 8'b11000100; // 2041 : 196 - 0xc4
      12'h7FA: dout <= 8'b11001100; // 2042 : 204 - 0xcc
      12'h7FB: dout <= 8'b11001100; // 2043 : 204 - 0xcc
      12'h7FC: dout <= 8'b10111000; // 2044 : 184 - 0xb8
      12'h7FD: dout <= 8'b01111100; // 2045 : 124 - 0x7c
      12'h7FE: dout <= 8'b11101100; // 2046 : 236 - 0xec
      12'h7FF: dout <= 8'b11001000; // 2047 : 200 - 0xc8
          // Background pattern Table
      12'h800: dout <= 8'b00111000; // 2048 :  56 - 0x38 -- Background 0x0
      12'h801: dout <= 8'b01001100; // 2049 :  76 - 0x4c
      12'h802: dout <= 8'b11000110; // 2050 : 198 - 0xc6
      12'h803: dout <= 8'b11000110; // 2051 : 198 - 0xc6
      12'h804: dout <= 8'b11000110; // 2052 : 198 - 0xc6
      12'h805: dout <= 8'b01100100; // 2053 : 100 - 0x64
      12'h806: dout <= 8'b00111000; // 2054 :  56 - 0x38
      12'h807: dout <= 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout <= 8'b00011000; // 2056 :  24 - 0x18 -- Background 0x1
      12'h809: dout <= 8'b00111000; // 2057 :  56 - 0x38
      12'h80A: dout <= 8'b00011000; // 2058 :  24 - 0x18
      12'h80B: dout <= 8'b00011000; // 2059 :  24 - 0x18
      12'h80C: dout <= 8'b00011000; // 2060 :  24 - 0x18
      12'h80D: dout <= 8'b00011000; // 2061 :  24 - 0x18
      12'h80E: dout <= 8'b01111110; // 2062 : 126 - 0x7e
      12'h80F: dout <= 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout <= 8'b01111100; // 2064 : 124 - 0x7c -- Background 0x2
      12'h811: dout <= 8'b11000110; // 2065 : 198 - 0xc6
      12'h812: dout <= 8'b00001110; // 2066 :  14 - 0xe
      12'h813: dout <= 8'b00111100; // 2067 :  60 - 0x3c
      12'h814: dout <= 8'b01111000; // 2068 : 120 - 0x78
      12'h815: dout <= 8'b11100000; // 2069 : 224 - 0xe0
      12'h816: dout <= 8'b11111110; // 2070 : 254 - 0xfe
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b01111110; // 2072 : 126 - 0x7e -- Background 0x3
      12'h819: dout <= 8'b00001100; // 2073 :  12 - 0xc
      12'h81A: dout <= 8'b00011000; // 2074 :  24 - 0x18
      12'h81B: dout <= 8'b00111100; // 2075 :  60 - 0x3c
      12'h81C: dout <= 8'b00000110; // 2076 :   6 - 0x6
      12'h81D: dout <= 8'b11000110; // 2077 : 198 - 0xc6
      12'h81E: dout <= 8'b01111100; // 2078 : 124 - 0x7c
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b00011100; // 2080 :  28 - 0x1c -- Background 0x4
      12'h821: dout <= 8'b00111100; // 2081 :  60 - 0x3c
      12'h822: dout <= 8'b01101100; // 2082 : 108 - 0x6c
      12'h823: dout <= 8'b11001100; // 2083 : 204 - 0xcc
      12'h824: dout <= 8'b11111110; // 2084 : 254 - 0xfe
      12'h825: dout <= 8'b00001100; // 2085 :  12 - 0xc
      12'h826: dout <= 8'b00001100; // 2086 :  12 - 0xc
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b11111100; // 2088 : 252 - 0xfc -- Background 0x5
      12'h829: dout <= 8'b11000000; // 2089 : 192 - 0xc0
      12'h82A: dout <= 8'b11111100; // 2090 : 252 - 0xfc
      12'h82B: dout <= 8'b00000110; // 2091 :   6 - 0x6
      12'h82C: dout <= 8'b00000110; // 2092 :   6 - 0x6
      12'h82D: dout <= 8'b11000110; // 2093 : 198 - 0xc6
      12'h82E: dout <= 8'b01111100; // 2094 : 124 - 0x7c
      12'h82F: dout <= 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout <= 8'b00111100; // 2096 :  60 - 0x3c -- Background 0x6
      12'h831: dout <= 8'b01100000; // 2097 :  96 - 0x60
      12'h832: dout <= 8'b11000000; // 2098 : 192 - 0xc0
      12'h833: dout <= 8'b11111100; // 2099 : 252 - 0xfc
      12'h834: dout <= 8'b11000110; // 2100 : 198 - 0xc6
      12'h835: dout <= 8'b11000110; // 2101 : 198 - 0xc6
      12'h836: dout <= 8'b01111100; // 2102 : 124 - 0x7c
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b11111110; // 2104 : 254 - 0xfe -- Background 0x7
      12'h839: dout <= 8'b11000110; // 2105 : 198 - 0xc6
      12'h83A: dout <= 8'b00001100; // 2106 :  12 - 0xc
      12'h83B: dout <= 8'b00011000; // 2107 :  24 - 0x18
      12'h83C: dout <= 8'b00110000; // 2108 :  48 - 0x30
      12'h83D: dout <= 8'b00110000; // 2109 :  48 - 0x30
      12'h83E: dout <= 8'b00110000; // 2110 :  48 - 0x30
      12'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout <= 8'b01111000; // 2112 : 120 - 0x78 -- Background 0x8
      12'h841: dout <= 8'b11000100; // 2113 : 196 - 0xc4
      12'h842: dout <= 8'b11100100; // 2114 : 228 - 0xe4
      12'h843: dout <= 8'b01111000; // 2115 : 120 - 0x78
      12'h844: dout <= 8'b10000110; // 2116 : 134 - 0x86
      12'h845: dout <= 8'b10000110; // 2117 : 134 - 0x86
      12'h846: dout <= 8'b01111100; // 2118 : 124 - 0x7c
      12'h847: dout <= 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout <= 8'b01111100; // 2120 : 124 - 0x7c -- Background 0x9
      12'h849: dout <= 8'b11000110; // 2121 : 198 - 0xc6
      12'h84A: dout <= 8'b11000110; // 2122 : 198 - 0xc6
      12'h84B: dout <= 8'b01111110; // 2123 : 126 - 0x7e
      12'h84C: dout <= 8'b00000110; // 2124 :   6 - 0x6
      12'h84D: dout <= 8'b00001100; // 2125 :  12 - 0xc
      12'h84E: dout <= 8'b01111000; // 2126 : 120 - 0x78
      12'h84F: dout <= 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout <= 8'b00111000; // 2128 :  56 - 0x38 -- Background 0xa
      12'h851: dout <= 8'b01101100; // 2129 : 108 - 0x6c
      12'h852: dout <= 8'b11000110; // 2130 : 198 - 0xc6
      12'h853: dout <= 8'b11000110; // 2131 : 198 - 0xc6
      12'h854: dout <= 8'b11111110; // 2132 : 254 - 0xfe
      12'h855: dout <= 8'b11000110; // 2133 : 198 - 0xc6
      12'h856: dout <= 8'b11000110; // 2134 : 198 - 0xc6
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b11111100; // 2136 : 252 - 0xfc -- Background 0xb
      12'h859: dout <= 8'b11000110; // 2137 : 198 - 0xc6
      12'h85A: dout <= 8'b11000110; // 2138 : 198 - 0xc6
      12'h85B: dout <= 8'b11111100; // 2139 : 252 - 0xfc
      12'h85C: dout <= 8'b11000110; // 2140 : 198 - 0xc6
      12'h85D: dout <= 8'b11000110; // 2141 : 198 - 0xc6
      12'h85E: dout <= 8'b11111100; // 2142 : 252 - 0xfc
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b00111100; // 2144 :  60 - 0x3c -- Background 0xc
      12'h861: dout <= 8'b01100110; // 2145 : 102 - 0x66
      12'h862: dout <= 8'b11000000; // 2146 : 192 - 0xc0
      12'h863: dout <= 8'b11000000; // 2147 : 192 - 0xc0
      12'h864: dout <= 8'b11000000; // 2148 : 192 - 0xc0
      12'h865: dout <= 8'b01100110; // 2149 : 102 - 0x66
      12'h866: dout <= 8'b00111100; // 2150 :  60 - 0x3c
      12'h867: dout <= 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout <= 8'b11111000; // 2152 : 248 - 0xf8 -- Background 0xd
      12'h869: dout <= 8'b11001100; // 2153 : 204 - 0xcc
      12'h86A: dout <= 8'b11000110; // 2154 : 198 - 0xc6
      12'h86B: dout <= 8'b11000110; // 2155 : 198 - 0xc6
      12'h86C: dout <= 8'b11000110; // 2156 : 198 - 0xc6
      12'h86D: dout <= 8'b11001100; // 2157 : 204 - 0xcc
      12'h86E: dout <= 8'b11111000; // 2158 : 248 - 0xf8
      12'h86F: dout <= 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout <= 8'b11111110; // 2160 : 254 - 0xfe -- Background 0xe
      12'h871: dout <= 8'b11000000; // 2161 : 192 - 0xc0
      12'h872: dout <= 8'b11000000; // 2162 : 192 - 0xc0
      12'h873: dout <= 8'b11111100; // 2163 : 252 - 0xfc
      12'h874: dout <= 8'b11000000; // 2164 : 192 - 0xc0
      12'h875: dout <= 8'b11000000; // 2165 : 192 - 0xc0
      12'h876: dout <= 8'b11111110; // 2166 : 254 - 0xfe
      12'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout <= 8'b11111110; // 2168 : 254 - 0xfe -- Background 0xf
      12'h879: dout <= 8'b11000000; // 2169 : 192 - 0xc0
      12'h87A: dout <= 8'b11000000; // 2170 : 192 - 0xc0
      12'h87B: dout <= 8'b11111100; // 2171 : 252 - 0xfc
      12'h87C: dout <= 8'b11000000; // 2172 : 192 - 0xc0
      12'h87D: dout <= 8'b11000000; // 2173 : 192 - 0xc0
      12'h87E: dout <= 8'b11000000; // 2174 : 192 - 0xc0
      12'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout <= 8'b00111110; // 2176 :  62 - 0x3e -- Background 0x10
      12'h881: dout <= 8'b01100000; // 2177 :  96 - 0x60
      12'h882: dout <= 8'b11000000; // 2178 : 192 - 0xc0
      12'h883: dout <= 8'b11011110; // 2179 : 222 - 0xde
      12'h884: dout <= 8'b11000110; // 2180 : 198 - 0xc6
      12'h885: dout <= 8'b01100110; // 2181 : 102 - 0x66
      12'h886: dout <= 8'b01111110; // 2182 : 126 - 0x7e
      12'h887: dout <= 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout <= 8'b11000110; // 2184 : 198 - 0xc6 -- Background 0x11
      12'h889: dout <= 8'b11000110; // 2185 : 198 - 0xc6
      12'h88A: dout <= 8'b11000110; // 2186 : 198 - 0xc6
      12'h88B: dout <= 8'b11111110; // 2187 : 254 - 0xfe
      12'h88C: dout <= 8'b11000110; // 2188 : 198 - 0xc6
      12'h88D: dout <= 8'b11000110; // 2189 : 198 - 0xc6
      12'h88E: dout <= 8'b11000110; // 2190 : 198 - 0xc6
      12'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout <= 8'b01111110; // 2192 : 126 - 0x7e -- Background 0x12
      12'h891: dout <= 8'b00011000; // 2193 :  24 - 0x18
      12'h892: dout <= 8'b00011000; // 2194 :  24 - 0x18
      12'h893: dout <= 8'b00011000; // 2195 :  24 - 0x18
      12'h894: dout <= 8'b00011000; // 2196 :  24 - 0x18
      12'h895: dout <= 8'b00011000; // 2197 :  24 - 0x18
      12'h896: dout <= 8'b01111110; // 2198 : 126 - 0x7e
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00011110; // 2200 :  30 - 0x1e -- Background 0x13
      12'h899: dout <= 8'b00000110; // 2201 :   6 - 0x6
      12'h89A: dout <= 8'b00000110; // 2202 :   6 - 0x6
      12'h89B: dout <= 8'b00000110; // 2203 :   6 - 0x6
      12'h89C: dout <= 8'b11000110; // 2204 : 198 - 0xc6
      12'h89D: dout <= 8'b11000110; // 2205 : 198 - 0xc6
      12'h89E: dout <= 8'b01111100; // 2206 : 124 - 0x7c
      12'h89F: dout <= 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout <= 8'b11000110; // 2208 : 198 - 0xc6 -- Background 0x14
      12'h8A1: dout <= 8'b11001100; // 2209 : 204 - 0xcc
      12'h8A2: dout <= 8'b11011000; // 2210 : 216 - 0xd8
      12'h8A3: dout <= 8'b11110000; // 2211 : 240 - 0xf0
      12'h8A4: dout <= 8'b11111000; // 2212 : 248 - 0xf8
      12'h8A5: dout <= 8'b11011100; // 2213 : 220 - 0xdc
      12'h8A6: dout <= 8'b11001110; // 2214 : 206 - 0xce
      12'h8A7: dout <= 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout <= 8'b01100000; // 2216 :  96 - 0x60 -- Background 0x15
      12'h8A9: dout <= 8'b01100000; // 2217 :  96 - 0x60
      12'h8AA: dout <= 8'b01100000; // 2218 :  96 - 0x60
      12'h8AB: dout <= 8'b01100000; // 2219 :  96 - 0x60
      12'h8AC: dout <= 8'b01100000; // 2220 :  96 - 0x60
      12'h8AD: dout <= 8'b01100000; // 2221 :  96 - 0x60
      12'h8AE: dout <= 8'b01111110; // 2222 : 126 - 0x7e
      12'h8AF: dout <= 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout <= 8'b11000110; // 2224 : 198 - 0xc6 -- Background 0x16
      12'h8B1: dout <= 8'b11101110; // 2225 : 238 - 0xee
      12'h8B2: dout <= 8'b11111110; // 2226 : 254 - 0xfe
      12'h8B3: dout <= 8'b11111110; // 2227 : 254 - 0xfe
      12'h8B4: dout <= 8'b11010110; // 2228 : 214 - 0xd6
      12'h8B5: dout <= 8'b11000110; // 2229 : 198 - 0xc6
      12'h8B6: dout <= 8'b11000110; // 2230 : 198 - 0xc6
      12'h8B7: dout <= 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout <= 8'b11000110; // 2232 : 198 - 0xc6 -- Background 0x17
      12'h8B9: dout <= 8'b11100110; // 2233 : 230 - 0xe6
      12'h8BA: dout <= 8'b11110110; // 2234 : 246 - 0xf6
      12'h8BB: dout <= 8'b11111110; // 2235 : 254 - 0xfe
      12'h8BC: dout <= 8'b11011110; // 2236 : 222 - 0xde
      12'h8BD: dout <= 8'b11001110; // 2237 : 206 - 0xce
      12'h8BE: dout <= 8'b11000110; // 2238 : 198 - 0xc6
      12'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout <= 8'b01111100; // 2240 : 124 - 0x7c -- Background 0x18
      12'h8C1: dout <= 8'b11000110; // 2241 : 198 - 0xc6
      12'h8C2: dout <= 8'b11000110; // 2242 : 198 - 0xc6
      12'h8C3: dout <= 8'b11000110; // 2243 : 198 - 0xc6
      12'h8C4: dout <= 8'b11000110; // 2244 : 198 - 0xc6
      12'h8C5: dout <= 8'b11000110; // 2245 : 198 - 0xc6
      12'h8C6: dout <= 8'b01111100; // 2246 : 124 - 0x7c
      12'h8C7: dout <= 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout <= 8'b11111100; // 2248 : 252 - 0xfc -- Background 0x19
      12'h8C9: dout <= 8'b11000110; // 2249 : 198 - 0xc6
      12'h8CA: dout <= 8'b11000110; // 2250 : 198 - 0xc6
      12'h8CB: dout <= 8'b11000110; // 2251 : 198 - 0xc6
      12'h8CC: dout <= 8'b11111100; // 2252 : 252 - 0xfc
      12'h8CD: dout <= 8'b11000000; // 2253 : 192 - 0xc0
      12'h8CE: dout <= 8'b11000000; // 2254 : 192 - 0xc0
      12'h8CF: dout <= 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout <= 8'b01111100; // 2256 : 124 - 0x7c -- Background 0x1a
      12'h8D1: dout <= 8'b11000110; // 2257 : 198 - 0xc6
      12'h8D2: dout <= 8'b11000110; // 2258 : 198 - 0xc6
      12'h8D3: dout <= 8'b11000110; // 2259 : 198 - 0xc6
      12'h8D4: dout <= 8'b11011110; // 2260 : 222 - 0xde
      12'h8D5: dout <= 8'b11001100; // 2261 : 204 - 0xcc
      12'h8D6: dout <= 8'b01111010; // 2262 : 122 - 0x7a
      12'h8D7: dout <= 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout <= 8'b11111100; // 2264 : 252 - 0xfc -- Background 0x1b
      12'h8D9: dout <= 8'b11000110; // 2265 : 198 - 0xc6
      12'h8DA: dout <= 8'b11000110; // 2266 : 198 - 0xc6
      12'h8DB: dout <= 8'b11001110; // 2267 : 206 - 0xce
      12'h8DC: dout <= 8'b11111000; // 2268 : 248 - 0xf8
      12'h8DD: dout <= 8'b11011100; // 2269 : 220 - 0xdc
      12'h8DE: dout <= 8'b11001110; // 2270 : 206 - 0xce
      12'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout <= 8'b01111000; // 2272 : 120 - 0x78 -- Background 0x1c
      12'h8E1: dout <= 8'b11001100; // 2273 : 204 - 0xcc
      12'h8E2: dout <= 8'b11000000; // 2274 : 192 - 0xc0
      12'h8E3: dout <= 8'b01111100; // 2275 : 124 - 0x7c
      12'h8E4: dout <= 8'b00000110; // 2276 :   6 - 0x6
      12'h8E5: dout <= 8'b11000110; // 2277 : 198 - 0xc6
      12'h8E6: dout <= 8'b01111100; // 2278 : 124 - 0x7c
      12'h8E7: dout <= 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout <= 8'b01111110; // 2280 : 126 - 0x7e -- Background 0x1d
      12'h8E9: dout <= 8'b00011000; // 2281 :  24 - 0x18
      12'h8EA: dout <= 8'b00011000; // 2282 :  24 - 0x18
      12'h8EB: dout <= 8'b00011000; // 2283 :  24 - 0x18
      12'h8EC: dout <= 8'b00011000; // 2284 :  24 - 0x18
      12'h8ED: dout <= 8'b00011000; // 2285 :  24 - 0x18
      12'h8EE: dout <= 8'b00011000; // 2286 :  24 - 0x18
      12'h8EF: dout <= 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout <= 8'b11000110; // 2288 : 198 - 0xc6 -- Background 0x1e
      12'h8F1: dout <= 8'b11000110; // 2289 : 198 - 0xc6
      12'h8F2: dout <= 8'b11000110; // 2290 : 198 - 0xc6
      12'h8F3: dout <= 8'b11000110; // 2291 : 198 - 0xc6
      12'h8F4: dout <= 8'b11000110; // 2292 : 198 - 0xc6
      12'h8F5: dout <= 8'b11000110; // 2293 : 198 - 0xc6
      12'h8F6: dout <= 8'b01111100; // 2294 : 124 - 0x7c
      12'h8F7: dout <= 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout <= 8'b11000110; // 2296 : 198 - 0xc6 -- Background 0x1f
      12'h8F9: dout <= 8'b11000110; // 2297 : 198 - 0xc6
      12'h8FA: dout <= 8'b11000110; // 2298 : 198 - 0xc6
      12'h8FB: dout <= 8'b11101110; // 2299 : 238 - 0xee
      12'h8FC: dout <= 8'b01111100; // 2300 : 124 - 0x7c
      12'h8FD: dout <= 8'b00111000; // 2301 :  56 - 0x38
      12'h8FE: dout <= 8'b00010000; // 2302 :  16 - 0x10
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b11000110; // 2304 : 198 - 0xc6 -- Background 0x20
      12'h901: dout <= 8'b11000110; // 2305 : 198 - 0xc6
      12'h902: dout <= 8'b11010110; // 2306 : 214 - 0xd6
      12'h903: dout <= 8'b11111110; // 2307 : 254 - 0xfe
      12'h904: dout <= 8'b11111110; // 2308 : 254 - 0xfe
      12'h905: dout <= 8'b11101110; // 2309 : 238 - 0xee
      12'h906: dout <= 8'b11000110; // 2310 : 198 - 0xc6
      12'h907: dout <= 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout <= 8'b11000110; // 2312 : 198 - 0xc6 -- Background 0x21
      12'h909: dout <= 8'b11101110; // 2313 : 238 - 0xee
      12'h90A: dout <= 8'b01111100; // 2314 : 124 - 0x7c
      12'h90B: dout <= 8'b00111000; // 2315 :  56 - 0x38
      12'h90C: dout <= 8'b01111100; // 2316 : 124 - 0x7c
      12'h90D: dout <= 8'b11101110; // 2317 : 238 - 0xee
      12'h90E: dout <= 8'b11000110; // 2318 : 198 - 0xc6
      12'h90F: dout <= 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout <= 8'b01100110; // 2320 : 102 - 0x66 -- Background 0x22
      12'h911: dout <= 8'b01100110; // 2321 : 102 - 0x66
      12'h912: dout <= 8'b01100110; // 2322 : 102 - 0x66
      12'h913: dout <= 8'b00111100; // 2323 :  60 - 0x3c
      12'h914: dout <= 8'b00011000; // 2324 :  24 - 0x18
      12'h915: dout <= 8'b00011000; // 2325 :  24 - 0x18
      12'h916: dout <= 8'b00011000; // 2326 :  24 - 0x18
      12'h917: dout <= 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout <= 8'b11111110; // 2328 : 254 - 0xfe -- Background 0x23
      12'h919: dout <= 8'b00001110; // 2329 :  14 - 0xe
      12'h91A: dout <= 8'b00011100; // 2330 :  28 - 0x1c
      12'h91B: dout <= 8'b00111000; // 2331 :  56 - 0x38
      12'h91C: dout <= 8'b01110000; // 2332 : 112 - 0x70
      12'h91D: dout <= 8'b11100000; // 2333 : 224 - 0xe0
      12'h91E: dout <= 8'b11111110; // 2334 : 254 - 0xfe
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout <= 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout <= 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout <= 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout <= 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout <= 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout <= 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0 -- Background 0x25
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00000110; // 2346 :   6 - 0x6
      12'h92B: dout <= 8'b00001110; // 2347 :  14 - 0xe
      12'h92C: dout <= 8'b00001000; // 2348 :   8 - 0x8
      12'h92D: dout <= 8'b00001000; // 2349 :   8 - 0x8
      12'h92E: dout <= 8'b00001000; // 2350 :   8 - 0x8
      12'h92F: dout <= 8'b00001000; // 2351 :   8 - 0x8
      12'h930: dout <= 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout <= 8'b01111000; // 2353 : 120 - 0x78
      12'h932: dout <= 8'b01100101; // 2354 : 101 - 0x65
      12'h933: dout <= 8'b01111001; // 2355 : 121 - 0x79
      12'h934: dout <= 8'b01100101; // 2356 : 101 - 0x65
      12'h935: dout <= 8'b01100101; // 2357 : 101 - 0x65
      12'h936: dout <= 8'b01111000; // 2358 : 120 - 0x78
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- Background 0x27
      12'h939: dout <= 8'b11100100; // 2361 : 228 - 0xe4
      12'h93A: dout <= 8'b10010110; // 2362 : 150 - 0x96
      12'h93B: dout <= 8'b10010110; // 2363 : 150 - 0x96
      12'h93C: dout <= 8'b10010111; // 2364 : 151 - 0x97
      12'h93D: dout <= 8'b10010110; // 2365 : 150 - 0x96
      12'h93E: dout <= 8'b11100110; // 2366 : 230 - 0xe6
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout <= 8'b01011001; // 2369 :  89 - 0x59
      12'h942: dout <= 8'b01011001; // 2370 :  89 - 0x59
      12'h943: dout <= 8'b01011001; // 2371 :  89 - 0x59
      12'h944: dout <= 8'b01011001; // 2372 :  89 - 0x59
      12'h945: dout <= 8'b11011001; // 2373 : 217 - 0xd9
      12'h946: dout <= 8'b01001110; // 2374 :  78 - 0x4e
      12'h947: dout <= 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- Background 0x29
      12'h949: dout <= 8'b00111100; // 2377 :  60 - 0x3c
      12'h94A: dout <= 8'b01110000; // 2378 : 112 - 0x70
      12'h94B: dout <= 8'b01110000; // 2379 : 112 - 0x70
      12'h94C: dout <= 8'b00111100; // 2380 :  60 - 0x3c
      12'h94D: dout <= 8'b00001100; // 2381 :  12 - 0xc
      12'h94E: dout <= 8'b01111000; // 2382 : 120 - 0x78
      12'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x2a
      12'h951: dout <= 8'b00000000; // 2385 :   0 - 0x0
      12'h952: dout <= 8'b11000110; // 2386 : 198 - 0xc6
      12'h953: dout <= 8'b11101110; // 2387 : 238 - 0xee
      12'h954: dout <= 8'b00101000; // 2388 :  40 - 0x28
      12'h955: dout <= 8'b00101000; // 2389 :  40 - 0x28
      12'h956: dout <= 8'b00101000; // 2390 :  40 - 0x28
      12'h957: dout <= 8'b00101000; // 2391 :  40 - 0x28
      12'h958: dout <= 8'b00001000; // 2392 :   8 - 0x8 -- Background 0x2b
      12'h959: dout <= 8'b00001000; // 2393 :   8 - 0x8
      12'h95A: dout <= 8'b00001000; // 2394 :   8 - 0x8
      12'h95B: dout <= 8'b00001000; // 2395 :   8 - 0x8
      12'h95C: dout <= 8'b00001110; // 2396 :  14 - 0xe
      12'h95D: dout <= 8'b00000110; // 2397 :   6 - 0x6
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00101000; // 2400 :  40 - 0x28 -- Background 0x2c
      12'h961: dout <= 8'b00101000; // 2401 :  40 - 0x28
      12'h962: dout <= 8'b00101000; // 2402 :  40 - 0x28
      12'h963: dout <= 8'b00101000; // 2403 :  40 - 0x28
      12'h964: dout <= 8'b11101110; // 2404 : 238 - 0xee
      12'h965: dout <= 8'b11000110; // 2405 : 198 - 0xc6
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- Background 0x2d
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b01100000; // 2410 :  96 - 0x60
      12'h96B: dout <= 8'b01110000; // 2411 : 112 - 0x70
      12'h96C: dout <= 8'b00010000; // 2412 :  16 - 0x10
      12'h96D: dout <= 8'b00010000; // 2413 :  16 - 0x10
      12'h96E: dout <= 8'b00010000; // 2414 :  16 - 0x10
      12'h96F: dout <= 8'b00010000; // 2415 :  16 - 0x10
      12'h970: dout <= 8'b00011100; // 2416 :  28 - 0x1c -- Background 0x2e
      12'h971: dout <= 8'b00111110; // 2417 :  62 - 0x3e
      12'h972: dout <= 8'b00111100; // 2418 :  60 - 0x3c
      12'h973: dout <= 8'b00111000; // 2419 :  56 - 0x38
      12'h974: dout <= 8'b00110000; // 2420 :  48 - 0x30
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b01100000; // 2422 :  96 - 0x60
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b00010000; // 2424 :  16 - 0x10 -- Background 0x2f
      12'h979: dout <= 8'b00010000; // 2425 :  16 - 0x10
      12'h97A: dout <= 8'b00010000; // 2426 :  16 - 0x10
      12'h97B: dout <= 8'b00010000; // 2427 :  16 - 0x10
      12'h97C: dout <= 8'b01110000; // 2428 : 112 - 0x70
      12'h97D: dout <= 8'b01100000; // 2429 :  96 - 0x60
      12'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Background 0x30
      12'h981: dout <= 8'b11111111; // 2433 : 255 - 0xff
      12'h982: dout <= 8'b00111000; // 2434 :  56 - 0x38
      12'h983: dout <= 8'b01101100; // 2435 : 108 - 0x6c
      12'h984: dout <= 8'b11000110; // 2436 : 198 - 0xc6
      12'h985: dout <= 8'b10000011; // 2437 : 131 - 0x83
      12'h986: dout <= 8'b11111111; // 2438 : 255 - 0xff
      12'h987: dout <= 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout <= 8'b11111111; // 2440 : 255 - 0xff -- Background 0x31
      12'h989: dout <= 8'b00111000; // 2441 :  56 - 0x38
      12'h98A: dout <= 8'b01101100; // 2442 : 108 - 0x6c
      12'h98B: dout <= 8'b11000110; // 2443 : 198 - 0xc6
      12'h98C: dout <= 8'b10000011; // 2444 : 131 - 0x83
      12'h98D: dout <= 8'b11111111; // 2445 : 255 - 0xff
      12'h98E: dout <= 8'b11111111; // 2446 : 255 - 0xff
      12'h98F: dout <= 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout <= 8'b00111000; // 2448 :  56 - 0x38 -- Background 0x32
      12'h991: dout <= 8'b01101100; // 2449 : 108 - 0x6c
      12'h992: dout <= 8'b11000110; // 2450 : 198 - 0xc6
      12'h993: dout <= 8'b10000011; // 2451 : 131 - 0x83
      12'h994: dout <= 8'b11111111; // 2452 : 255 - 0xff
      12'h995: dout <= 8'b11111111; // 2453 : 255 - 0xff
      12'h996: dout <= 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout <= 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout <= 8'b01101100; // 2456 : 108 - 0x6c -- Background 0x33
      12'h999: dout <= 8'b11000110; // 2457 : 198 - 0xc6
      12'h99A: dout <= 8'b10000011; // 2458 : 131 - 0x83
      12'h99B: dout <= 8'b11111111; // 2459 : 255 - 0xff
      12'h99C: dout <= 8'b11111111; // 2460 : 255 - 0xff
      12'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b11000110; // 2464 : 198 - 0xc6 -- Background 0x34
      12'h9A1: dout <= 8'b10000011; // 2465 : 131 - 0x83
      12'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout <= 8'b11111111; // 2467 : 255 - 0xff
      12'h9A4: dout <= 8'b00000000; // 2468 :   0 - 0x0
      12'h9A5: dout <= 8'b00000000; // 2469 :   0 - 0x0
      12'h9A6: dout <= 8'b00000000; // 2470 :   0 - 0x0
      12'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout <= 8'b10000011; // 2472 : 131 - 0x83 -- Background 0x35
      12'h9A9: dout <= 8'b11111111; // 2473 : 255 - 0xff
      12'h9AA: dout <= 8'b11111111; // 2474 : 255 - 0xff
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout <= 8'b11111111; // 2480 : 255 - 0xff -- Background 0x36
      12'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      12'h9B2: dout <= 8'b00000000; // 2482 :   0 - 0x0
      12'h9B3: dout <= 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout <= 8'b00000000; // 2484 :   0 - 0x0
      12'h9B5: dout <= 8'b00000000; // 2485 :   0 - 0x0
      12'h9B6: dout <= 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b11111111; // 2488 : 255 - 0xff -- Background 0x37
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b00000000; // 2492 :   0 - 0x0
      12'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout <= 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout <= 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout <= 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout <= 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout <= 8'b11111111; // 2503 : 255 - 0xff
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b11111111; // 2510 : 255 - 0xff
      12'h9CF: dout <= 8'b11111111; // 2511 : 255 - 0xff
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout <= 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout <= 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout <= 8'b11111111; // 2517 : 255 - 0xff
      12'h9D6: dout <= 8'b11111111; // 2518 : 255 - 0xff
      12'h9D7: dout <= 8'b00111000; // 2519 :  56 - 0x38
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b11111111; // 2524 : 255 - 0xff
      12'h9DD: dout <= 8'b11111111; // 2525 : 255 - 0xff
      12'h9DE: dout <= 8'b00111000; // 2526 :  56 - 0x38
      12'h9DF: dout <= 8'b01101100; // 2527 : 108 - 0x6c
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b11111111; // 2531 : 255 - 0xff
      12'h9E4: dout <= 8'b11111111; // 2532 : 255 - 0xff
      12'h9E5: dout <= 8'b00111000; // 2533 :  56 - 0x38
      12'h9E6: dout <= 8'b01101100; // 2534 : 108 - 0x6c
      12'h9E7: dout <= 8'b11000110; // 2535 : 198 - 0xc6
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b11111111; // 2538 : 255 - 0xff
      12'h9EB: dout <= 8'b11111111; // 2539 : 255 - 0xff
      12'h9EC: dout <= 8'b00111000; // 2540 :  56 - 0x38
      12'h9ED: dout <= 8'b01101100; // 2541 : 108 - 0x6c
      12'h9EE: dout <= 8'b11000110; // 2542 : 198 - 0xc6
      12'h9EF: dout <= 8'b10000011; // 2543 : 131 - 0x83
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b11111111; // 2545 : 255 - 0xff
      12'h9F2: dout <= 8'b11111111; // 2546 : 255 - 0xff
      12'h9F3: dout <= 8'b00111000; // 2547 :  56 - 0x38
      12'h9F4: dout <= 8'b01101100; // 2548 : 108 - 0x6c
      12'h9F5: dout <= 8'b11000110; // 2549 : 198 - 0xc6
      12'h9F6: dout <= 8'b10000011; // 2550 : 131 - 0x83
      12'h9F7: dout <= 8'b11111111; // 2551 : 255 - 0xff
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout <= 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout <= 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout <= 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout <= 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout <= 8'b11111111; // 2567 : 255 - 0xff
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b11111111; // 2573 : 255 - 0xff
      12'hA0E: dout <= 8'b11111111; // 2574 : 255 - 0xff
      12'hA0F: dout <= 8'b00111000; // 2575 :  56 - 0x38
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout <= 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout <= 8'b11111111; // 2580 : 255 - 0xff
      12'hA15: dout <= 8'b11111111; // 2581 : 255 - 0xff
      12'hA16: dout <= 8'b00111000; // 2582 :  56 - 0x38
      12'hA17: dout <= 8'b01101100; // 2583 : 108 - 0x6c
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b11111111; // 2587 : 255 - 0xff
      12'hA1C: dout <= 8'b11111111; // 2588 : 255 - 0xff
      12'hA1D: dout <= 8'b00111000; // 2589 :  56 - 0x38
      12'hA1E: dout <= 8'b01101100; // 2590 : 108 - 0x6c
      12'hA1F: dout <= 8'b11000110; // 2591 : 198 - 0xc6
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout <= 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout <= 8'b11111111; // 2594 : 255 - 0xff
      12'hA23: dout <= 8'b11111111; // 2595 : 255 - 0xff
      12'hA24: dout <= 8'b00111000; // 2596 :  56 - 0x38
      12'hA25: dout <= 8'b01101100; // 2597 : 108 - 0x6c
      12'hA26: dout <= 8'b11000110; // 2598 : 198 - 0xc6
      12'hA27: dout <= 8'b10000011; // 2599 : 131 - 0x83
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout <= 8'b11111111; // 2601 : 255 - 0xff
      12'hA2A: dout <= 8'b11111111; // 2602 : 255 - 0xff
      12'hA2B: dout <= 8'b00111000; // 2603 :  56 - 0x38
      12'hA2C: dout <= 8'b01101100; // 2604 : 108 - 0x6c
      12'hA2D: dout <= 8'b11000110; // 2605 : 198 - 0xc6
      12'hA2E: dout <= 8'b10000011; // 2606 : 131 - 0x83
      12'hA2F: dout <= 8'b11111111; // 2607 : 255 - 0xff
      12'hA30: dout <= 8'b11111111; // 2608 : 255 - 0xff -- Background 0x46
      12'hA31: dout <= 8'b00111000; // 2609 :  56 - 0x38
      12'hA32: dout <= 8'b01101100; // 2610 : 108 - 0x6c
      12'hA33: dout <= 8'b11000110; // 2611 : 198 - 0xc6
      12'hA34: dout <= 8'b10000011; // 2612 : 131 - 0x83
      12'hA35: dout <= 8'b11111111; // 2613 : 255 - 0xff
      12'hA36: dout <= 8'b11111111; // 2614 : 255 - 0xff
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00111000; // 2616 :  56 - 0x38 -- Background 0x47
      12'hA39: dout <= 8'b01101100; // 2617 : 108 - 0x6c
      12'hA3A: dout <= 8'b11000110; // 2618 : 198 - 0xc6
      12'hA3B: dout <= 8'b10000011; // 2619 : 131 - 0x83
      12'hA3C: dout <= 8'b11111111; // 2620 : 255 - 0xff
      12'hA3D: dout <= 8'b11111111; // 2621 : 255 - 0xff
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b01101100; // 2624 : 108 - 0x6c -- Background 0x48
      12'hA41: dout <= 8'b11000110; // 2625 : 198 - 0xc6
      12'hA42: dout <= 8'b10000011; // 2626 : 131 - 0x83
      12'hA43: dout <= 8'b11111111; // 2627 : 255 - 0xff
      12'hA44: dout <= 8'b11111111; // 2628 : 255 - 0xff
      12'hA45: dout <= 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout <= 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b11000110; // 2632 : 198 - 0xc6 -- Background 0x49
      12'hA49: dout <= 8'b10000011; // 2633 : 131 - 0x83
      12'hA4A: dout <= 8'b11111111; // 2634 : 255 - 0xff
      12'hA4B: dout <= 8'b11111111; // 2635 : 255 - 0xff
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b10000011; // 2640 : 131 - 0x83 -- Background 0x4a
      12'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout <= 8'b11111111; // 2642 : 255 - 0xff
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout <= 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout <= 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout <= 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout <= 8'b11111111; // 2648 : 255 - 0xff -- Background 0x4b
      12'hA59: dout <= 8'b11111111; // 2649 : 255 - 0xff
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b10111111; // 2656 : 191 - 0xbf -- Background 0x4c
      12'hA61: dout <= 8'b01011111; // 2657 :  95 - 0x5f
      12'hA62: dout <= 8'b01011111; // 2658 :  95 - 0x5f
      12'hA63: dout <= 8'b01011111; // 2659 :  95 - 0x5f
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b01011111; // 2661 :  95 - 0x5f
      12'hA66: dout <= 8'b01010001; // 2662 :  81 - 0x51
      12'hA67: dout <= 8'b01010101; // 2663 :  85 - 0x55
      12'hA68: dout <= 8'b01010001; // 2664 :  81 - 0x51 -- Background 0x4d
      12'hA69: dout <= 8'b01011111; // 2665 :  95 - 0x5f
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b01011111; // 2667 :  95 - 0x5f
      12'hA6C: dout <= 8'b01011111; // 2668 :  95 - 0x5f
      12'hA6D: dout <= 8'b01011111; // 2669 :  95 - 0x5f
      12'hA6E: dout <= 8'b01011111; // 2670 :  95 - 0x5f
      12'hA6F: dout <= 8'b10111111; // 2671 : 191 - 0xbf
      12'hA70: dout <= 8'b11111111; // 2672 : 255 - 0xff -- Background 0x4e
      12'hA71: dout <= 8'b11111110; // 2673 : 254 - 0xfe
      12'hA72: dout <= 8'b11111110; // 2674 : 254 - 0xfe
      12'hA73: dout <= 8'b11111110; // 2675 : 254 - 0xfe
      12'hA74: dout <= 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout <= 8'b11111110; // 2677 : 254 - 0xfe
      12'hA76: dout <= 8'b00100110; // 2678 :  38 - 0x26
      12'hA77: dout <= 8'b00100110; // 2679 :  38 - 0x26
      12'hA78: dout <= 8'b00100010; // 2680 :  34 - 0x22 -- Background 0x4f
      12'hA79: dout <= 8'b11111110; // 2681 : 254 - 0xfe
      12'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout <= 8'b11111110; // 2683 : 254 - 0xfe
      12'hA7C: dout <= 8'b11111110; // 2684 : 254 - 0xfe
      12'hA7D: dout <= 8'b11111110; // 2685 : 254 - 0xfe
      12'hA7E: dout <= 8'b11111110; // 2686 : 254 - 0xfe
      12'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout <= 8'b00000111; // 2688 :   7 - 0x7 -- Background 0x50
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00001111; // 2690 :  15 - 0xf
      12'hA83: dout <= 8'b00011111; // 2691 :  31 - 0x1f
      12'hA84: dout <= 8'b00011111; // 2692 :  31 - 0x1f
      12'hA85: dout <= 8'b00011111; // 2693 :  31 - 0x1f
      12'hA86: dout <= 8'b00011111; // 2694 :  31 - 0x1f
      12'hA87: dout <= 8'b00011111; // 2695 :  31 - 0x1f
      12'hA88: dout <= 8'b00011111; // 2696 :  31 - 0x1f -- Background 0x51
      12'hA89: dout <= 8'b00011111; // 2697 :  31 - 0x1f
      12'hA8A: dout <= 8'b00011111; // 2698 :  31 - 0x1f
      12'hA8B: dout <= 8'b00011111; // 2699 :  31 - 0x1f
      12'hA8C: dout <= 8'b00011111; // 2700 :  31 - 0x1f
      12'hA8D: dout <= 8'b00001111; // 2701 :  15 - 0xf
      12'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout <= 8'b00000111; // 2703 :   7 - 0x7
      12'hA90: dout <= 8'b00000111; // 2704 :   7 - 0x7 -- Background 0x52
      12'hA91: dout <= 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout <= 8'b00001111; // 2706 :  15 - 0xf
      12'hA93: dout <= 8'b00011111; // 2707 :  31 - 0x1f
      12'hA94: dout <= 8'b00011111; // 2708 :  31 - 0x1f
      12'hA95: dout <= 8'b00011111; // 2709 :  31 - 0x1f
      12'hA96: dout <= 8'b00011111; // 2710 :  31 - 0x1f
      12'hA97: dout <= 8'b00011111; // 2711 :  31 - 0x1f
      12'hA98: dout <= 8'b00011111; // 2712 :  31 - 0x1f -- Background 0x53
      12'hA99: dout <= 8'b00011111; // 2713 :  31 - 0x1f
      12'hA9A: dout <= 8'b00011111; // 2714 :  31 - 0x1f
      12'hA9B: dout <= 8'b00011111; // 2715 :  31 - 0x1f
      12'hA9C: dout <= 8'b00011111; // 2716 :  31 - 0x1f
      12'hA9D: dout <= 8'b00001111; // 2717 :  15 - 0xf
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000111; // 2719 :   7 - 0x7
      12'hAA0: dout <= 8'b11100000; // 2720 : 224 - 0xe0 -- Background 0x54
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b11110001; // 2722 : 241 - 0xf1
      12'hAA3: dout <= 8'b11111011; // 2723 : 251 - 0xfb
      12'hAA4: dout <= 8'b11111011; // 2724 : 251 - 0xfb
      12'hAA5: dout <= 8'b11111011; // 2725 : 251 - 0xfb
      12'hAA6: dout <= 8'b11111011; // 2726 : 251 - 0xfb
      12'hAA7: dout <= 8'b11111011; // 2727 : 251 - 0xfb
      12'hAA8: dout <= 8'b11111011; // 2728 : 251 - 0xfb -- Background 0x55
      12'hAA9: dout <= 8'b11111011; // 2729 : 251 - 0xfb
      12'hAAA: dout <= 8'b11111011; // 2730 : 251 - 0xfb
      12'hAAB: dout <= 8'b11111011; // 2731 : 251 - 0xfb
      12'hAAC: dout <= 8'b11111011; // 2732 : 251 - 0xfb
      12'hAAD: dout <= 8'b11110001; // 2733 : 241 - 0xf1
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b11100000; // 2735 : 224 - 0xe0
      12'hAB0: dout <= 8'b11100000; // 2736 : 224 - 0xe0 -- Background 0x56
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b11110001; // 2738 : 241 - 0xf1
      12'hAB3: dout <= 8'b11111011; // 2739 : 251 - 0xfb
      12'hAB4: dout <= 8'b11111011; // 2740 : 251 - 0xfb
      12'hAB5: dout <= 8'b11111011; // 2741 : 251 - 0xfb
      12'hAB6: dout <= 8'b11111011; // 2742 : 251 - 0xfb
      12'hAB7: dout <= 8'b11111011; // 2743 : 251 - 0xfb
      12'hAB8: dout <= 8'b11111011; // 2744 : 251 - 0xfb -- Background 0x57
      12'hAB9: dout <= 8'b11111011; // 2745 : 251 - 0xfb
      12'hABA: dout <= 8'b11111011; // 2746 : 251 - 0xfb
      12'hABB: dout <= 8'b11111011; // 2747 : 251 - 0xfb
      12'hABC: dout <= 8'b11111011; // 2748 : 251 - 0xfb
      12'hABD: dout <= 8'b11110001; // 2749 : 241 - 0xf1
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b11100000; // 2751 : 224 - 0xe0
      12'hAC0: dout <= 8'b11111100; // 2752 : 252 - 0xfc -- Background 0x58
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b11111110; // 2754 : 254 - 0xfe
      12'hAC3: dout <= 8'b11111111; // 2755 : 255 - 0xff
      12'hAC4: dout <= 8'b11111111; // 2756 : 255 - 0xff
      12'hAC5: dout <= 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout <= 8'b11111111; // 2758 : 255 - 0xff
      12'hAC7: dout <= 8'b11111111; // 2759 : 255 - 0xff
      12'hAC8: dout <= 8'b11111111; // 2760 : 255 - 0xff -- Background 0x59
      12'hAC9: dout <= 8'b11111111; // 2761 : 255 - 0xff
      12'hACA: dout <= 8'b11111111; // 2762 : 255 - 0xff
      12'hACB: dout <= 8'b11111111; // 2763 : 255 - 0xff
      12'hACC: dout <= 8'b11111111; // 2764 : 255 - 0xff
      12'hACD: dout <= 8'b11111110; // 2765 : 254 - 0xfe
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b11111100; // 2767 : 252 - 0xfc
      12'hAD0: dout <= 8'b11111100; // 2768 : 252 - 0xfc -- Background 0x5a
      12'hAD1: dout <= 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout <= 8'b11111110; // 2770 : 254 - 0xfe
      12'hAD3: dout <= 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout <= 8'b11111111; // 2772 : 255 - 0xff
      12'hAD5: dout <= 8'b11111111; // 2773 : 255 - 0xff
      12'hAD6: dout <= 8'b11111111; // 2774 : 255 - 0xff
      12'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      12'hAD8: dout <= 8'b11111111; // 2776 : 255 - 0xff -- Background 0x5b
      12'hAD9: dout <= 8'b11111111; // 2777 : 255 - 0xff
      12'hADA: dout <= 8'b11111111; // 2778 : 255 - 0xff
      12'hADB: dout <= 8'b11111111; // 2779 : 255 - 0xff
      12'hADC: dout <= 8'b11111111; // 2780 : 255 - 0xff
      12'hADD: dout <= 8'b11111110; // 2781 : 254 - 0xfe
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b11111100; // 2783 : 252 - 0xfc
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00011111; // 2786 :  31 - 0x1f
      12'hAE3: dout <= 8'b00010000; // 2787 :  16 - 0x10
      12'hAE4: dout <= 8'b00010000; // 2788 :  16 - 0x10
      12'hAE5: dout <= 8'b00011111; // 2789 :  31 - 0x1f
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b11111000; // 2794 : 248 - 0xf8
      12'hAEB: dout <= 8'b00001000; // 2795 :   8 - 0x8
      12'hAEC: dout <= 8'b00001000; // 2796 :   8 - 0x8
      12'hAED: dout <= 8'b11111000; // 2797 : 248 - 0xf8
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout <= 8'b00000001; // 2801 :   1 - 0x1
      12'hAF2: dout <= 8'b00000010; // 2802 :   2 - 0x2
      12'hAF3: dout <= 8'b00000010; // 2803 :   2 - 0x2
      12'hAF4: dout <= 8'b11110001; // 2804 : 241 - 0xf1
      12'hAF5: dout <= 8'b00001000; // 2805 :   8 - 0x8
      12'hAF6: dout <= 8'b00000100; // 2806 :   4 - 0x4
      12'hAF7: dout <= 8'b00000011; // 2807 :   3 - 0x3
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout <= 8'b10000000; // 2809 : 128 - 0x80
      12'hAFA: dout <= 8'b01000000; // 2810 :  64 - 0x40
      12'hAFB: dout <= 8'b01000000; // 2811 :  64 - 0x40
      12'hAFC: dout <= 8'b10001111; // 2812 : 143 - 0x8f
      12'hAFD: dout <= 8'b00010000; // 2813 :  16 - 0x10
      12'hAFE: dout <= 8'b00100000; // 2814 :  32 - 0x20
      12'hAFF: dout <= 8'b11000000; // 2815 : 192 - 0xc0
      12'hB00: dout <= 8'b00000011; // 2816 :   3 - 0x3 -- Background 0x60
      12'hB01: dout <= 8'b00000100; // 2817 :   4 - 0x4
      12'hB02: dout <= 8'b00001000; // 2818 :   8 - 0x8
      12'hB03: dout <= 8'b11110001; // 2819 : 241 - 0xf1
      12'hB04: dout <= 8'b00000010; // 2820 :   2 - 0x2
      12'hB05: dout <= 8'b00000010; // 2821 :   2 - 0x2
      12'hB06: dout <= 8'b00000001; // 2822 :   1 - 0x1
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b11000000; // 2824 : 192 - 0xc0 -- Background 0x61
      12'hB09: dout <= 8'b00100000; // 2825 :  32 - 0x20
      12'hB0A: dout <= 8'b00010000; // 2826 :  16 - 0x10
      12'hB0B: dout <= 8'b10001111; // 2827 : 143 - 0x8f
      12'hB0C: dout <= 8'b01000000; // 2828 :  64 - 0x40
      12'hB0D: dout <= 8'b01000000; // 2829 :  64 - 0x40
      12'hB0E: dout <= 8'b10000000; // 2830 : 128 - 0x80
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b11111111; // 2832 : 255 - 0xff -- Background 0x62
      12'hB11: dout <= 8'b11111111; // 2833 : 255 - 0xff
      12'hB12: dout <= 8'b11000011; // 2834 : 195 - 0xc3
      12'hB13: dout <= 8'b10000001; // 2835 : 129 - 0x81
      12'hB14: dout <= 8'b10000001; // 2836 : 129 - 0x81
      12'hB15: dout <= 8'b11000011; // 2837 : 195 - 0xc3
      12'hB16: dout <= 8'b11111111; // 2838 : 255 - 0xff
      12'hB17: dout <= 8'b11111111; // 2839 : 255 - 0xff
      12'hB18: dout <= 8'b11111111; // 2840 : 255 - 0xff -- Background 0x63
      12'hB19: dout <= 8'b10011001; // 2841 : 153 - 0x99
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b10000001; // 2845 : 129 - 0x81
      12'hB1E: dout <= 8'b10000001; // 2846 : 129 - 0x81
      12'hB1F: dout <= 8'b10000001; // 2847 : 129 - 0x81
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout <= 8'b01100000; // 2852 :  96 - 0x60
      12'hB25: dout <= 8'b01100000; // 2853 :  96 - 0x60
      12'hB26: dout <= 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- Background 0x65
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout <= 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout <= 8'b01101100; // 2860 : 108 - 0x6c
      12'hB2D: dout <= 8'b01101100; // 2861 : 108 - 0x6c
      12'hB2E: dout <= 8'b00001000; // 2862 :   8 - 0x8
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00111100; // 2864 :  60 - 0x3c -- Background 0x66
      12'hB31: dout <= 8'b00011000; // 2865 :  24 - 0x18
      12'hB32: dout <= 8'b00011000; // 2866 :  24 - 0x18
      12'hB33: dout <= 8'b00011000; // 2867 :  24 - 0x18
      12'hB34: dout <= 8'b00011000; // 2868 :  24 - 0x18
      12'hB35: dout <= 8'b00011000; // 2869 :  24 - 0x18
      12'hB36: dout <= 8'b00111100; // 2870 :  60 - 0x3c
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b11111111; // 2872 : 255 - 0xff -- Background 0x67
      12'hB39: dout <= 8'b01100110; // 2873 : 102 - 0x66
      12'hB3A: dout <= 8'b01100110; // 2874 : 102 - 0x66
      12'hB3B: dout <= 8'b01100110; // 2875 : 102 - 0x66
      12'hB3C: dout <= 8'b01100110; // 2876 : 102 - 0x66
      12'hB3D: dout <= 8'b01100110; // 2877 : 102 - 0x66
      12'hB3E: dout <= 8'b01100110; // 2878 : 102 - 0x66
      12'hB3F: dout <= 8'b11111111; // 2879 : 255 - 0xff
      12'hB40: dout <= 8'b00000011; // 2880 :   3 - 0x3 -- Background 0x68
      12'hB41: dout <= 8'b00000001; // 2881 :   1 - 0x1
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b10000011; // 2888 : 131 - 0x83 -- Background 0x69
      12'hB49: dout <= 8'b11010001; // 2889 : 209 - 0xd1
      12'hB4A: dout <= 8'b11100001; // 2890 : 225 - 0xe1
      12'hB4B: dout <= 8'b11010001; // 2891 : 209 - 0xd1
      12'hB4C: dout <= 8'b00000010; // 2892 :   2 - 0x2
      12'hB4D: dout <= 8'b10000100; // 2893 : 132 - 0x84
      12'hB4E: dout <= 8'b11110000; // 2894 : 240 - 0xf0
      12'hB4F: dout <= 8'b11001110; // 2895 : 206 - 0xce
      12'hB50: dout <= 8'b11000000; // 2896 : 192 - 0xc0 -- Background 0x6a
      12'hB51: dout <= 8'b10000000; // 2897 : 128 - 0x80
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b11000001; // 2904 : 193 - 0xc1 -- Background 0x6b
      12'hB59: dout <= 8'b10001011; // 2905 : 139 - 0x8b
      12'hB5A: dout <= 8'b10000111; // 2906 : 135 - 0x87
      12'hB5B: dout <= 8'b10001011; // 2907 : 139 - 0x8b
      12'hB5C: dout <= 8'b01000000; // 2908 :  64 - 0x40
      12'hB5D: dout <= 8'b00100001; // 2909 :  33 - 0x21
      12'hB5E: dout <= 8'b00001111; // 2910 :  15 - 0xf
      12'hB5F: dout <= 8'b11010011; // 2911 : 211 - 0xd3
      12'hB60: dout <= 8'b11111111; // 2912 : 255 - 0xff -- Background 0x6c
      12'hB61: dout <= 8'b11111111; // 2913 : 255 - 0xff
      12'hB62: dout <= 8'b11111111; // 2914 : 255 - 0xff
      12'hB63: dout <= 8'b00011111; // 2915 :  31 - 0x1f
      12'hB64: dout <= 8'b00001111; // 2916 :  15 - 0xf
      12'hB65: dout <= 8'b00011110; // 2917 :  30 - 0x1e
      12'hB66: dout <= 8'b00111111; // 2918 :  63 - 0x3f
      12'hB67: dout <= 8'b01111111; // 2919 : 127 - 0x7f
      12'hB68: dout <= 8'b11111111; // 2920 : 255 - 0xff -- Background 0x6d
      12'hB69: dout <= 8'b11111111; // 2921 : 255 - 0xff
      12'hB6A: dout <= 8'b11111111; // 2922 : 255 - 0xff
      12'hB6B: dout <= 8'b11111000; // 2923 : 248 - 0xf8
      12'hB6C: dout <= 8'b11110000; // 2924 : 240 - 0xf0
      12'hB6D: dout <= 8'b01111000; // 2925 : 120 - 0x78
      12'hB6E: dout <= 8'b11111100; // 2926 : 252 - 0xfc
      12'hB6F: dout <= 8'b11111110; // 2927 : 254 - 0xfe
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00111100; // 2933 :  60 - 0x3c
      12'hB76: dout <= 8'b01000010; // 2934 :  66 - 0x42
      12'hB77: dout <= 8'b10000001; // 2935 : 129 - 0x81
      12'hB78: dout <= 8'b10000001; // 2936 : 129 - 0x81 -- Background 0x6f
      12'hB79: dout <= 8'b10111101; // 2937 : 189 - 0xbd
      12'hB7A: dout <= 8'b01111110; // 2938 : 126 - 0x7e
      12'hB7B: dout <= 8'b11111111; // 2939 : 255 - 0xff
      12'hB7C: dout <= 8'b11100111; // 2940 : 231 - 0xe7
      12'hB7D: dout <= 8'b11111111; // 2941 : 255 - 0xff
      12'hB7E: dout <= 8'b11111111; // 2942 : 255 - 0xff
      12'hB7F: dout <= 8'b11111111; // 2943 : 255 - 0xff
      12'hB80: dout <= 8'b00000001; // 2944 :   1 - 0x1 -- Background 0x70
      12'hB81: dout <= 8'b00000111; // 2945 :   7 - 0x7
      12'hB82: dout <= 8'b00011111; // 2946 :  31 - 0x1f
      12'hB83: dout <= 8'b00111111; // 2947 :  63 - 0x3f
      12'hB84: dout <= 8'b01111111; // 2948 : 127 - 0x7f
      12'hB85: dout <= 8'b11111111; // 2949 : 255 - 0xff
      12'hB86: dout <= 8'b11111111; // 2950 : 255 - 0xff
      12'hB87: dout <= 8'b11011101; // 2951 : 221 - 0xdd
      12'hB88: dout <= 8'b10001001; // 2952 : 137 - 0x89 -- Background 0x71
      12'hB89: dout <= 8'b00000001; // 2953 :   1 - 0x1
      12'hB8A: dout <= 8'b00000001; // 2954 :   1 - 0x1
      12'hB8B: dout <= 8'b00000001; // 2955 :   1 - 0x1
      12'hB8C: dout <= 8'b00000001; // 2956 :   1 - 0x1
      12'hB8D: dout <= 8'b00000001; // 2957 :   1 - 0x1
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b10000000; // 2960 : 128 - 0x80 -- Background 0x72
      12'hB91: dout <= 8'b11100000; // 2961 : 224 - 0xe0
      12'hB92: dout <= 8'b11111000; // 2962 : 248 - 0xf8
      12'hB93: dout <= 8'b11111100; // 2963 : 252 - 0xfc
      12'hB94: dout <= 8'b11111110; // 2964 : 254 - 0xfe
      12'hB95: dout <= 8'b11111111; // 2965 : 255 - 0xff
      12'hB96: dout <= 8'b11111111; // 2966 : 255 - 0xff
      12'hB97: dout <= 8'b00111011; // 2967 :  59 - 0x3b
      12'hB98: dout <= 8'b00010001; // 2968 :  17 - 0x11 -- Background 0x73
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b01000000; // 2973 :  64 - 0x40
      12'hB9E: dout <= 8'b10000000; // 2974 : 128 - 0x80
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000001; // 2976 :   1 - 0x1 -- Background 0x74
      12'hBA1: dout <= 8'b00000001; // 2977 :   1 - 0x1
      12'hBA2: dout <= 8'b00000001; // 2978 :   1 - 0x1
      12'hBA3: dout <= 8'b00000001; // 2979 :   1 - 0x1
      12'hBA4: dout <= 8'b00000001; // 2980 :   1 - 0x1
      12'hBA5: dout <= 8'b00000001; // 2981 :   1 - 0x1
      12'hBA6: dout <= 8'b00000001; // 2982 :   1 - 0x1
      12'hBA7: dout <= 8'b00000001; // 2983 :   1 - 0x1
      12'hBA8: dout <= 8'b10000000; // 2984 : 128 - 0x80 -- Background 0x75
      12'hBA9: dout <= 8'b10000000; // 2985 : 128 - 0x80
      12'hBAA: dout <= 8'b10000000; // 2986 : 128 - 0x80
      12'hBAB: dout <= 8'b10000000; // 2987 : 128 - 0x80
      12'hBAC: dout <= 8'b10000000; // 2988 : 128 - 0x80
      12'hBAD: dout <= 8'b10000000; // 2989 : 128 - 0x80
      12'hBAE: dout <= 8'b10000000; // 2990 : 128 - 0x80
      12'hBAF: dout <= 8'b10000000; // 2991 : 128 - 0x80
      12'hBB0: dout <= 8'b00000001; // 2992 :   1 - 0x1 -- Background 0x76
      12'hBB1: dout <= 8'b00000011; // 2993 :   3 - 0x3
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000011; // 2996 :   3 - 0x3
      12'hBB5: dout <= 8'b00011001; // 2997 :  25 - 0x19
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b01111100; // 3002 : 124 - 0x7c
      12'hBBB: dout <= 8'b00000010; // 3003 :   2 - 0x2
      12'hBBC: dout <= 8'b00000001; // 3004 :   1 - 0x1
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000001; // 3010 :   1 - 0x1
      12'hBC3: dout <= 8'b00000001; // 3011 :   1 - 0x1
      12'hBC4: dout <= 8'b00000011; // 3012 :   3 - 0x3
      12'hBC5: dout <= 8'b00000111; // 3013 :   7 - 0x7
      12'hBC6: dout <= 8'b00000111; // 3014 :   7 - 0x7
      12'hBC7: dout <= 8'b00001111; // 3015 :  15 - 0xf
      12'hBC8: dout <= 8'b00001111; // 3016 :  15 - 0xf -- Background 0x79
      12'hBC9: dout <= 8'b00000111; // 3017 :   7 - 0x7
      12'hBCA: dout <= 8'b00001111; // 3018 :  15 - 0xf
      12'hBCB: dout <= 8'b00000111; // 3019 :   7 - 0x7
      12'hBCC: dout <= 8'b00000001; // 3020 :   1 - 0x1
      12'hBCD: dout <= 8'b00010000; // 3021 :  16 - 0x10
      12'hBCE: dout <= 8'b00100000; // 3022 :  32 - 0x20
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b11111000; // 3024 : 248 - 0xf8 -- Background 0x7a
      12'hBD1: dout <= 8'b11111110; // 3025 : 254 - 0xfe
      12'hBD2: dout <= 8'b01111111; // 3026 : 127 - 0x7f
      12'hBD3: dout <= 8'b00011111; // 3027 :  31 - 0x1f
      12'hBD4: dout <= 8'b00001111; // 3028 :  15 - 0xf
      12'hBD5: dout <= 8'b00011001; // 3029 :  25 - 0x19
      12'hBD6: dout <= 8'b00110000; // 3030 :  48 - 0x30
      12'hBD7: dout <= 8'b01110000; // 3031 : 112 - 0x70
      12'hBD8: dout <= 8'b11111011; // 3032 : 251 - 0xfb -- Background 0x7b
      12'hBD9: dout <= 8'b01110011; // 3033 : 115 - 0x73
      12'hBDA: dout <= 8'b00100111; // 3034 :  39 - 0x27
      12'hBDB: dout <= 8'b00001111; // 3035 :  15 - 0xf
      12'hBDC: dout <= 8'b00011111; // 3036 :  31 - 0x1f
      12'hBDD: dout <= 8'b00011111; // 3037 :  31 - 0x1f
      12'hBDE: dout <= 8'b00111111; // 3038 :  63 - 0x3f
      12'hBDF: dout <= 8'b01111111; // 3039 : 127 - 0x7f
      12'hBE0: dout <= 8'b11111111; // 3040 : 255 - 0xff -- Background 0x7c
      12'hBE1: dout <= 8'b11111111; // 3041 : 255 - 0xff
      12'hBE2: dout <= 8'b11111111; // 3042 : 255 - 0xff
      12'hBE3: dout <= 8'b11111111; // 3043 : 255 - 0xff
      12'hBE4: dout <= 8'b11111110; // 3044 : 254 - 0xfe
      12'hBE5: dout <= 8'b11111101; // 3045 : 253 - 0xfd
      12'hBE6: dout <= 8'b11111000; // 3046 : 248 - 0xf8
      12'hBE7: dout <= 8'b11110110; // 3047 : 246 - 0xf6
      12'hBE8: dout <= 8'b11101111; // 3048 : 239 - 0xef -- Background 0x7d
      12'hBE9: dout <= 8'b11001111; // 3049 : 207 - 0xcf
      12'hBEA: dout <= 8'b10011111; // 3050 : 159 - 0x9f
      12'hBEB: dout <= 8'b00011111; // 3051 :  31 - 0x1f
      12'hBEC: dout <= 8'b00001111; // 3052 :  15 - 0xf
      12'hBED: dout <= 8'b00101101; // 3053 :  45 - 0x2d
      12'hBEE: dout <= 8'b01010000; // 3054 :  80 - 0x50
      12'hBEF: dout <= 8'b01000000; // 3055 :  64 - 0x40
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0x7e
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b11100000; // 3060 : 224 - 0xe0
      12'hBF5: dout <= 8'b11111110; // 3061 : 254 - 0xfe
      12'hBF6: dout <= 8'b11111111; // 3062 : 255 - 0xff
      12'hBF7: dout <= 8'b11110011; // 3063 : 243 - 0xf3
      12'hBF8: dout <= 8'b11111011; // 3064 : 251 - 0xfb -- Background 0x7f
      12'hBF9: dout <= 8'b11111011; // 3065 : 251 - 0xfb
      12'hBFA: dout <= 8'b11111011; // 3066 : 251 - 0xfb
      12'hBFB: dout <= 8'b11111011; // 3067 : 251 - 0xfb
      12'hBFC: dout <= 8'b11111011; // 3068 : 251 - 0xfb
      12'hBFD: dout <= 8'b11110011; // 3069 : 243 - 0xf3
      12'hBFE: dout <= 8'b11110111; // 3070 : 247 - 0xf7
      12'hBFF: dout <= 8'b11100111; // 3071 : 231 - 0xe7
      12'hC00: dout <= 8'b11001111; // 3072 : 207 - 0xcf -- Background 0x80
      12'hC01: dout <= 8'b10011111; // 3073 : 159 - 0x9f
      12'hC02: dout <= 8'b00111111; // 3074 :  63 - 0x3f
      12'hC03: dout <= 8'b00111111; // 3075 :  63 - 0x3f
      12'hC04: dout <= 8'b00111111; // 3076 :  63 - 0x3f
      12'hC05: dout <= 8'b00001111; // 3077 :  15 - 0xf
      12'hC06: dout <= 8'b00000011; // 3078 :   3 - 0x3
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b11000000; // 3080 : 192 - 0xc0 -- Background 0x81
      12'hC09: dout <= 8'b11110000; // 3081 : 240 - 0xf0
      12'hC0A: dout <= 8'b11111100; // 3082 : 252 - 0xfc
      12'hC0B: dout <= 8'b11110000; // 3083 : 240 - 0xf0
      12'hC0C: dout <= 8'b11110000; // 3084 : 240 - 0xf0
      12'hC0D: dout <= 8'b10011000; // 3085 : 152 - 0x98
      12'hC0E: dout <= 8'b00001000; // 3086 :   8 - 0x8
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00000000; // 3088 :   0 - 0x0 -- Background 0x82
      12'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout <= 8'b10000000; // 3094 : 128 - 0x80
      12'hC17: dout <= 8'b11000000; // 3095 : 192 - 0xc0
      12'hC18: dout <= 8'b11100000; // 3096 : 224 - 0xe0 -- Background 0x83
      12'hC19: dout <= 8'b11100000; // 3097 : 224 - 0xe0
      12'hC1A: dout <= 8'b11110000; // 3098 : 240 - 0xf0
      12'hC1B: dout <= 8'b11110000; // 3099 : 240 - 0xf0
      12'hC1C: dout <= 8'b11110000; // 3100 : 240 - 0xf0
      12'hC1D: dout <= 8'b11110000; // 3101 : 240 - 0xf0
      12'hC1E: dout <= 8'b11111000; // 3102 : 248 - 0xf8
      12'hC1F: dout <= 8'b11111000; // 3103 : 248 - 0xf8
      12'hC20: dout <= 8'b11111110; // 3104 : 254 - 0xfe -- Background 0x84
      12'hC21: dout <= 8'b11111111; // 3105 : 255 - 0xff
      12'hC22: dout <= 8'b11111111; // 3106 : 255 - 0xff
      12'hC23: dout <= 8'b11111111; // 3107 : 255 - 0xff
      12'hC24: dout <= 8'b11111111; // 3108 : 255 - 0xff
      12'hC25: dout <= 8'b11111111; // 3109 : 255 - 0xff
      12'hC26: dout <= 8'b11111111; // 3110 : 255 - 0xff
      12'hC27: dout <= 8'b11111111; // 3111 : 255 - 0xff
      12'hC28: dout <= 8'b00111111; // 3112 :  63 - 0x3f -- Background 0x85
      12'hC29: dout <= 8'b00011111; // 3113 :  31 - 0x1f
      12'hC2A: dout <= 8'b00011111; // 3114 :  31 - 0x1f
      12'hC2B: dout <= 8'b00001111; // 3115 :  15 - 0xf
      12'hC2C: dout <= 8'b00000111; // 3116 :   7 - 0x7
      12'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Background 0x86
      12'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout <= 8'b11000000; // 3122 : 192 - 0xc0
      12'hC33: dout <= 8'b11100000; // 3123 : 224 - 0xe0
      12'hC34: dout <= 8'b11110000; // 3124 : 240 - 0xf0
      12'hC35: dout <= 8'b11110000; // 3125 : 240 - 0xf0
      12'hC36: dout <= 8'b11110000; // 3126 : 240 - 0xf0
      12'hC37: dout <= 8'b11111000; // 3127 : 248 - 0xf8
      12'hC38: dout <= 8'b11111001; // 3128 : 249 - 0xf9 -- Background 0x87
      12'hC39: dout <= 8'b11111111; // 3129 : 255 - 0xff
      12'hC3A: dout <= 8'b11111111; // 3130 : 255 - 0xff
      12'hC3B: dout <= 8'b11111111; // 3131 : 255 - 0xff
      12'hC3C: dout <= 8'b11111111; // 3132 : 255 - 0xff
      12'hC3D: dout <= 8'b00001110; // 3133 :  14 - 0xe
      12'hC3E: dout <= 8'b00000010; // 3134 :   2 - 0x2
      12'hC3F: dout <= 8'b00010100; // 3135 :  20 - 0x14
      12'hC40: dout <= 8'b10000000; // 3136 : 128 - 0x80 -- Background 0x88
      12'hC41: dout <= 8'b10100000; // 3137 : 160 - 0xa0
      12'hC42: dout <= 8'b00100000; // 3138 :  32 - 0x20
      12'hC43: dout <= 8'b00100000; // 3139 :  32 - 0x20
      12'hC44: dout <= 8'b10100000; // 3140 : 160 - 0xa0
      12'hC45: dout <= 8'b10000000; // 3141 : 128 - 0x80
      12'hC46: dout <= 8'b00000000; // 3142 :   0 - 0x0
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00000001; // 3144 :   1 - 0x1 -- Background 0x89
      12'hC49: dout <= 8'b00000101; // 3145 :   5 - 0x5
      12'hC4A: dout <= 8'b00000100; // 3146 :   4 - 0x4
      12'hC4B: dout <= 8'b00000100; // 3147 :   4 - 0x4
      12'hC4C: dout <= 8'b00000101; // 3148 :   5 - 0x5
      12'hC4D: dout <= 8'b00000001; // 3149 :   1 - 0x1
      12'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Background 0x8a
      12'hC51: dout <= 8'b00000000; // 3153 :   0 - 0x0
      12'hC52: dout <= 8'b00000011; // 3154 :   3 - 0x3
      12'hC53: dout <= 8'b00000111; // 3155 :   7 - 0x7
      12'hC54: dout <= 8'b00001111; // 3156 :  15 - 0xf
      12'hC55: dout <= 8'b00001111; // 3157 :  15 - 0xf
      12'hC56: dout <= 8'b00001111; // 3158 :  15 - 0xf
      12'hC57: dout <= 8'b00001111; // 3159 :  15 - 0xf
      12'hC58: dout <= 8'b10011111; // 3160 : 159 - 0x9f -- Background 0x8b
      12'hC59: dout <= 8'b11111111; // 3161 : 255 - 0xff
      12'hC5A: dout <= 8'b11111111; // 3162 : 255 - 0xff
      12'hC5B: dout <= 8'b11111111; // 3163 : 255 - 0xff
      12'hC5C: dout <= 8'b11111111; // 3164 : 255 - 0xff
      12'hC5D: dout <= 8'b01110000; // 3165 : 112 - 0x70
      12'hC5E: dout <= 8'b01000000; // 3166 :  64 - 0x40
      12'hC5F: dout <= 8'b00101000; // 3167 :  40 - 0x28
      12'hC60: dout <= 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout <= 8'b00000000; // 3169 :   0 - 0x0
      12'hC62: dout <= 8'b00000000; // 3170 :   0 - 0x0
      12'hC63: dout <= 8'b00000000; // 3171 :   0 - 0x0
      12'hC64: dout <= 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout <= 8'b00000000; // 3173 :   0 - 0x0
      12'hC66: dout <= 8'b00000001; // 3174 :   1 - 0x1
      12'hC67: dout <= 8'b00000011; // 3175 :   3 - 0x3
      12'hC68: dout <= 8'b00000111; // 3176 :   7 - 0x7 -- Background 0x8d
      12'hC69: dout <= 8'b00000111; // 3177 :   7 - 0x7
      12'hC6A: dout <= 8'b00001111; // 3178 :  15 - 0xf
      12'hC6B: dout <= 8'b00001111; // 3179 :  15 - 0xf
      12'hC6C: dout <= 8'b00001111; // 3180 :  15 - 0xf
      12'hC6D: dout <= 8'b00001111; // 3181 :  15 - 0xf
      12'hC6E: dout <= 8'b00011111; // 3182 :  31 - 0x1f
      12'hC6F: dout <= 8'b00011111; // 3183 :  31 - 0x1f
      12'hC70: dout <= 8'b01111111; // 3184 : 127 - 0x7f -- Background 0x8e
      12'hC71: dout <= 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout <= 8'b11111111; // 3186 : 255 - 0xff
      12'hC73: dout <= 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout <= 8'b11111111; // 3188 : 255 - 0xff
      12'hC75: dout <= 8'b11111111; // 3189 : 255 - 0xff
      12'hC76: dout <= 8'b11111111; // 3190 : 255 - 0xff
      12'hC77: dout <= 8'b11111111; // 3191 : 255 - 0xff
      12'hC78: dout <= 8'b11111100; // 3192 : 252 - 0xfc -- Background 0x8f
      12'hC79: dout <= 8'b11111000; // 3193 : 248 - 0xf8
      12'hC7A: dout <= 8'b11111000; // 3194 : 248 - 0xf8
      12'hC7B: dout <= 8'b11110000; // 3195 : 240 - 0xf0
      12'hC7C: dout <= 8'b11100000; // 3196 : 224 - 0xe0
      12'hC7D: dout <= 8'b00000000; // 3197 :   0 - 0x0
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000111; // 3204 :   7 - 0x7
      12'hC85: dout <= 8'b01111111; // 3205 : 127 - 0x7f
      12'hC86: dout <= 8'b11111111; // 3206 : 255 - 0xff
      12'hC87: dout <= 8'b11001111; // 3207 : 207 - 0xcf
      12'hC88: dout <= 8'b11011111; // 3208 : 223 - 0xdf -- Background 0x91
      12'hC89: dout <= 8'b11011111; // 3209 : 223 - 0xdf
      12'hC8A: dout <= 8'b11011111; // 3210 : 223 - 0xdf
      12'hC8B: dout <= 8'b11011111; // 3211 : 223 - 0xdf
      12'hC8C: dout <= 8'b11011111; // 3212 : 223 - 0xdf
      12'hC8D: dout <= 8'b11001111; // 3213 : 207 - 0xcf
      12'hC8E: dout <= 8'b11101111; // 3214 : 239 - 0xef
      12'hC8F: dout <= 8'b11100111; // 3215 : 231 - 0xe7
      12'hC90: dout <= 8'b11110011; // 3216 : 243 - 0xf3 -- Background 0x92
      12'hC91: dout <= 8'b11111001; // 3217 : 249 - 0xf9
      12'hC92: dout <= 8'b11111100; // 3218 : 252 - 0xfc
      12'hC93: dout <= 8'b11111100; // 3219 : 252 - 0xfc
      12'hC94: dout <= 8'b11111100; // 3220 : 252 - 0xfc
      12'hC95: dout <= 8'b11110000; // 3221 : 240 - 0xf0
      12'hC96: dout <= 8'b11000000; // 3222 : 192 - 0xc0
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b00000011; // 3224 :   3 - 0x3 -- Background 0x93
      12'hC99: dout <= 8'b00001111; // 3225 :  15 - 0xf
      12'hC9A: dout <= 8'b00111111; // 3226 :  63 - 0x3f
      12'hC9B: dout <= 8'b00001111; // 3227 :  15 - 0xf
      12'hC9C: dout <= 8'b00001111; // 3228 :  15 - 0xf
      12'hC9D: dout <= 8'b00011001; // 3229 :  25 - 0x19
      12'hC9E: dout <= 8'b00010000; // 3230 :  16 - 0x10
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00011111; // 3232 :  31 - 0x1f -- Background 0x94
      12'hCA1: dout <= 8'b01111111; // 3233 : 127 - 0x7f
      12'hCA2: dout <= 8'b11111110; // 3234 : 254 - 0xfe
      12'hCA3: dout <= 8'b11111000; // 3235 : 248 - 0xf8
      12'hCA4: dout <= 8'b11110000; // 3236 : 240 - 0xf0
      12'hCA5: dout <= 8'b10011000; // 3237 : 152 - 0x98
      12'hCA6: dout <= 8'b00001100; // 3238 :  12 - 0xc
      12'hCA7: dout <= 8'b00001110; // 3239 :  14 - 0xe
      12'hCA8: dout <= 8'b11011111; // 3240 : 223 - 0xdf -- Background 0x95
      12'hCA9: dout <= 8'b11001110; // 3241 : 206 - 0xce
      12'hCAA: dout <= 8'b11100100; // 3242 : 228 - 0xe4
      12'hCAB: dout <= 8'b11110000; // 3243 : 240 - 0xf0
      12'hCAC: dout <= 8'b11111000; // 3244 : 248 - 0xf8
      12'hCAD: dout <= 8'b11111000; // 3245 : 248 - 0xf8
      12'hCAE: dout <= 8'b11111100; // 3246 : 252 - 0xfc
      12'hCAF: dout <= 8'b11111110; // 3247 : 254 - 0xfe
      12'hCB0: dout <= 8'b11111111; // 3248 : 255 - 0xff -- Background 0x96
      12'hCB1: dout <= 8'b11111111; // 3249 : 255 - 0xff
      12'hCB2: dout <= 8'b11111111; // 3250 : 255 - 0xff
      12'hCB3: dout <= 8'b11111111; // 3251 : 255 - 0xff
      12'hCB4: dout <= 8'b01111111; // 3252 : 127 - 0x7f
      12'hCB5: dout <= 8'b10111111; // 3253 : 191 - 0xbf
      12'hCB6: dout <= 8'b00011111; // 3254 :  31 - 0x1f
      12'hCB7: dout <= 8'b01101111; // 3255 : 111 - 0x6f
      12'hCB8: dout <= 8'b11110111; // 3256 : 247 - 0xf7 -- Background 0x97
      12'hCB9: dout <= 8'b11110011; // 3257 : 243 - 0xf3
      12'hCBA: dout <= 8'b11111001; // 3258 : 249 - 0xf9
      12'hCBB: dout <= 8'b11111000; // 3259 : 248 - 0xf8
      12'hCBC: dout <= 8'b11110000; // 3260 : 240 - 0xf0
      12'hCBD: dout <= 8'b10110100; // 3261 : 180 - 0xb4
      12'hCBE: dout <= 8'b00001010; // 3262 :  10 - 0xa
      12'hCBF: dout <= 8'b00000010; // 3263 :   2 - 0x2
      12'hCC0: dout <= 8'b10000000; // 3264 : 128 - 0x80 -- Background 0x98
      12'hCC1: dout <= 8'b11000000; // 3265 : 192 - 0xc0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b11000000; // 3268 : 192 - 0xc0
      12'hCC5: dout <= 8'b10011000; // 3269 : 152 - 0x98
      12'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- Background 0x99
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00111110; // 3274 :  62 - 0x3e
      12'hCCB: dout <= 8'b01000000; // 3275 :  64 - 0x40
      12'hCCC: dout <= 8'b10000000; // 3276 : 128 - 0x80
      12'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Background 0x9a
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b10000000; // 3282 : 128 - 0x80
      12'hCD3: dout <= 8'b10000000; // 3283 : 128 - 0x80
      12'hCD4: dout <= 8'b11000000; // 3284 : 192 - 0xc0
      12'hCD5: dout <= 8'b11100000; // 3285 : 224 - 0xe0
      12'hCD6: dout <= 8'b11100000; // 3286 : 224 - 0xe0
      12'hCD7: dout <= 8'b11110000; // 3287 : 240 - 0xf0
      12'hCD8: dout <= 8'b11110000; // 3288 : 240 - 0xf0 -- Background 0x9b
      12'hCD9: dout <= 8'b11100000; // 3289 : 224 - 0xe0
      12'hCDA: dout <= 8'b11110000; // 3290 : 240 - 0xf0
      12'hCDB: dout <= 8'b11100000; // 3291 : 224 - 0xe0
      12'hCDC: dout <= 8'b10000000; // 3292 : 128 - 0x80
      12'hCDD: dout <= 8'b00001000; // 3293 :   8 - 0x8
      12'hCDE: dout <= 8'b00000100; // 3294 :   4 - 0x4
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Background 0x9c
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000001; // 3298 :   1 - 0x1
      12'hCE3: dout <= 8'b00000011; // 3299 :   3 - 0x3
      12'hCE4: dout <= 8'b00000011; // 3300 :   3 - 0x3
      12'hCE5: dout <= 8'b00000011; // 3301 :   3 - 0x3
      12'hCE6: dout <= 8'b00000111; // 3302 :   7 - 0x7
      12'hCE7: dout <= 8'b00000111; // 3303 :   7 - 0x7
      12'hCE8: dout <= 8'b00000111; // 3304 :   7 - 0x7 -- Background 0x9d
      12'hCE9: dout <= 8'b00000011; // 3305 :   3 - 0x3
      12'hCEA: dout <= 8'b00000011; // 3306 :   3 - 0x3
      12'hCEB: dout <= 8'b00000011; // 3307 :   3 - 0x3
      12'hCEC: dout <= 8'b00000011; // 3308 :   3 - 0x3
      12'hCED: dout <= 8'b00000011; // 3309 :   3 - 0x3
      12'hCEE: dout <= 8'b00000011; // 3310 :   3 - 0x3
      12'hCEF: dout <= 8'b00000001; // 3311 :   1 - 0x1
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Background 0x9e
      12'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      12'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      12'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      12'hCF5: dout <= 8'b00000001; // 3317 :   1 - 0x1
      12'hCF6: dout <= 8'b00000010; // 3318 :   2 - 0x2
      12'hCF7: dout <= 8'b00000100; // 3319 :   4 - 0x4
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- Background 0x9f
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout <= 8'b00011100; // 3326 :  28 - 0x1c
      12'hCFF: dout <= 8'b00111011; // 3327 :  59 - 0x3b
      12'hD00: dout <= 8'b01111110; // 3328 : 126 - 0x7e -- Background 0xa0
      12'hD01: dout <= 8'b11111110; // 3329 : 254 - 0xfe
      12'hD02: dout <= 8'b11111111; // 3330 : 255 - 0xff
      12'hD03: dout <= 8'b11111111; // 3331 : 255 - 0xff
      12'hD04: dout <= 8'b11111111; // 3332 : 255 - 0xff
      12'hD05: dout <= 8'b11111111; // 3333 : 255 - 0xff
      12'hD06: dout <= 8'b11111101; // 3334 : 253 - 0xfd
      12'hD07: dout <= 8'b11111001; // 3335 : 249 - 0xf9
      12'hD08: dout <= 8'b11110011; // 3336 : 243 - 0xf3 -- Background 0xa1
      12'hD09: dout <= 8'b11110111; // 3337 : 247 - 0xf7
      12'hD0A: dout <= 8'b11110110; // 3338 : 246 - 0xf6
      12'hD0B: dout <= 8'b11101110; // 3339 : 238 - 0xee
      12'hD0C: dout <= 8'b11111101; // 3340 : 253 - 0xfd
      12'hD0D: dout <= 8'b11111100; // 3341 : 252 - 0xfc
      12'hD0E: dout <= 8'b11111000; // 3342 : 248 - 0xf8
      12'hD0F: dout <= 8'b11100001; // 3343 : 225 - 0xe1
      12'hD10: dout <= 8'b11010011; // 3344 : 211 - 0xd3 -- Background 0xa2
      12'hD11: dout <= 8'b11001011; // 3345 : 203 - 0xcb
      12'hD12: dout <= 8'b11000011; // 3346 : 195 - 0xc3
      12'hD13: dout <= 8'b11100001; // 3347 : 225 - 0xe1
      12'hD14: dout <= 8'b11111001; // 3348 : 249 - 0xf9
      12'hD15: dout <= 8'b00111001; // 3349 :  57 - 0x39
      12'hD16: dout <= 8'b01000010; // 3350 :  66 - 0x42
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000111; // 3352 :   7 - 0x7 -- Background 0xa3
      12'hD19: dout <= 8'b00001111; // 3353 :  15 - 0xf
      12'hD1A: dout <= 8'b00011001; // 3354 :  25 - 0x19
      12'hD1B: dout <= 8'b00110000; // 3355 :  48 - 0x30
      12'hD1C: dout <= 8'b01100011; // 3356 :  99 - 0x63
      12'hD1D: dout <= 8'b01110010; // 3357 : 114 - 0x72
      12'hD1E: dout <= 8'b01110000; // 3358 : 112 - 0x70
      12'hD1F: dout <= 8'b00000001; // 3359 :   1 - 0x1
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout <= 8'b00011111; // 3361 :  31 - 0x1f
      12'hD22: dout <= 8'b00100000; // 3362 :  32 - 0x20
      12'hD23: dout <= 8'b11000000; // 3363 : 192 - 0xc0
      12'hD24: dout <= 8'b11000000; // 3364 : 192 - 0xc0
      12'hD25: dout <= 8'b11110000; // 3365 : 240 - 0xf0
      12'hD26: dout <= 8'b11111111; // 3366 : 255 - 0xff
      12'hD27: dout <= 8'b11111111; // 3367 : 255 - 0xff
      12'hD28: dout <= 8'b10101011; // 3368 : 171 - 0xab -- Background 0xa5
      12'hD29: dout <= 8'b11000001; // 3369 : 193 - 0xc1
      12'hD2A: dout <= 8'b10000001; // 3370 : 129 - 0x81
      12'hD2B: dout <= 8'b10010001; // 3371 : 145 - 0x91
      12'hD2C: dout <= 8'b10000010; // 3372 : 130 - 0x82
      12'hD2D: dout <= 8'b11111100; // 3373 : 252 - 0xfc
      12'hD2E: dout <= 8'b11100000; // 3374 : 224 - 0xe0
      12'hD2F: dout <= 8'b11001110; // 3375 : 206 - 0xce
      12'hD30: dout <= 8'b11100101; // 3376 : 229 - 0xe5 -- Background 0xa6
      12'hD31: dout <= 8'b11011010; // 3377 : 218 - 0xda
      12'hD32: dout <= 8'b11110000; // 3378 : 240 - 0xf0
      12'hD33: dout <= 8'b11100000; // 3379 : 224 - 0xe0
      12'hD34: dout <= 8'b11000000; // 3380 : 192 - 0xc0
      12'hD35: dout <= 8'b00000000; // 3381 :   0 - 0x0
      12'hD36: dout <= 8'b00000000; // 3382 :   0 - 0x0
      12'hD37: dout <= 8'b00000000; // 3383 :   0 - 0x0
      12'hD38: dout <= 8'b11110000; // 3384 : 240 - 0xf0 -- Background 0xa7
      12'hD39: dout <= 8'b11111000; // 3385 : 248 - 0xf8
      12'hD3A: dout <= 8'b11001100; // 3386 : 204 - 0xcc
      12'hD3B: dout <= 8'b10000110; // 3387 : 134 - 0x86
      12'hD3C: dout <= 8'b01100010; // 3388 :  98 - 0x62
      12'hD3D: dout <= 8'b00100110; // 3389 :  38 - 0x26
      12'hD3E: dout <= 8'b00000110; // 3390 :   6 - 0x6
      12'hD3F: dout <= 8'b11000000; // 3391 : 192 - 0xc0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xa8
      12'hD41: dout <= 8'b11111100; // 3393 : 252 - 0xfc
      12'hD42: dout <= 8'b00000110; // 3394 :   6 - 0x6
      12'hD43: dout <= 8'b00000011; // 3395 :   3 - 0x3
      12'hD44: dout <= 8'b00000001; // 3396 :   1 - 0x1
      12'hD45: dout <= 8'b00000111; // 3397 :   7 - 0x7
      12'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      12'hD47: dout <= 8'b11111111; // 3399 : 255 - 0xff
      12'hD48: dout <= 8'b11010101; // 3400 : 213 - 0xd5 -- Background 0xa9
      12'hD49: dout <= 8'b10000011; // 3401 : 131 - 0x83
      12'hD4A: dout <= 8'b10000001; // 3402 : 129 - 0x81
      12'hD4B: dout <= 8'b10001001; // 3403 : 137 - 0x89
      12'hD4C: dout <= 8'b01000001; // 3404 :  65 - 0x41
      12'hD4D: dout <= 8'b00111111; // 3405 :  63 - 0x3f
      12'hD4E: dout <= 8'b00000111; // 3406 :   7 - 0x7
      12'hD4F: dout <= 8'b11010011; // 3407 : 211 - 0xd3
      12'hD50: dout <= 8'b01101111; // 3408 : 111 - 0x6f -- Background 0xaa
      12'hD51: dout <= 8'b11011011; // 3409 : 219 - 0xdb
      12'hD52: dout <= 8'b00001111; // 3410 :  15 - 0xf
      12'hD53: dout <= 8'b00000111; // 3411 :   7 - 0x7
      12'hD54: dout <= 8'b00000011; // 3412 :   3 - 0x3
      12'hD55: dout <= 8'b00000000; // 3413 :   0 - 0x0
      12'hD56: dout <= 8'b00000000; // 3414 :   0 - 0x0
      12'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- Background 0xab
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout <= 8'b00000000; // 3419 :   0 - 0x0
      12'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout <= 8'b00111000; // 3422 :  56 - 0x38
      12'hD5F: dout <= 8'b11011100; // 3423 : 220 - 0xdc
      12'hD60: dout <= 8'b01111110; // 3424 : 126 - 0x7e -- Background 0xac
      12'hD61: dout <= 8'b01111111; // 3425 : 127 - 0x7f
      12'hD62: dout <= 8'b01111111; // 3426 : 127 - 0x7f
      12'hD63: dout <= 8'b11111111; // 3427 : 255 - 0xff
      12'hD64: dout <= 8'b11111111; // 3428 : 255 - 0xff
      12'hD65: dout <= 8'b11111111; // 3429 : 255 - 0xff
      12'hD66: dout <= 8'b10111111; // 3430 : 191 - 0xbf
      12'hD67: dout <= 8'b10011111; // 3431 : 159 - 0x9f
      12'hD68: dout <= 8'b11001111; // 3432 : 207 - 0xcf -- Background 0xad
      12'hD69: dout <= 8'b11101111; // 3433 : 239 - 0xef
      12'hD6A: dout <= 8'b01101111; // 3434 : 111 - 0x6f
      12'hD6B: dout <= 8'b01110111; // 3435 : 119 - 0x77
      12'hD6C: dout <= 8'b10111111; // 3436 : 191 - 0xbf
      12'hD6D: dout <= 8'b00111111; // 3437 :  63 - 0x3f
      12'hD6E: dout <= 8'b00011111; // 3438 :  31 - 0x1f
      12'hD6F: dout <= 8'b10000111; // 3439 : 135 - 0x87
      12'hD70: dout <= 8'b11001011; // 3440 : 203 - 0xcb -- Background 0xae
      12'hD71: dout <= 8'b11010011; // 3441 : 211 - 0xd3
      12'hD72: dout <= 8'b11000011; // 3442 : 195 - 0xc3
      12'hD73: dout <= 8'b10000111; // 3443 : 135 - 0x87
      12'hD74: dout <= 8'b10011111; // 3444 : 159 - 0x9f
      12'hD75: dout <= 8'b10011100; // 3445 : 156 - 0x9c
      12'hD76: dout <= 8'b01000010; // 3446 :  66 - 0x42
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0 -- Background 0xaf
      12'hD79: dout <= 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout <= 8'b10000000; // 3450 : 128 - 0x80
      12'hD7B: dout <= 8'b11000000; // 3451 : 192 - 0xc0
      12'hD7C: dout <= 8'b11000000; // 3452 : 192 - 0xc0
      12'hD7D: dout <= 8'b11000000; // 3453 : 192 - 0xc0
      12'hD7E: dout <= 8'b11100000; // 3454 : 224 - 0xe0
      12'hD7F: dout <= 8'b11100000; // 3455 : 224 - 0xe0
      12'hD80: dout <= 8'b11100000; // 3456 : 224 - 0xe0 -- Background 0xb0
      12'hD81: dout <= 8'b11000000; // 3457 : 192 - 0xc0
      12'hD82: dout <= 8'b11000000; // 3458 : 192 - 0xc0
      12'hD83: dout <= 8'b11000000; // 3459 : 192 - 0xc0
      12'hD84: dout <= 8'b11000000; // 3460 : 192 - 0xc0
      12'hD85: dout <= 8'b11000000; // 3461 : 192 - 0xc0
      12'hD86: dout <= 8'b11000000; // 3462 : 192 - 0xc0
      12'hD87: dout <= 8'b10000000; // 3463 : 128 - 0x80
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- Background 0xb1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b00000000; // 3466 :   0 - 0x0
      12'hD8B: dout <= 8'b00000000; // 3467 :   0 - 0x0
      12'hD8C: dout <= 8'b00000000; // 3468 :   0 - 0x0
      12'hD8D: dout <= 8'b10000000; // 3469 : 128 - 0x80
      12'hD8E: dout <= 8'b01000000; // 3470 :  64 - 0x40
      12'hD8F: dout <= 8'b00100000; // 3471 :  32 - 0x20
      12'hD90: dout <= 8'b00000000; // 3472 :   0 - 0x0 -- Background 0xb2
      12'hD91: dout <= 8'b00000000; // 3473 :   0 - 0x0
      12'hD92: dout <= 8'b00000000; // 3474 :   0 - 0x0
      12'hD93: dout <= 8'b00000001; // 3475 :   1 - 0x1
      12'hD94: dout <= 8'b00000011; // 3476 :   3 - 0x3
      12'hD95: dout <= 8'b00000111; // 3477 :   7 - 0x7
      12'hD96: dout <= 8'b00000111; // 3478 :   7 - 0x7
      12'hD97: dout <= 8'b00000111; // 3479 :   7 - 0x7
      12'hD98: dout <= 8'b00000011; // 3480 :   3 - 0x3 -- Background 0xb3
      12'hD99: dout <= 8'b00000001; // 3481 :   1 - 0x1
      12'hD9A: dout <= 8'b00000000; // 3482 :   0 - 0x0
      12'hD9B: dout <= 8'b00000000; // 3483 :   0 - 0x0
      12'hD9C: dout <= 8'b00000000; // 3484 :   0 - 0x0
      12'hD9D: dout <= 8'b00000000; // 3485 :   0 - 0x0
      12'hD9E: dout <= 8'b00000001; // 3486 :   1 - 0x1
      12'hD9F: dout <= 8'b00000001; // 3487 :   1 - 0x1
      12'hDA0: dout <= 8'b00000001; // 3488 :   1 - 0x1 -- Background 0xb4
      12'hDA1: dout <= 8'b00000001; // 3489 :   1 - 0x1
      12'hDA2: dout <= 8'b00000111; // 3490 :   7 - 0x7
      12'hDA3: dout <= 8'b00000011; // 3491 :   3 - 0x3
      12'hDA4: dout <= 8'b00000100; // 3492 :   4 - 0x4
      12'hDA5: dout <= 8'b00000000; // 3493 :   0 - 0x0
      12'hDA6: dout <= 8'b00000000; // 3494 :   0 - 0x0
      12'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- Background 0xb5
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b00000000; // 3499 :   0 - 0x0
      12'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      12'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      12'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout <= 8'b00000111; // 3503 :   7 - 0x7
      12'hDB0: dout <= 8'b00001110; // 3504 :  14 - 0xe -- Background 0xb6
      12'hDB1: dout <= 8'b00111110; // 3505 :  62 - 0x3e
      12'hDB2: dout <= 8'b01111111; // 3506 : 127 - 0x7f
      12'hDB3: dout <= 8'b11111111; // 3507 : 255 - 0xff
      12'hDB4: dout <= 8'b11111111; // 3508 : 255 - 0xff
      12'hDB5: dout <= 8'b11101111; // 3509 : 239 - 0xef
      12'hDB6: dout <= 8'b11110111; // 3510 : 247 - 0xf7
      12'hDB7: dout <= 8'b11111000; // 3511 : 248 - 0xf8
      12'hDB8: dout <= 8'b11111111; // 3512 : 255 - 0xff -- Background 0xb7
      12'hDB9: dout <= 8'b11111111; // 3513 : 255 - 0xff
      12'hDBA: dout <= 8'b11111111; // 3514 : 255 - 0xff
      12'hDBB: dout <= 8'b00011111; // 3515 :  31 - 0x1f
      12'hDBC: dout <= 8'b00011111; // 3516 :  31 - 0x1f
      12'hDBD: dout <= 8'b01111111; // 3517 : 127 - 0x7f
      12'hDBE: dout <= 8'b11111111; // 3518 : 255 - 0xff
      12'hDBF: dout <= 8'b11111110; // 3519 : 254 - 0xfe
      12'hDC0: dout <= 8'b11111111; // 3520 : 255 - 0xff -- Background 0xb8
      12'hDC1: dout <= 8'b11111111; // 3521 : 255 - 0xff
      12'hDC2: dout <= 8'b11111111; // 3522 : 255 - 0xff
      12'hDC3: dout <= 8'b11111100; // 3523 : 252 - 0xfc
      12'hDC4: dout <= 8'b11111000; // 3524 : 248 - 0xf8
      12'hDC5: dout <= 8'b10000000; // 3525 : 128 - 0x80
      12'hDC6: dout <= 8'b00000000; // 3526 :   0 - 0x0
      12'hDC7: dout <= 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout <= 8'b00110000; // 3528 :  48 - 0x30 -- Background 0xb9
      12'hDC9: dout <= 8'b01111111; // 3529 : 127 - 0x7f
      12'hDCA: dout <= 8'b01111111; // 3530 : 127 - 0x7f
      12'hDCB: dout <= 8'b00111111; // 3531 :  63 - 0x3f
      12'hDCC: dout <= 8'b10000111; // 3532 : 135 - 0x87
      12'hDCD: dout <= 8'b11110000; // 3533 : 240 - 0xf0
      12'hDCE: dout <= 8'b11111111; // 3534 : 255 - 0xff
      12'hDCF: dout <= 8'b11111111; // 3535 : 255 - 0xff
      12'hDD0: dout <= 8'b11100101; // 3536 : 229 - 0xe5 -- Background 0xba
      12'hDD1: dout <= 8'b11011010; // 3537 : 218 - 0xda
      12'hDD2: dout <= 8'b11000000; // 3538 : 192 - 0xc0
      12'hDD3: dout <= 8'b00000000; // 3539 :   0 - 0x0
      12'hDD4: dout <= 8'b00000000; // 3540 :   0 - 0x0
      12'hDD5: dout <= 8'b00000000; // 3541 :   0 - 0x0
      12'hDD6: dout <= 8'b00000000; // 3542 :   0 - 0x0
      12'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout <= 8'b00000110; // 3544 :   6 - 0x6 -- Background 0xbb
      12'hDD9: dout <= 8'b11111111; // 3545 : 255 - 0xff
      12'hDDA: dout <= 8'b11111111; // 3546 : 255 - 0xff
      12'hDDB: dout <= 8'b11111110; // 3547 : 254 - 0xfe
      12'hDDC: dout <= 8'b11110001; // 3548 : 241 - 0xf1
      12'hDDD: dout <= 8'b00000111; // 3549 :   7 - 0x7
      12'hDDE: dout <= 8'b11111111; // 3550 : 255 - 0xff
      12'hDDF: dout <= 8'b11111111; // 3551 : 255 - 0xff
      12'hDE0: dout <= 8'b00000000; // 3552 :   0 - 0x0 -- Background 0xbc
      12'hDE1: dout <= 8'b00000001; // 3553 :   1 - 0x1
      12'hDE2: dout <= 8'b00000010; // 3554 :   2 - 0x2
      12'hDE3: dout <= 8'b00000111; // 3555 :   7 - 0x7
      12'hDE4: dout <= 8'b00000000; // 3556 :   0 - 0x0
      12'hDE5: dout <= 8'b00000000; // 3557 :   0 - 0x0
      12'hDE6: dout <= 8'b00100000; // 3558 :  32 - 0x20
      12'hDE7: dout <= 8'b11111111; // 3559 : 255 - 0xff
      12'hDE8: dout <= 8'b01111111; // 3560 : 127 - 0x7f -- Background 0xbd
      12'hDE9: dout <= 8'b01111111; // 3561 : 127 - 0x7f
      12'hDEA: dout <= 8'b01111111; // 3562 : 127 - 0x7f
      12'hDEB: dout <= 8'b11111111; // 3563 : 255 - 0xff
      12'hDEC: dout <= 8'b11111111; // 3564 : 255 - 0xff
      12'hDED: dout <= 8'b11111111; // 3565 : 255 - 0xff
      12'hDEE: dout <= 8'b11111111; // 3566 : 255 - 0xff
      12'hDEF: dout <= 8'b11111110; // 3567 : 254 - 0xfe
      12'hDF0: dout <= 8'b11111100; // 3568 : 252 - 0xfc -- Background 0xbe
      12'hDF1: dout <= 8'b10111000; // 3569 : 184 - 0xb8
      12'hDF2: dout <= 8'b01111000; // 3570 : 120 - 0x78
      12'hDF3: dout <= 8'b01111000; // 3571 : 120 - 0x78
      12'hDF4: dout <= 8'b10110000; // 3572 : 176 - 0xb0
      12'hDF5: dout <= 8'b01111000; // 3573 : 120 - 0x78
      12'hDF6: dout <= 8'b11111100; // 3574 : 252 - 0xfc
      12'hDF7: dout <= 8'b11111110; // 3575 : 254 - 0xfe
      12'hDF8: dout <= 8'b11111111; // 3576 : 255 - 0xff -- Background 0xbf
      12'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      12'hDFA: dout <= 8'b11111111; // 3578 : 255 - 0xff
      12'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout <= 8'b11111111; // 3580 : 255 - 0xff
      12'hDFD: dout <= 8'b10011100; // 3581 : 156 - 0x9c
      12'hDFE: dout <= 8'b01000010; // 3582 :  66 - 0x42
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout <= 8'b00100000; // 3586 :  32 - 0x20
      12'hE03: dout <= 8'b01000000; // 3587 :  64 - 0x40
      12'hE04: dout <= 8'b10001010; // 3588 : 138 - 0x8a
      12'hE05: dout <= 8'b00011110; // 3589 :  30 - 0x1e
      12'hE06: dout <= 8'b01111110; // 3590 : 126 - 0x7e
      12'hE07: dout <= 8'b10111110; // 3591 : 190 - 0xbe
      12'hE08: dout <= 8'b11011111; // 3592 : 223 - 0xdf -- Background 0xc1
      12'hE09: dout <= 8'b11111111; // 3593 : 255 - 0xff
      12'hE0A: dout <= 8'b11111110; // 3594 : 254 - 0xfe
      12'hE0B: dout <= 8'b11111100; // 3595 : 252 - 0xfc
      12'hE0C: dout <= 8'b11110000; // 3596 : 240 - 0xf0
      12'hE0D: dout <= 8'b11100000; // 3597 : 224 - 0xe0
      12'hE0E: dout <= 8'b10000000; // 3598 : 128 - 0x80
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout <= 8'b00000100; // 3602 :   4 - 0x4
      12'hE13: dout <= 8'b00000010; // 3603 :   2 - 0x2
      12'hE14: dout <= 8'b01010001; // 3604 :  81 - 0x51
      12'hE15: dout <= 8'b01111000; // 3605 : 120 - 0x78
      12'hE16: dout <= 8'b01111110; // 3606 : 126 - 0x7e
      12'hE17: dout <= 8'b11111101; // 3607 : 253 - 0xfd
      12'hE18: dout <= 8'b11111011; // 3608 : 251 - 0xfb -- Background 0xc3
      12'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout <= 8'b01111111; // 3610 : 127 - 0x7f
      12'hE1B: dout <= 8'b00111111; // 3611 :  63 - 0x3f
      12'hE1C: dout <= 8'b00001111; // 3612 :  15 - 0xf
      12'hE1D: dout <= 8'b00000111; // 3613 :   7 - 0x7
      12'hE1E: dout <= 8'b00000001; // 3614 :   1 - 0x1
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout <= 8'b10000000; // 3617 : 128 - 0x80
      12'hE22: dout <= 8'b01000000; // 3618 :  64 - 0x40
      12'hE23: dout <= 8'b11100000; // 3619 : 224 - 0xe0
      12'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout <= 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout <= 8'b00000100; // 3622 :   4 - 0x4
      12'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout <= 8'b11111110; // 3624 : 254 - 0xfe -- Background 0xc5
      12'hE29: dout <= 8'b11111110; // 3625 : 254 - 0xfe
      12'hE2A: dout <= 8'b11111110; // 3626 : 254 - 0xfe
      12'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout <= 8'b11111111; // 3628 : 255 - 0xff
      12'hE2D: dout <= 8'b11111111; // 3629 : 255 - 0xff
      12'hE2E: dout <= 8'b11111111; // 3630 : 255 - 0xff
      12'hE2F: dout <= 8'b01111111; // 3631 : 127 - 0x7f
      12'hE30: dout <= 8'b00111111; // 3632 :  63 - 0x3f -- Background 0xc6
      12'hE31: dout <= 8'b00011101; // 3633 :  29 - 0x1d
      12'hE32: dout <= 8'b00011110; // 3634 :  30 - 0x1e
      12'hE33: dout <= 8'b00011110; // 3635 :  30 - 0x1e
      12'hE34: dout <= 8'b00001101; // 3636 :  13 - 0xd
      12'hE35: dout <= 8'b00011110; // 3637 :  30 - 0x1e
      12'hE36: dout <= 8'b00111111; // 3638 :  63 - 0x3f
      12'hE37: dout <= 8'b01111111; // 3639 : 127 - 0x7f
      12'hE38: dout <= 8'b11111111; // 3640 : 255 - 0xff -- Background 0xc7
      12'hE39: dout <= 8'b11111111; // 3641 : 255 - 0xff
      12'hE3A: dout <= 8'b11111111; // 3642 : 255 - 0xff
      12'hE3B: dout <= 8'b11111111; // 3643 : 255 - 0xff
      12'hE3C: dout <= 8'b11111111; // 3644 : 255 - 0xff
      12'hE3D: dout <= 8'b00111001; // 3645 :  57 - 0x39
      12'hE3E: dout <= 8'b01000010; // 3646 :  66 - 0x42
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b01101111; // 3648 : 111 - 0x6f -- Background 0xc8
      12'hE41: dout <= 8'b11011011; // 3649 : 219 - 0xdb
      12'hE42: dout <= 8'b00000011; // 3650 :   3 - 0x3
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout <= 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- Background 0xc9
      12'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      12'hE4C: dout <= 8'b00000000; // 3660 :   0 - 0x0
      12'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b11100000; // 3663 : 224 - 0xe0
      12'hE50: dout <= 8'b01110000; // 3664 : 112 - 0x70 -- Background 0xca
      12'hE51: dout <= 8'b01111100; // 3665 : 124 - 0x7c
      12'hE52: dout <= 8'b01111110; // 3666 : 126 - 0x7e
      12'hE53: dout <= 8'b11111111; // 3667 : 255 - 0xff
      12'hE54: dout <= 8'b11111111; // 3668 : 255 - 0xff
      12'hE55: dout <= 8'b11110111; // 3669 : 247 - 0xf7
      12'hE56: dout <= 8'b11101111; // 3670 : 239 - 0xef
      12'hE57: dout <= 8'b00011111; // 3671 :  31 - 0x1f
      12'hE58: dout <= 8'b11111111; // 3672 : 255 - 0xff -- Background 0xcb
      12'hE59: dout <= 8'b11111111; // 3673 : 255 - 0xff
      12'hE5A: dout <= 8'b11111111; // 3674 : 255 - 0xff
      12'hE5B: dout <= 8'b11111000; // 3675 : 248 - 0xf8
      12'hE5C: dout <= 8'b11111000; // 3676 : 248 - 0xf8
      12'hE5D: dout <= 8'b11111110; // 3677 : 254 - 0xfe
      12'hE5E: dout <= 8'b11111111; // 3678 : 255 - 0xff
      12'hE5F: dout <= 8'b11111111; // 3679 : 255 - 0xff
      12'hE60: dout <= 8'b11111111; // 3680 : 255 - 0xff -- Background 0xcc
      12'hE61: dout <= 8'b11111111; // 3681 : 255 - 0xff
      12'hE62: dout <= 8'b11111111; // 3682 : 255 - 0xff
      12'hE63: dout <= 8'b00111111; // 3683 :  63 - 0x3f
      12'hE64: dout <= 8'b00011110; // 3684 :  30 - 0x1e
      12'hE65: dout <= 8'b00000001; // 3685 :   1 - 0x1
      12'hE66: dout <= 8'b00000000; // 3686 :   0 - 0x0
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b10000000; // 3691 : 128 - 0x80
      12'hE6C: dout <= 8'b11000000; // 3692 : 192 - 0xc0
      12'hE6D: dout <= 8'b11100000; // 3693 : 224 - 0xe0
      12'hE6E: dout <= 8'b11100000; // 3694 : 224 - 0xe0
      12'hE6F: dout <= 8'b11100000; // 3695 : 224 - 0xe0
      12'hE70: dout <= 8'b11000000; // 3696 : 192 - 0xc0 -- Background 0xce
      12'hE71: dout <= 8'b10000000; // 3697 : 128 - 0x80
      12'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout <= 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout <= 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout <= 8'b10000000; // 3702 : 128 - 0x80
      12'hE77: dout <= 8'b10000000; // 3703 : 128 - 0x80
      12'hE78: dout <= 8'b10000000; // 3704 : 128 - 0x80 -- Background 0xcf
      12'hE79: dout <= 8'b10000000; // 3705 : 128 - 0x80
      12'hE7A: dout <= 8'b11100000; // 3706 : 224 - 0xe0
      12'hE7B: dout <= 8'b11000000; // 3707 : 192 - 0xc0
      12'hE7C: dout <= 8'b00100000; // 3708 :  32 - 0x20
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b00011111; // 3712 :  31 - 0x1f -- Background 0xd0
      12'hE81: dout <= 8'b00000110; // 3713 :   6 - 0x6
      12'hE82: dout <= 8'b00000110; // 3714 :   6 - 0x6
      12'hE83: dout <= 8'b00000110; // 3715 :   6 - 0x6
      12'hE84: dout <= 8'b00000110; // 3716 :   6 - 0x6
      12'hE85: dout <= 8'b00000110; // 3717 :   6 - 0x6
      12'hE86: dout <= 8'b00000110; // 3718 :   6 - 0x6
      12'hE87: dout <= 8'b00000000; // 3719 :   0 - 0x0
      12'hE88: dout <= 8'b00111001; // 3720 :  57 - 0x39 -- Background 0xd1
      12'hE89: dout <= 8'b01100101; // 3721 : 101 - 0x65
      12'hE8A: dout <= 8'b01100101; // 3722 : 101 - 0x65
      12'hE8B: dout <= 8'b01100101; // 3723 : 101 - 0x65
      12'hE8C: dout <= 8'b01100101; // 3724 : 101 - 0x65
      12'hE8D: dout <= 8'b01100101; // 3725 : 101 - 0x65
      12'hE8E: dout <= 8'b00111001; // 3726 :  57 - 0x39
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b11100000; // 3728 : 224 - 0xe0 -- Background 0xd2
      12'hE91: dout <= 8'b10110000; // 3729 : 176 - 0xb0
      12'hE92: dout <= 8'b10110000; // 3730 : 176 - 0xb0
      12'hE93: dout <= 8'b10110110; // 3731 : 182 - 0xb6
      12'hE94: dout <= 8'b11100110; // 3732 : 230 - 0xe6
      12'hE95: dout <= 8'b10000000; // 3733 : 128 - 0x80
      12'hE96: dout <= 8'b10000000; // 3734 : 128 - 0x80
      12'hE97: dout <= 8'b00000000; // 3735 :   0 - 0x0
      12'hE98: dout <= 8'b00111100; // 3736 :  60 - 0x3c -- Background 0xd3
      12'hE99: dout <= 8'b01000010; // 3737 :  66 - 0x42
      12'hE9A: dout <= 8'b10011001; // 3738 : 153 - 0x99
      12'hE9B: dout <= 8'b10100001; // 3739 : 161 - 0xa1
      12'hE9C: dout <= 8'b10100001; // 3740 : 161 - 0xa1
      12'hE9D: dout <= 8'b10011001; // 3741 : 153 - 0x99
      12'hE9E: dout <= 8'b01000010; // 3742 :  66 - 0x42
      12'hE9F: dout <= 8'b00111100; // 3743 :  60 - 0x3c
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout <= 8'b00000011; // 3747 :   3 - 0x3
      12'hEA4: dout <= 8'b00000110; // 3748 :   6 - 0x6
      12'hEA5: dout <= 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout <= 8'b00000001; // 3750 :   1 - 0x1
      12'hEA7: dout <= 8'b00000111; // 3751 :   7 - 0x7
      12'hEA8: dout <= 8'b00001111; // 3752 :  15 - 0xf -- Background 0xd5
      12'hEA9: dout <= 8'b00011111; // 3753 :  31 - 0x1f
      12'hEAA: dout <= 8'b00111111; // 3754 :  63 - 0x3f
      12'hEAB: dout <= 8'b01111111; // 3755 : 127 - 0x7f
      12'hEAC: dout <= 8'b01111111; // 3756 : 127 - 0x7f
      12'hEAD: dout <= 8'b01111111; // 3757 : 127 - 0x7f
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b01111111; // 3759 : 127 - 0x7f
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout <= 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout <= 8'b00000000; // 3762 :   0 - 0x0
      12'hEB3: dout <= 8'b10000000; // 3763 : 128 - 0x80
      12'hEB4: dout <= 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout <= 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout <= 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout <= 8'b10100000; // 3767 : 160 - 0xa0
      12'hEB8: dout <= 8'b11100000; // 3768 : 224 - 0xe0 -- Background 0xd7
      12'hEB9: dout <= 8'b11110000; // 3769 : 240 - 0xf0
      12'hEBA: dout <= 8'b11100000; // 3770 : 224 - 0xe0
      12'hEBB: dout <= 8'b11011101; // 3771 : 221 - 0xdd
      12'hEBC: dout <= 8'b11111010; // 3772 : 250 - 0xfa
      12'hEBD: dout <= 8'b11101011; // 3773 : 235 - 0xeb
      12'hEBE: dout <= 8'b10000000; // 3774 : 128 - 0x80
      12'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xd8
      12'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout <= 8'b00000011; // 3779 :   3 - 0x3
      12'hEC4: dout <= 8'b00000110; // 3780 :   6 - 0x6
      12'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout <= 8'b00000001; // 3782 :   1 - 0x1
      12'hEC7: dout <= 8'b00000001; // 3783 :   1 - 0x1
      12'hEC8: dout <= 8'b00001011; // 3784 :  11 - 0xb -- Background 0xd9
      12'hEC9: dout <= 8'b00000111; // 3785 :   7 - 0x7
      12'hECA: dout <= 8'b00000011; // 3786 :   3 - 0x3
      12'hECB: dout <= 8'b01011101; // 3787 :  93 - 0x5d
      12'hECC: dout <= 8'b10101111; // 3788 : 175 - 0xaf
      12'hECD: dout <= 8'b01010011; // 3789 :  83 - 0x53
      12'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xda
      12'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      12'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      12'hED3: dout <= 8'b10000000; // 3795 : 128 - 0x80
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout <= 8'b01100000; // 3798 :  96 - 0x60
      12'hED7: dout <= 8'b11110000; // 3799 : 240 - 0xf0
      12'hED8: dout <= 8'b11111000; // 3800 : 248 - 0xf8 -- Background 0xdb
      12'hED9: dout <= 8'b11111100; // 3801 : 252 - 0xfc
      12'hEDA: dout <= 8'b11111100; // 3802 : 252 - 0xfc
      12'hEDB: dout <= 8'b11111110; // 3803 : 254 - 0xfe
      12'hEDC: dout <= 8'b11111110; // 3804 : 254 - 0xfe
      12'hEDD: dout <= 8'b11111111; // 3805 : 255 - 0xff
      12'hEDE: dout <= 8'b11111111; // 3806 : 255 - 0xff
      12'hEDF: dout <= 8'b01111110; // 3807 : 126 - 0x7e
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout <= 8'b00100001; // 3814 :  33 - 0x21
      12'hEE7: dout <= 8'b00111111; // 3815 :  63 - 0x3f
      12'hEE8: dout <= 8'b00111111; // 3816 :  63 - 0x3f -- Background 0xdd
      12'hEE9: dout <= 8'b00011111; // 3817 :  31 - 0x1f
      12'hEEA: dout <= 8'b00011111; // 3818 :  31 - 0x1f
      12'hEEB: dout <= 8'b00001111; // 3819 :  15 - 0xf
      12'hEEC: dout <= 8'b00000111; // 3820 :   7 - 0x7
      12'hEED: dout <= 8'b00000011; // 3821 :   3 - 0x3
      12'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b00111110; // 3824 :  62 - 0x3e -- Background 0xde
      12'hEF1: dout <= 8'b00011110; // 3825 :  30 - 0x1e
      12'hEF2: dout <= 8'b00011110; // 3826 :  30 - 0x1e
      12'hEF3: dout <= 8'b00001110; // 3827 :  14 - 0xe
      12'hEF4: dout <= 8'b00001111; // 3828 :  15 - 0xf
      12'hEF5: dout <= 8'b00011111; // 3829 :  31 - 0x1f
      12'hEF6: dout <= 8'b10011111; // 3830 : 159 - 0x9f
      12'hEF7: dout <= 8'b10011111; // 3831 : 159 - 0x9f
      12'hEF8: dout <= 8'b11011111; // 3832 : 223 - 0xdf -- Background 0xdf
      12'hEF9: dout <= 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout <= 8'b11111111; // 3834 : 255 - 0xff
      12'hEFB: dout <= 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout <= 8'b11111111; // 3836 : 255 - 0xff
      12'hEFD: dout <= 8'b11011111; // 3837 : 223 - 0xdf
      12'hEFE: dout <= 8'b11100111; // 3838 : 231 - 0xe7
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b00100000; // 3840 :  32 - 0x20 -- Background 0xe0
      12'hF01: dout <= 8'b00001111; // 3841 :  15 - 0xf
      12'hF02: dout <= 8'b00110000; // 3842 :  48 - 0x30
      12'hF03: dout <= 8'b01000000; // 3843 :  64 - 0x40
      12'hF04: dout <= 8'b10011000; // 3844 : 152 - 0x98
      12'hF05: dout <= 8'b00111110; // 3845 :  62 - 0x3e
      12'hF06: dout <= 8'b00011111; // 3846 :  31 - 0x1f
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b10000001; // 3848 : 129 - 0x81 -- Background 0xe1
      12'hF09: dout <= 8'b00110110; // 3849 :  54 - 0x36
      12'hF0A: dout <= 8'b00101110; // 3850 :  46 - 0x2e
      12'hF0B: dout <= 8'b10101111; // 3851 : 175 - 0xaf
      12'hF0C: dout <= 8'b10101110; // 3852 : 174 - 0xae
      12'hF0D: dout <= 8'b11010001; // 3853 : 209 - 0xd1
      12'hF0E: dout <= 8'b11101111; // 3854 : 239 - 0xef
      12'hF0F: dout <= 8'b10000111; // 3855 : 135 - 0x87
      12'hF10: dout <= 8'b00000010; // 3856 :   2 - 0x2 -- Background 0xe2
      12'hF11: dout <= 8'b11111000; // 3857 : 248 - 0xf8
      12'hF12: dout <= 8'b00000110; // 3858 :   6 - 0x6
      12'hF13: dout <= 8'b00000001; // 3859 :   1 - 0x1
      12'hF14: dout <= 8'b00001100; // 3860 :  12 - 0xc
      12'hF15: dout <= 8'b00111110; // 3861 :  62 - 0x3e
      12'hF16: dout <= 8'b11111100; // 3862 : 252 - 0xfc
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b11000000; // 3864 : 192 - 0xc0 -- Background 0xe3
      12'hF19: dout <= 8'b00110110; // 3865 :  54 - 0x36
      12'hF1A: dout <= 8'b00111110; // 3866 :  62 - 0x3e
      12'hF1B: dout <= 8'b01111010; // 3867 : 122 - 0x7a
      12'hF1C: dout <= 8'b10110110; // 3868 : 182 - 0xb6
      12'hF1D: dout <= 8'b11001101; // 3869 : 205 - 0xcd
      12'hF1E: dout <= 8'b11111011; // 3870 : 251 - 0xfb
      12'hF1F: dout <= 8'b11110000; // 3871 : 240 - 0xf0
      12'hF20: dout <= 8'b00111110; // 3872 :  62 - 0x3e -- Background 0xe4
      12'hF21: dout <= 8'b00111100; // 3873 :  60 - 0x3c
      12'hF22: dout <= 8'b00111100; // 3874 :  60 - 0x3c
      12'hF23: dout <= 8'b00111000; // 3875 :  56 - 0x38
      12'hF24: dout <= 8'b11111000; // 3876 : 248 - 0xf8
      12'hF25: dout <= 8'b01111100; // 3877 : 124 - 0x7c
      12'hF26: dout <= 8'b01111110; // 3878 : 126 - 0x7e
      12'hF27: dout <= 8'b01111000; // 3879 : 120 - 0x78
      12'hF28: dout <= 8'b11111000; // 3880 : 248 - 0xf8 -- Background 0xe5
      12'hF29: dout <= 8'b01111111; // 3881 : 127 - 0x7f
      12'hF2A: dout <= 8'b01111111; // 3882 : 127 - 0x7f
      12'hF2B: dout <= 8'b11111110; // 3883 : 254 - 0xfe
      12'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      12'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      12'hF2E: dout <= 8'b11110011; // 3886 : 243 - 0xf3
      12'hF2F: dout <= 8'b10000001; // 3887 : 129 - 0x81
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xe6
      12'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout <= 8'b00010000; // 3891 :  16 - 0x10
      12'hF34: dout <= 8'b01000000; // 3892 :  64 - 0x40
      12'hF35: dout <= 8'b00100000; // 3893 :  32 - 0x20
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b00000110; // 3896 :   6 - 0x6 -- Background 0xe7
      12'hF39: dout <= 8'b00001110; // 3897 :  14 - 0xe
      12'hF3A: dout <= 8'b01111110; // 3898 : 126 - 0x7e
      12'hF3B: dout <= 8'b11111110; // 3899 : 254 - 0xfe
      12'hF3C: dout <= 8'b11111110; // 3900 : 254 - 0xfe
      12'hF3D: dout <= 8'b11111100; // 3901 : 252 - 0xfc
      12'hF3E: dout <= 8'b11111000; // 3902 : 248 - 0xf8
      12'hF3F: dout <= 8'b11110000; // 3903 : 240 - 0xf0
      12'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xe8
      12'hF41: dout <= 8'b00000000; // 3905 :   0 - 0x0
      12'hF42: dout <= 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout <= 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b00000001; // 3911 :   1 - 0x1
      12'hF48: dout <= 8'b00000010; // 3912 :   2 - 0x2 -- Background 0xe9
      12'hF49: dout <= 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout <= 8'b00001000; // 3914 :   8 - 0x8
      12'hF4B: dout <= 8'b00000001; // 3915 :   1 - 0x1
      12'hF4C: dout <= 8'b00010011; // 3916 :  19 - 0x13
      12'hF4D: dout <= 8'b00000001; // 3917 :   1 - 0x1
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xea
      12'hF51: dout <= 8'b00000000; // 3921 :   0 - 0x0
      12'hF52: dout <= 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout <= 8'b01000011; // 3929 :  67 - 0x43
      12'hF5A: dout <= 8'b01111111; // 3930 : 127 - 0x7f
      12'hF5B: dout <= 8'b01111111; // 3931 : 127 - 0x7f
      12'hF5C: dout <= 8'b01111111; // 3932 : 127 - 0x7f
      12'hF5D: dout <= 8'b00111111; // 3933 :  63 - 0x3f
      12'hF5E: dout <= 8'b00011111; // 3934 :  31 - 0x1f
      12'hF5F: dout <= 8'b00000111; // 3935 :   7 - 0x7
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout <= 8'b11000000; // 3942 : 192 - 0xc0
      12'hF67: dout <= 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout <= 8'b00010000; // 3944 :  16 - 0x10 -- Background 0xed
      12'hF69: dout <= 8'b00111000; // 3945 :  56 - 0x38
      12'hF6A: dout <= 8'b10111111; // 3946 : 191 - 0xbf
      12'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      12'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      12'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      12'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      12'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      12'hF70: dout <= 8'b01111110; // 3952 : 126 - 0x7e -- Background 0xee
      12'hF71: dout <= 8'b00011110; // 3953 :  30 - 0x1e
      12'hF72: dout <= 8'b00011110; // 3954 :  30 - 0x1e
      12'hF73: dout <= 8'b00001110; // 3955 :  14 - 0xe
      12'hF74: dout <= 8'b00001111; // 3956 :  15 - 0xf
      12'hF75: dout <= 8'b00011110; // 3957 :  30 - 0x1e
      12'hF76: dout <= 8'b00011110; // 3958 :  30 - 0x1e
      12'hF77: dout <= 8'b00111110; // 3959 :  62 - 0x3e
      12'hF78: dout <= 8'b01111111; // 3960 : 127 - 0x7f -- Background 0xef
      12'hF79: dout <= 8'b01111111; // 3961 : 127 - 0x7f
      12'hF7A: dout <= 8'b10111111; // 3962 : 191 - 0xbf
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11100111; // 3966 : 231 - 0xe7
      12'hF7F: dout <= 8'b11000000; // 3967 : 192 - 0xc0
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00010000; // 3970 :  16 - 0x10
      12'hF83: dout <= 8'b11111101; // 3971 : 253 - 0xfd
      12'hF84: dout <= 8'b11111010; // 3972 : 250 - 0xfa
      12'hF85: dout <= 8'b11101011; // 3973 : 235 - 0xeb
      12'hF86: dout <= 8'b10000000; // 3974 : 128 - 0x80
      12'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout <= 8'b00100000; // 3976 :  32 - 0x20 -- Background 0xf1
      12'hF89: dout <= 8'b00011111; // 3977 :  31 - 0x1f
      12'hF8A: dout <= 8'b01100000; // 3978 :  96 - 0x60
      12'hF8B: dout <= 8'b10001110; // 3979 : 142 - 0x8e
      12'hF8C: dout <= 8'b00111111; // 3980 :  63 - 0x3f
      12'hF8D: dout <= 8'b01111111; // 3981 : 127 - 0x7f
      12'hF8E: dout <= 8'b01111111; // 3982 : 127 - 0x7f
      12'hF8F: dout <= 8'b01111100; // 3983 : 124 - 0x7c
      12'hF90: dout <= 8'b00111001; // 3984 :  57 - 0x39 -- Background 0xf2
      12'hF91: dout <= 8'b00110110; // 3985 :  54 - 0x36
      12'hF92: dout <= 8'b00101110; // 3986 :  46 - 0x2e
      12'hF93: dout <= 8'b10101111; // 3987 : 175 - 0xaf
      12'hF94: dout <= 8'b10101110; // 3988 : 174 - 0xae
      12'hF95: dout <= 8'b11010001; // 3989 : 209 - 0xd1
      12'hF96: dout <= 8'b11101111; // 3990 : 239 - 0xef
      12'hF97: dout <= 8'b10000111; // 3991 : 135 - 0x87
      12'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0 -- Background 0xf3
      12'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout <= 8'b00000100; // 3994 :   4 - 0x4
      12'hF9B: dout <= 8'b01011111; // 3995 :  95 - 0x5f
      12'hF9C: dout <= 8'b10101111; // 3996 : 175 - 0xaf
      12'hF9D: dout <= 8'b01010011; // 3997 :  83 - 0x53
      12'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b00000010; // 4000 :   2 - 0x2 -- Background 0xf4
      12'hFA1: dout <= 8'b11111100; // 4001 : 252 - 0xfc
      12'hFA2: dout <= 8'b00000011; // 4002 :   3 - 0x3
      12'hFA3: dout <= 8'b00111000; // 4003 :  56 - 0x38
      12'hFA4: dout <= 8'b11111110; // 4004 : 254 - 0xfe
      12'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      12'hFA7: dout <= 8'b00011110; // 4007 :  30 - 0x1e
      12'hFA8: dout <= 8'b11000000; // 4008 : 192 - 0xc0 -- Background 0xf5
      12'hFA9: dout <= 8'b00110110; // 4009 :  54 - 0x36
      12'hFAA: dout <= 8'b00111110; // 4010 :  62 - 0x3e
      12'hFAB: dout <= 8'b01111010; // 4011 : 122 - 0x7a
      12'hFAC: dout <= 8'b10110110; // 4012 : 182 - 0xb6
      12'hFAD: dout <= 8'b11001101; // 4013 : 205 - 0xcd
      12'hFAE: dout <= 8'b11111011; // 4014 : 251 - 0xfb
      12'hFAF: dout <= 8'b11110000; // 4015 : 240 - 0xf0
      12'hFB0: dout <= 8'b00000000; // 4016 :   0 - 0x0 -- Background 0xf6
      12'hFB1: dout <= 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout <= 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout <= 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout <= 8'b00001110; // 4021 :  14 - 0xe
      12'hFB6: dout <= 8'b00001000; // 4022 :   8 - 0x8
      12'hFB7: dout <= 8'b00001000; // 4023 :   8 - 0x8
      12'hFB8: dout <= 8'b00011111; // 4024 :  31 - 0x1f -- Background 0xf7
      12'hFB9: dout <= 8'b00111111; // 4025 :  63 - 0x3f
      12'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      12'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      12'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      12'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      12'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      12'hFBF: dout <= 8'b01111111; // 4031 : 127 - 0x7f
      12'hFC0: dout <= 8'b00111111; // 4032 :  63 - 0x3f -- Background 0xf8
      12'hFC1: dout <= 8'b00111110; // 4033 :  62 - 0x3e
      12'hFC2: dout <= 8'b00111100; // 4034 :  60 - 0x3c
      12'hFC3: dout <= 8'b10111000; // 4035 : 184 - 0xb8
      12'hFC4: dout <= 8'b01111000; // 4036 : 120 - 0x78
      12'hFC5: dout <= 8'b01111000; // 4037 : 120 - 0x78
      12'hFC6: dout <= 8'b01111110; // 4038 : 126 - 0x7e
      12'hFC7: dout <= 8'b01111110; // 4039 : 126 - 0x7e
      12'hFC8: dout <= 8'b11111101; // 4040 : 253 - 0xfd -- Background 0xf9
      12'hFC9: dout <= 8'b01111001; // 4041 : 121 - 0x79
      12'hFCA: dout <= 8'b01111011; // 4042 : 123 - 0x7b
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout <= 8'b11110011; // 4046 : 243 - 0xf3
      12'hFCF: dout <= 8'b10000000; // 4047 : 128 - 0x80
      12'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Background 0xfa
      12'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout <= 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout <= 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout <= 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout <= 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout <= 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout <= 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout <= 8'b00010000; // 4056 :  16 - 0x10 -- Background 0xfb
      12'hFD9: dout <= 8'b10000100; // 4057 : 132 - 0x84
      12'hFDA: dout <= 8'b11100000; // 4058 : 224 - 0xe0
      12'hFDB: dout <= 8'b11000000; // 4059 : 192 - 0xc0
      12'hFDC: dout <= 8'b10000000; // 4060 : 128 - 0x80
      12'hFDD: dout <= 8'b10000000; // 4061 : 128 - 0x80
      12'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b00000000; // 4064 :   0 - 0x0 -- Background 0xfc
      12'hFE1: dout <= 8'b01001000; // 4065 :  72 - 0x48
      12'hFE2: dout <= 8'b00100000; // 4066 :  32 - 0x20
      12'hFE3: dout <= 8'b00000000; // 4067 :   0 - 0x0
      12'hFE4: dout <= 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout <= 8'b00000100; // 4069 :   4 - 0x4
      12'hFE6: dout <= 8'b00001110; // 4070 :  14 - 0xe
      12'hFE7: dout <= 8'b11111110; // 4071 : 254 - 0xfe
      12'hFE8: dout <= 8'b11111110; // 4072 : 254 - 0xfe -- Background 0xfd
      12'hFE9: dout <= 8'b11111100; // 4073 : 252 - 0xfc
      12'hFEA: dout <= 8'b11111100; // 4074 : 252 - 0xfc
      12'hFEB: dout <= 8'b11111000; // 4075 : 248 - 0xf8
      12'hFEC: dout <= 8'b11110000; // 4076 : 240 - 0xf0
      12'hFED: dout <= 8'b11100000; // 4077 : 224 - 0xe0
      12'hFEE: dout <= 8'b10000000; // 4078 : 128 - 0x80
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b00001111; // 4080 :  15 - 0xf -- Background 0xfe
      12'hFF1: dout <= 8'b00000110; // 4081 :   6 - 0x6
      12'hFF2: dout <= 8'b00000110; // 4082 :   6 - 0x6
      12'hFF3: dout <= 8'b00000110; // 4083 :   6 - 0x6
      12'hFF4: dout <= 8'b00000110; // 4084 :   6 - 0x6
      12'hFF5: dout <= 8'b00000110; // 4085 :   6 - 0x6
      12'hFF6: dout <= 8'b00001111; // 4086 :  15 - 0xf
      12'hFF7: dout <= 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout <= 8'b11110000; // 4088 : 240 - 0xf0 -- Background 0xff
      12'hFF9: dout <= 8'b01100000; // 4089 :  96 - 0x60
      12'hFFA: dout <= 8'b01100000; // 4090 :  96 - 0x60
      12'hFFB: dout <= 8'b01100110; // 4091 : 102 - 0x66
      12'hFFC: dout <= 8'b01100110; // 4092 : 102 - 0x66
      12'hFFD: dout <= 8'b01100000; // 4093 :  96 - 0x60
      12'hFFE: dout <= 8'b11110000; // 4094 : 240 - 0xf0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
