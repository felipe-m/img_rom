//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables


//-  Original memory dump file name: lawnmower_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE_LAWN_00
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      11'h0: dout <= 8'b10101001; //    0 : 169 - 0xa9 -- line 0x0
      11'h1: dout <= 8'b10101001; //    1 : 169 - 0xa9
      11'h2: dout <= 8'b10101001; //    2 : 169 - 0xa9
      11'h3: dout <= 8'b10101001; //    3 : 169 - 0xa9
      11'h4: dout <= 8'b10101001; //    4 : 169 - 0xa9
      11'h5: dout <= 8'b10101001; //    5 : 169 - 0xa9
      11'h6: dout <= 8'b10101001; //    6 : 169 - 0xa9
      11'h7: dout <= 8'b10101001; //    7 : 169 - 0xa9
      11'h8: dout <= 8'b10101001; //    8 : 169 - 0xa9
      11'h9: dout <= 8'b10101001; //    9 : 169 - 0xa9
      11'hA: dout <= 8'b10101001; //   10 : 169 - 0xa9
      11'hB: dout <= 8'b10101001; //   11 : 169 - 0xa9
      11'hC: dout <= 8'b10101001; //   12 : 169 - 0xa9
      11'hD: dout <= 8'b10101001; //   13 : 169 - 0xa9
      11'hE: dout <= 8'b10101001; //   14 : 169 - 0xa9
      11'hF: dout <= 8'b10101001; //   15 : 169 - 0xa9
      11'h10: dout <= 8'b10101001; //   16 : 169 - 0xa9
      11'h11: dout <= 8'b10101001; //   17 : 169 - 0xa9
      11'h12: dout <= 8'b10101001; //   18 : 169 - 0xa9
      11'h13: dout <= 8'b10101001; //   19 : 169 - 0xa9
      11'h14: dout <= 8'b10101001; //   20 : 169 - 0xa9
      11'h15: dout <= 8'b10101001; //   21 : 169 - 0xa9
      11'h16: dout <= 8'b10101001; //   22 : 169 - 0xa9
      11'h17: dout <= 8'b10101001; //   23 : 169 - 0xa9
      11'h18: dout <= 8'b10101001; //   24 : 169 - 0xa9
      11'h19: dout <= 8'b10101001; //   25 : 169 - 0xa9
      11'h1A: dout <= 8'b10101001; //   26 : 169 - 0xa9
      11'h1B: dout <= 8'b10101001; //   27 : 169 - 0xa9
      11'h1C: dout <= 8'b10101001; //   28 : 169 - 0xa9
      11'h1D: dout <= 8'b10101001; //   29 : 169 - 0xa9
      11'h1E: dout <= 8'b10101001; //   30 : 169 - 0xa9
      11'h1F: dout <= 8'b10101001; //   31 : 169 - 0xa9
      11'h20: dout <= 8'b10101001; //   32 : 169 - 0xa9 -- line 0x1
      11'h21: dout <= 8'b10101001; //   33 : 169 - 0xa9
      11'h22: dout <= 8'b10101001; //   34 : 169 - 0xa9
      11'h23: dout <= 8'b10101001; //   35 : 169 - 0xa9
      11'h24: dout <= 8'b10101001; //   36 : 169 - 0xa9
      11'h25: dout <= 8'b10101001; //   37 : 169 - 0xa9
      11'h26: dout <= 8'b10101001; //   38 : 169 - 0xa9
      11'h27: dout <= 8'b10101001; //   39 : 169 - 0xa9
      11'h28: dout <= 8'b10101001; //   40 : 169 - 0xa9
      11'h29: dout <= 8'b10101001; //   41 : 169 - 0xa9
      11'h2A: dout <= 8'b10101001; //   42 : 169 - 0xa9
      11'h2B: dout <= 8'b10101001; //   43 : 169 - 0xa9
      11'h2C: dout <= 8'b10101001; //   44 : 169 - 0xa9
      11'h2D: dout <= 8'b10101001; //   45 : 169 - 0xa9
      11'h2E: dout <= 8'b10101001; //   46 : 169 - 0xa9
      11'h2F: dout <= 8'b10101001; //   47 : 169 - 0xa9
      11'h30: dout <= 8'b10101001; //   48 : 169 - 0xa9
      11'h31: dout <= 8'b10101001; //   49 : 169 - 0xa9
      11'h32: dout <= 8'b10101001; //   50 : 169 - 0xa9
      11'h33: dout <= 8'b10101001; //   51 : 169 - 0xa9
      11'h34: dout <= 8'b10101001; //   52 : 169 - 0xa9
      11'h35: dout <= 8'b10101001; //   53 : 169 - 0xa9
      11'h36: dout <= 8'b10101001; //   54 : 169 - 0xa9
      11'h37: dout <= 8'b10101001; //   55 : 169 - 0xa9
      11'h38: dout <= 8'b10101001; //   56 : 169 - 0xa9
      11'h39: dout <= 8'b10101001; //   57 : 169 - 0xa9
      11'h3A: dout <= 8'b10101001; //   58 : 169 - 0xa9
      11'h3B: dout <= 8'b10101001; //   59 : 169 - 0xa9
      11'h3C: dout <= 8'b10101001; //   60 : 169 - 0xa9
      11'h3D: dout <= 8'b10101001; //   61 : 169 - 0xa9
      11'h3E: dout <= 8'b10101001; //   62 : 169 - 0xa9
      11'h3F: dout <= 8'b10101001; //   63 : 169 - 0xa9
      11'h40: dout <= 8'b10101001; //   64 : 169 - 0xa9 -- line 0x2
      11'h41: dout <= 8'b10101001; //   65 : 169 - 0xa9
      11'h42: dout <= 8'b01010110; //   66 :  86 - 0x56
      11'h43: dout <= 8'b01010101; //   67 :  85 - 0x55
      11'h44: dout <= 8'b01010111; //   68 :  87 - 0x57
      11'h45: dout <= 8'b01011000; //   69 :  88 - 0x58
      11'h46: dout <= 8'b11010000; //   70 : 208 - 0xd0
      11'h47: dout <= 8'b11010001; //   71 : 209 - 0xd1
      11'h48: dout <= 8'b10101001; //   72 : 169 - 0xa9
      11'h49: dout <= 8'b01011101; //   73 :  93 - 0x5d
      11'h4A: dout <= 8'b01011110; //   74 :  94 - 0x5e
      11'h4B: dout <= 8'b01011011; //   75 :  91 - 0x5b
      11'h4C: dout <= 8'b01010110; //   76 :  86 - 0x56
      11'h4D: dout <= 8'b11111001; //   77 : 249 - 0xf9
      11'h4E: dout <= 8'b11111010; //   78 : 250 - 0xfa
      11'h4F: dout <= 8'b11111010; //   79 : 250 - 0xfa
      11'h50: dout <= 8'b11111010; //   80 : 250 - 0xfa
      11'h51: dout <= 8'b11111010; //   81 : 250 - 0xfa
      11'h52: dout <= 8'b11111010; //   82 : 250 - 0xfa
      11'h53: dout <= 8'b11111010; //   83 : 250 - 0xfa
      11'h54: dout <= 8'b11111011; //   84 : 251 - 0xfb
      11'h55: dout <= 8'b10101001; //   85 : 169 - 0xa9
      11'h56: dout <= 8'b01011001; //   86 :  89 - 0x59
      11'h57: dout <= 8'b01011010; //   87 :  90 - 0x5a
      11'h58: dout <= 8'b01011000; //   88 :  88 - 0x58
      11'h59: dout <= 8'b01011011; //   89 :  91 - 0x5b
      11'h5A: dout <= 8'b11010000; //   90 : 208 - 0xd0
      11'h5B: dout <= 8'b11010000; //   91 : 208 - 0xd0
      11'h5C: dout <= 8'b11010000; //   92 : 208 - 0xd0
      11'h5D: dout <= 8'b01011100; //   93 :  92 - 0x5c
      11'h5E: dout <= 8'b10101001; //   94 : 169 - 0xa9
      11'h5F: dout <= 8'b10101001; //   95 : 169 - 0xa9
      11'h60: dout <= 8'b10101001; //   96 : 169 - 0xa9 -- line 0x3
      11'h61: dout <= 8'b10101001; //   97 : 169 - 0xa9
      11'h62: dout <= 8'b01100110; //   98 : 102 - 0x66
      11'h63: dout <= 8'b01100101; //   99 : 101 - 0x65
      11'h64: dout <= 8'b01100111; //  100 : 103 - 0x67
      11'h65: dout <= 8'b01101000; //  101 : 104 - 0x68
      11'h66: dout <= 8'b11100000; //  102 : 224 - 0xe0
      11'h67: dout <= 8'b11100001; //  103 : 225 - 0xe1
      11'h68: dout <= 8'b10101001; //  104 : 169 - 0xa9
      11'h69: dout <= 8'b01101101; //  105 : 109 - 0x6d
      11'h6A: dout <= 8'b01101110; //  106 : 110 - 0x6e
      11'h6B: dout <= 8'b01101011; //  107 : 107 - 0x6b
      11'h6C: dout <= 8'b01100110; //  108 : 102 - 0x66
      11'h6D: dout <= 8'b11111100; //  109 : 252 - 0xfc
      11'h6E: dout <= 8'b11111101; //  110 : 253 - 0xfd
      11'h6F: dout <= 8'b11111101; //  111 : 253 - 0xfd
      11'h70: dout <= 8'b11111101; //  112 : 253 - 0xfd
      11'h71: dout <= 8'b11111101; //  113 : 253 - 0xfd
      11'h72: dout <= 8'b11111101; //  114 : 253 - 0xfd
      11'h73: dout <= 8'b11111101; //  115 : 253 - 0xfd
      11'h74: dout <= 8'b11111110; //  116 : 254 - 0xfe
      11'h75: dout <= 8'b10101001; //  117 : 169 - 0xa9
      11'h76: dout <= 8'b01101001; //  118 : 105 - 0x69
      11'h77: dout <= 8'b01101010; //  119 : 106 - 0x6a
      11'h78: dout <= 8'b01101000; //  120 : 104 - 0x68
      11'h79: dout <= 8'b01101011; //  121 : 107 - 0x6b
      11'h7A: dout <= 8'b11100000; //  122 : 224 - 0xe0
      11'h7B: dout <= 8'b11100000; //  123 : 224 - 0xe0
      11'h7C: dout <= 8'b11100000; //  124 : 224 - 0xe0
      11'h7D: dout <= 8'b01101100; //  125 : 108 - 0x6c
      11'h7E: dout <= 8'b10101001; //  126 : 169 - 0xa9
      11'h7F: dout <= 8'b10101001; //  127 : 169 - 0xa9
      11'h80: dout <= 8'b10101010; //  128 : 170 - 0xaa -- line 0x4
      11'h81: dout <= 8'b10101010; //  129 : 170 - 0xaa
      11'h82: dout <= 8'b10101010; //  130 : 170 - 0xaa
      11'h83: dout <= 8'b10101010; //  131 : 170 - 0xaa
      11'h84: dout <= 8'b10101010; //  132 : 170 - 0xaa
      11'h85: dout <= 8'b10101010; //  133 : 170 - 0xaa
      11'h86: dout <= 8'b10101010; //  134 : 170 - 0xaa
      11'h87: dout <= 8'b10101010; //  135 : 170 - 0xaa
      11'h88: dout <= 8'b10101010; //  136 : 170 - 0xaa
      11'h89: dout <= 8'b10101010; //  137 : 170 - 0xaa
      11'h8A: dout <= 8'b10101010; //  138 : 170 - 0xaa
      11'h8B: dout <= 8'b10101010; //  139 : 170 - 0xaa
      11'h8C: dout <= 8'b10101010; //  140 : 170 - 0xaa
      11'h8D: dout <= 8'b10101010; //  141 : 170 - 0xaa
      11'h8E: dout <= 8'b10101010; //  142 : 170 - 0xaa
      11'h8F: dout <= 8'b10101010; //  143 : 170 - 0xaa
      11'h90: dout <= 8'b10101010; //  144 : 170 - 0xaa
      11'h91: dout <= 8'b10101010; //  145 : 170 - 0xaa
      11'h92: dout <= 8'b10101010; //  146 : 170 - 0xaa
      11'h93: dout <= 8'b10101010; //  147 : 170 - 0xaa
      11'h94: dout <= 8'b10101010; //  148 : 170 - 0xaa
      11'h95: dout <= 8'b10101010; //  149 : 170 - 0xaa
      11'h96: dout <= 8'b10101010; //  150 : 170 - 0xaa
      11'h97: dout <= 8'b10101010; //  151 : 170 - 0xaa
      11'h98: dout <= 8'b10101010; //  152 : 170 - 0xaa
      11'h99: dout <= 8'b10101010; //  153 : 170 - 0xaa
      11'h9A: dout <= 8'b10101010; //  154 : 170 - 0xaa
      11'h9B: dout <= 8'b10101010; //  155 : 170 - 0xaa
      11'h9C: dout <= 8'b10101010; //  156 : 170 - 0xaa
      11'h9D: dout <= 8'b10101010; //  157 : 170 - 0xaa
      11'h9E: dout <= 8'b10101010; //  158 : 170 - 0xaa
      11'h9F: dout <= 8'b10101010; //  159 : 170 - 0xaa
      11'hA0: dout <= 8'b10100000; //  160 : 160 - 0xa0 -- line 0x5
      11'hA1: dout <= 8'b10100001; //  161 : 161 - 0xa1
      11'hA2: dout <= 8'b10100010; //  162 : 162 - 0xa2
      11'hA3: dout <= 8'b10100010; //  163 : 162 - 0xa2
      11'hA4: dout <= 8'b10100010; //  164 : 162 - 0xa2
      11'hA5: dout <= 8'b10100010; //  165 : 162 - 0xa2
      11'hA6: dout <= 8'b10100010; //  166 : 162 - 0xa2
      11'hA7: dout <= 8'b10100010; //  167 : 162 - 0xa2
      11'hA8: dout <= 8'b10100010; //  168 : 162 - 0xa2
      11'hA9: dout <= 8'b10100010; //  169 : 162 - 0xa2
      11'hAA: dout <= 8'b10100010; //  170 : 162 - 0xa2
      11'hAB: dout <= 8'b10100010; //  171 : 162 - 0xa2
      11'hAC: dout <= 8'b10100010; //  172 : 162 - 0xa2
      11'hAD: dout <= 8'b10100010; //  173 : 162 - 0xa2
      11'hAE: dout <= 8'b10100010; //  174 : 162 - 0xa2
      11'hAF: dout <= 8'b10100010; //  175 : 162 - 0xa2
      11'hB0: dout <= 8'b10100010; //  176 : 162 - 0xa2
      11'hB1: dout <= 8'b10100010; //  177 : 162 - 0xa2
      11'hB2: dout <= 8'b10100010; //  178 : 162 - 0xa2
      11'hB3: dout <= 8'b10100010; //  179 : 162 - 0xa2
      11'hB4: dout <= 8'b10100010; //  180 : 162 - 0xa2
      11'hB5: dout <= 8'b10100010; //  181 : 162 - 0xa2
      11'hB6: dout <= 8'b10100010; //  182 : 162 - 0xa2
      11'hB7: dout <= 8'b10100010; //  183 : 162 - 0xa2
      11'hB8: dout <= 8'b10100010; //  184 : 162 - 0xa2
      11'hB9: dout <= 8'b10100010; //  185 : 162 - 0xa2
      11'hBA: dout <= 8'b10100010; //  186 : 162 - 0xa2
      11'hBB: dout <= 8'b10100010; //  187 : 162 - 0xa2
      11'hBC: dout <= 8'b10100010; //  188 : 162 - 0xa2
      11'hBD: dout <= 8'b10100010; //  189 : 162 - 0xa2
      11'hBE: dout <= 8'b10100110; //  190 : 166 - 0xa6
      11'hBF: dout <= 8'b10100000; //  191 : 160 - 0xa0
      11'hC0: dout <= 8'b10100000; //  192 : 160 - 0xa0 -- line 0x6
      11'hC1: dout <= 8'b10100011; //  193 : 163 - 0xa3
      11'hC2: dout <= 8'b10000000; //  194 : 128 - 0x80
      11'hC3: dout <= 8'b10000001; //  195 : 129 - 0x81
      11'hC4: dout <= 8'b10000000; //  196 : 128 - 0x80
      11'hC5: dout <= 8'b10000001; //  197 : 129 - 0x81
      11'hC6: dout <= 8'b10000000; //  198 : 128 - 0x80
      11'hC7: dout <= 8'b10000010; //  199 : 130 - 0x82
      11'hC8: dout <= 8'b10000000; //  200 : 128 - 0x80
      11'hC9: dout <= 8'b10000001; //  201 : 129 - 0x81
      11'hCA: dout <= 8'b10000001; //  202 : 129 - 0x81
      11'hCB: dout <= 8'b10000000; //  203 : 128 - 0x80
      11'hCC: dout <= 8'b10000000; //  204 : 128 - 0x80
      11'hCD: dout <= 8'b10000001; //  205 : 129 - 0x81
      11'hCE: dout <= 8'b10000010; //  206 : 130 - 0x82
      11'hCF: dout <= 8'b10000011; //  207 : 131 - 0x83
      11'hD0: dout <= 8'b10000010; //  208 : 130 - 0x82
      11'hD1: dout <= 8'b10000011; //  209 : 131 - 0x83
      11'hD2: dout <= 8'b10000000; //  210 : 128 - 0x80
      11'hD3: dout <= 8'b10000010; //  211 : 130 - 0x82
      11'hD4: dout <= 8'b10000000; //  212 : 128 - 0x80
      11'hD5: dout <= 8'b10000010; //  213 : 130 - 0x82
      11'hD6: dout <= 8'b10000010; //  214 : 130 - 0x82
      11'hD7: dout <= 8'b10000011; //  215 : 131 - 0x83
      11'hD8: dout <= 8'b10000010; //  216 : 130 - 0x82
      11'hD9: dout <= 8'b10000011; //  217 : 131 - 0x83
      11'hDA: dout <= 8'b10000001; //  218 : 129 - 0x81
      11'hDB: dout <= 8'b10000000; //  219 : 128 - 0x80
      11'hDC: dout <= 8'b10000000; //  220 : 128 - 0x80
      11'hDD: dout <= 8'b10000001; //  221 : 129 - 0x81
      11'hDE: dout <= 8'b10100111; //  222 : 167 - 0xa7
      11'hDF: dout <= 8'b10100000; //  223 : 160 - 0xa0
      11'hE0: dout <= 8'b10100000; //  224 : 160 - 0xa0 -- line 0x7
      11'hE1: dout <= 8'b10100011; //  225 : 163 - 0xa3
      11'hE2: dout <= 8'b10010000; //  226 : 144 - 0x90
      11'hE3: dout <= 8'b10010001; //  227 : 145 - 0x91
      11'hE4: dout <= 8'b10010000; //  228 : 144 - 0x90
      11'hE5: dout <= 8'b10010001; //  229 : 145 - 0x91
      11'hE6: dout <= 8'b10010010; //  230 : 146 - 0x92
      11'hE7: dout <= 8'b10010001; //  231 : 145 - 0x91
      11'hE8: dout <= 8'b10010000; //  232 : 144 - 0x90
      11'hE9: dout <= 8'b10010001; //  233 : 145 - 0x91
      11'hEA: dout <= 8'b10010011; //  234 : 147 - 0x93
      11'hEB: dout <= 8'b10010010; //  235 : 146 - 0x92
      11'hEC: dout <= 8'b10010000; //  236 : 144 - 0x90
      11'hED: dout <= 8'b10010001; //  237 : 145 - 0x91
      11'hEE: dout <= 8'b10010010; //  238 : 146 - 0x92
      11'hEF: dout <= 8'b10010011; //  239 : 147 - 0x93
      11'hF0: dout <= 8'b10010010; //  240 : 146 - 0x92
      11'hF1: dout <= 8'b10010011; //  241 : 147 - 0x93
      11'hF2: dout <= 8'b10010010; //  242 : 146 - 0x92
      11'hF3: dout <= 8'b10010001; //  243 : 145 - 0x91
      11'hF4: dout <= 8'b10010010; //  244 : 146 - 0x92
      11'hF5: dout <= 8'b10010001; //  245 : 145 - 0x91
      11'hF6: dout <= 8'b10010010; //  246 : 146 - 0x92
      11'hF7: dout <= 8'b10010011; //  247 : 147 - 0x93
      11'hF8: dout <= 8'b10010010; //  248 : 146 - 0x92
      11'hF9: dout <= 8'b10010011; //  249 : 147 - 0x93
      11'hFA: dout <= 8'b10010011; //  250 : 147 - 0x93
      11'hFB: dout <= 8'b10010010; //  251 : 146 - 0x92
      11'hFC: dout <= 8'b10010000; //  252 : 144 - 0x90
      11'hFD: dout <= 8'b10010001; //  253 : 145 - 0x91
      11'hFE: dout <= 8'b10100111; //  254 : 167 - 0xa7
      11'hFF: dout <= 8'b10100000; //  255 : 160 - 0xa0
      11'h100: dout <= 8'b10100000; //  256 : 160 - 0xa0 -- line 0x8
      11'h101: dout <= 8'b10100011; //  257 : 163 - 0xa3
      11'h102: dout <= 8'b10000010; //  258 : 130 - 0x82
      11'h103: dout <= 8'b10000011; //  259 : 131 - 0x83
      11'h104: dout <= 8'b10000101; //  260 : 133 - 0x85
      11'h105: dout <= 8'b10000110; //  261 : 134 - 0x86
      11'h106: dout <= 8'b10000101; //  262 : 133 - 0x85
      11'h107: dout <= 8'b10000110; //  263 : 134 - 0x86
      11'h108: dout <= 8'b10000101; //  264 : 133 - 0x85
      11'h109: dout <= 8'b10000110; //  265 : 134 - 0x86
      11'h10A: dout <= 8'b10000101; //  266 : 133 - 0x85
      11'h10B: dout <= 8'b10000110; //  267 : 134 - 0x86
      11'h10C: dout <= 8'b10000100; //  268 : 132 - 0x84
      11'h10D: dout <= 8'b10000111; //  269 : 135 - 0x87
      11'h10E: dout <= 8'b10000110; //  270 : 134 - 0x86
      11'h10F: dout <= 8'b10000111; //  271 : 135 - 0x87
      11'h110: dout <= 8'b10000100; //  272 : 132 - 0x84
      11'h111: dout <= 8'b10000101; //  273 : 133 - 0x85
      11'h112: dout <= 8'b10000101; //  274 : 133 - 0x85
      11'h113: dout <= 8'b10000110; //  275 : 134 - 0x86
      11'h114: dout <= 8'b10000101; //  276 : 133 - 0x85
      11'h115: dout <= 8'b10000110; //  277 : 134 - 0x86
      11'h116: dout <= 8'b10000110; //  278 : 134 - 0x86
      11'h117: dout <= 8'b10000111; //  279 : 135 - 0x87
      11'h118: dout <= 8'b10000110; //  280 : 134 - 0x86
      11'h119: dout <= 8'b10000111; //  281 : 135 - 0x87
      11'h11A: dout <= 8'b10000100; //  282 : 132 - 0x84
      11'h11B: dout <= 8'b10000101; //  283 : 133 - 0x85
      11'h11C: dout <= 8'b10000010; //  284 : 130 - 0x82
      11'h11D: dout <= 8'b10000011; //  285 : 131 - 0x83
      11'h11E: dout <= 8'b10100111; //  286 : 167 - 0xa7
      11'h11F: dout <= 8'b10100000; //  287 : 160 - 0xa0
      11'h120: dout <= 8'b10100000; //  288 : 160 - 0xa0 -- line 0x9
      11'h121: dout <= 8'b10100011; //  289 : 163 - 0xa3
      11'h122: dout <= 8'b10010010; //  290 : 146 - 0x92
      11'h123: dout <= 8'b10010011; //  291 : 147 - 0x93
      11'h124: dout <= 8'b10010111; //  292 : 151 - 0x97
      11'h125: dout <= 8'b10010100; //  293 : 148 - 0x94
      11'h126: dout <= 8'b10010111; //  294 : 151 - 0x97
      11'h127: dout <= 8'b10010100; //  295 : 148 - 0x94
      11'h128: dout <= 8'b10010111; //  296 : 151 - 0x97
      11'h129: dout <= 8'b10010100; //  297 : 148 - 0x94
      11'h12A: dout <= 8'b10010111; //  298 : 151 - 0x97
      11'h12B: dout <= 8'b10010100; //  299 : 148 - 0x94
      11'h12C: dout <= 8'b10010110; //  300 : 150 - 0x96
      11'h12D: dout <= 8'b10010101; //  301 : 149 - 0x95
      11'h12E: dout <= 8'b10010110; //  302 : 150 - 0x96
      11'h12F: dout <= 8'b10010111; //  303 : 151 - 0x97
      11'h130: dout <= 8'b10010100; //  304 : 148 - 0x94
      11'h131: dout <= 8'b10010101; //  305 : 149 - 0x95
      11'h132: dout <= 8'b10010111; //  306 : 151 - 0x97
      11'h133: dout <= 8'b10010100; //  307 : 148 - 0x94
      11'h134: dout <= 8'b10010111; //  308 : 151 - 0x97
      11'h135: dout <= 8'b10010100; //  309 : 148 - 0x94
      11'h136: dout <= 8'b10010110; //  310 : 150 - 0x96
      11'h137: dout <= 8'b10010111; //  311 : 151 - 0x97
      11'h138: dout <= 8'b10010110; //  312 : 150 - 0x96
      11'h139: dout <= 8'b10010111; //  313 : 151 - 0x97
      11'h13A: dout <= 8'b10010100; //  314 : 148 - 0x94
      11'h13B: dout <= 8'b10010101; //  315 : 149 - 0x95
      11'h13C: dout <= 8'b10010010; //  316 : 146 - 0x92
      11'h13D: dout <= 8'b10010011; //  317 : 147 - 0x93
      11'h13E: dout <= 8'b10100111; //  318 : 167 - 0xa7
      11'h13F: dout <= 8'b10100000; //  319 : 160 - 0xa0
      11'h140: dout <= 8'b10100000; //  320 : 160 - 0xa0 -- line 0xa
      11'h141: dout <= 8'b10100011; //  321 : 163 - 0xa3
      11'h142: dout <= 8'b10000000; //  322 : 128 - 0x80
      11'h143: dout <= 8'b10000010; //  323 : 130 - 0x82
      11'h144: dout <= 8'b10000100; //  324 : 132 - 0x84
      11'h145: dout <= 8'b10000111; //  325 : 135 - 0x87
      11'h146: dout <= 8'b10000101; //  326 : 133 - 0x85
      11'h147: dout <= 8'b10000110; //  327 : 134 - 0x86
      11'h148: dout <= 8'b10000100; //  328 : 132 - 0x84
      11'h149: dout <= 8'b10000111; //  329 : 135 - 0x87
      11'h14A: dout <= 8'b10000100; //  330 : 132 - 0x84
      11'h14B: dout <= 8'b10000111; //  331 : 135 - 0x87
      11'h14C: dout <= 8'b10000110; //  332 : 134 - 0x86
      11'h14D: dout <= 8'b10000111; //  333 : 135 - 0x87
      11'h14E: dout <= 8'b10000100; //  334 : 132 - 0x84
      11'h14F: dout <= 8'b10000101; //  335 : 133 - 0x85
      11'h150: dout <= 8'b10000100; //  336 : 132 - 0x84
      11'h151: dout <= 8'b10000101; //  337 : 133 - 0x85
      11'h152: dout <= 8'b10000110; //  338 : 134 - 0x86
      11'h153: dout <= 8'b10000111; //  339 : 135 - 0x87
      11'h154: dout <= 8'b10000100; //  340 : 132 - 0x84
      11'h155: dout <= 8'b10000101; //  341 : 133 - 0x85
      11'h156: dout <= 8'b10000101; //  342 : 133 - 0x85
      11'h157: dout <= 8'b10000110; //  343 : 134 - 0x86
      11'h158: dout <= 8'b10000100; //  344 : 132 - 0x84
      11'h159: dout <= 8'b10000111; //  345 : 135 - 0x87
      11'h15A: dout <= 8'b10000100; //  346 : 132 - 0x84
      11'h15B: dout <= 8'b10000111; //  347 : 135 - 0x87
      11'h15C: dout <= 8'b10000000; //  348 : 128 - 0x80
      11'h15D: dout <= 8'b10000001; //  349 : 129 - 0x81
      11'h15E: dout <= 8'b10100111; //  350 : 167 - 0xa7
      11'h15F: dout <= 8'b10100000; //  351 : 160 - 0xa0
      11'h160: dout <= 8'b10100000; //  352 : 160 - 0xa0 -- line 0xb
      11'h161: dout <= 8'b10100011; //  353 : 163 - 0xa3
      11'h162: dout <= 8'b10010010; //  354 : 146 - 0x92
      11'h163: dout <= 8'b10010001; //  355 : 145 - 0x91
      11'h164: dout <= 8'b10010110; //  356 : 150 - 0x96
      11'h165: dout <= 8'b10010101; //  357 : 149 - 0x95
      11'h166: dout <= 8'b10010111; //  358 : 151 - 0x97
      11'h167: dout <= 8'b10010100; //  359 : 148 - 0x94
      11'h168: dout <= 8'b10010110; //  360 : 150 - 0x96
      11'h169: dout <= 8'b10010101; //  361 : 149 - 0x95
      11'h16A: dout <= 8'b10010110; //  362 : 150 - 0x96
      11'h16B: dout <= 8'b10010101; //  363 : 149 - 0x95
      11'h16C: dout <= 8'b10010110; //  364 : 150 - 0x96
      11'h16D: dout <= 8'b10010111; //  365 : 151 - 0x97
      11'h16E: dout <= 8'b10010100; //  366 : 148 - 0x94
      11'h16F: dout <= 8'b10010101; //  367 : 149 - 0x95
      11'h170: dout <= 8'b10010100; //  368 : 148 - 0x94
      11'h171: dout <= 8'b10010101; //  369 : 149 - 0x95
      11'h172: dout <= 8'b10010110; //  370 : 150 - 0x96
      11'h173: dout <= 8'b10010111; //  371 : 151 - 0x97
      11'h174: dout <= 8'b10010100; //  372 : 148 - 0x94
      11'h175: dout <= 8'b10010101; //  373 : 149 - 0x95
      11'h176: dout <= 8'b10010111; //  374 : 151 - 0x97
      11'h177: dout <= 8'b10010100; //  375 : 148 - 0x94
      11'h178: dout <= 8'b10010110; //  376 : 150 - 0x96
      11'h179: dout <= 8'b10010101; //  377 : 149 - 0x95
      11'h17A: dout <= 8'b10010110; //  378 : 150 - 0x96
      11'h17B: dout <= 8'b10010101; //  379 : 149 - 0x95
      11'h17C: dout <= 8'b10010000; //  380 : 144 - 0x90
      11'h17D: dout <= 8'b10010001; //  381 : 145 - 0x91
      11'h17E: dout <= 8'b10100111; //  382 : 167 - 0xa7
      11'h17F: dout <= 8'b10100000; //  383 : 160 - 0xa0
      11'h180: dout <= 8'b10100000; //  384 : 160 - 0xa0 -- line 0xc
      11'h181: dout <= 8'b10100011; //  385 : 163 - 0xa3
      11'h182: dout <= 8'b10000010; //  386 : 130 - 0x82
      11'h183: dout <= 8'b10000011; //  387 : 131 - 0x83
      11'h184: dout <= 8'b10000110; //  388 : 134 - 0x86
      11'h185: dout <= 8'b10000111; //  389 : 135 - 0x87
      11'h186: dout <= 8'b10000100; //  390 : 132 - 0x84
      11'h187: dout <= 8'b10000101; //  391 : 133 - 0x85
      11'h188: dout <= 8'b10000100; //  392 : 132 - 0x84
      11'h189: dout <= 8'b10000111; //  393 : 135 - 0x87
      11'h18A: dout <= 8'b10000100; //  394 : 132 - 0x84
      11'h18B: dout <= 8'b10000111; //  395 : 135 - 0x87
      11'h18C: dout <= 8'b10000110; //  396 : 134 - 0x86
      11'h18D: dout <= 8'b10000111; //  397 : 135 - 0x87
      11'h18E: dout <= 8'b10000100; //  398 : 132 - 0x84
      11'h18F: dout <= 8'b10000111; //  399 : 135 - 0x87
      11'h190: dout <= 8'b10000110; //  400 : 134 - 0x86
      11'h191: dout <= 8'b10000111; //  401 : 135 - 0x87
      11'h192: dout <= 8'b10000110; //  402 : 134 - 0x86
      11'h193: dout <= 8'b10000111; //  403 : 135 - 0x87
      11'h194: dout <= 8'b10000110; //  404 : 134 - 0x86
      11'h195: dout <= 8'b10000111; //  405 : 135 - 0x87
      11'h196: dout <= 8'b10000110; //  406 : 134 - 0x86
      11'h197: dout <= 8'b10000111; //  407 : 135 - 0x87
      11'h198: dout <= 8'b10000101; //  408 : 133 - 0x85
      11'h199: dout <= 8'b10000110; //  409 : 134 - 0x86
      11'h19A: dout <= 8'b10000100; //  410 : 132 - 0x84
      11'h19B: dout <= 8'b10000111; //  411 : 135 - 0x87
      11'h19C: dout <= 8'b10000000; //  412 : 128 - 0x80
      11'h19D: dout <= 8'b10000010; //  413 : 130 - 0x82
      11'h19E: dout <= 8'b10100111; //  414 : 167 - 0xa7
      11'h19F: dout <= 8'b10100000; //  415 : 160 - 0xa0
      11'h1A0: dout <= 8'b10100000; //  416 : 160 - 0xa0 -- line 0xd
      11'h1A1: dout <= 8'b10100011; //  417 : 163 - 0xa3
      11'h1A2: dout <= 8'b10010010; //  418 : 146 - 0x92
      11'h1A3: dout <= 8'b10010011; //  419 : 147 - 0x93
      11'h1A4: dout <= 8'b10010110; //  420 : 150 - 0x96
      11'h1A5: dout <= 8'b10010111; //  421 : 151 - 0x97
      11'h1A6: dout <= 8'b10010100; //  422 : 148 - 0x94
      11'h1A7: dout <= 8'b10010101; //  423 : 149 - 0x95
      11'h1A8: dout <= 8'b10010110; //  424 : 150 - 0x96
      11'h1A9: dout <= 8'b10010101; //  425 : 149 - 0x95
      11'h1AA: dout <= 8'b10010110; //  426 : 150 - 0x96
      11'h1AB: dout <= 8'b10010101; //  427 : 149 - 0x95
      11'h1AC: dout <= 8'b10010110; //  428 : 150 - 0x96
      11'h1AD: dout <= 8'b10010111; //  429 : 151 - 0x97
      11'h1AE: dout <= 8'b10010110; //  430 : 150 - 0x96
      11'h1AF: dout <= 8'b10010101; //  431 : 149 - 0x95
      11'h1B0: dout <= 8'b10010110; //  432 : 150 - 0x96
      11'h1B1: dout <= 8'b10010111; //  433 : 151 - 0x97
      11'h1B2: dout <= 8'b10010110; //  434 : 150 - 0x96
      11'h1B3: dout <= 8'b10010111; //  435 : 151 - 0x97
      11'h1B4: dout <= 8'b10010110; //  436 : 150 - 0x96
      11'h1B5: dout <= 8'b10010111; //  437 : 151 - 0x97
      11'h1B6: dout <= 8'b10010110; //  438 : 150 - 0x96
      11'h1B7: dout <= 8'b10010111; //  439 : 151 - 0x97
      11'h1B8: dout <= 8'b10010111; //  440 : 151 - 0x97
      11'h1B9: dout <= 8'b10010100; //  441 : 148 - 0x94
      11'h1BA: dout <= 8'b10010110; //  442 : 150 - 0x96
      11'h1BB: dout <= 8'b10010101; //  443 : 149 - 0x95
      11'h1BC: dout <= 8'b10010010; //  444 : 146 - 0x92
      11'h1BD: dout <= 8'b10010001; //  445 : 145 - 0x91
      11'h1BE: dout <= 8'b10100111; //  446 : 167 - 0xa7
      11'h1BF: dout <= 8'b10100000; //  447 : 160 - 0xa0
      11'h1C0: dout <= 8'b10100000; //  448 : 160 - 0xa0 -- line 0xe
      11'h1C1: dout <= 8'b10100011; //  449 : 163 - 0xa3
      11'h1C2: dout <= 8'b10000000; //  450 : 128 - 0x80
      11'h1C3: dout <= 8'b10000001; //  451 : 129 - 0x81
      11'h1C4: dout <= 8'b10000101; //  452 : 133 - 0x85
      11'h1C5: dout <= 8'b10000110; //  453 : 134 - 0x86
      11'h1C6: dout <= 8'b10000100; //  454 : 132 - 0x84
      11'h1C7: dout <= 8'b10000101; //  455 : 133 - 0x85
      11'h1C8: dout <= 8'b10000100; //  456 : 132 - 0x84
      11'h1C9: dout <= 8'b10000101; //  457 : 133 - 0x85
      11'h1CA: dout <= 8'b10000100; //  458 : 132 - 0x84
      11'h1CB: dout <= 8'b10000111; //  459 : 135 - 0x87
      11'h1CC: dout <= 8'b10000001; //  460 : 129 - 0x81
      11'h1CD: dout <= 8'b10000000; //  461 : 128 - 0x80
      11'h1CE: dout <= 8'b10000010; //  462 : 130 - 0x82
      11'h1CF: dout <= 8'b10000011; //  463 : 131 - 0x83
      11'h1D0: dout <= 8'b10000010; //  464 : 130 - 0x82
      11'h1D1: dout <= 8'b10000011; //  465 : 131 - 0x83
      11'h1D2: dout <= 8'b10000001; //  466 : 129 - 0x81
      11'h1D3: dout <= 8'b10000000; //  467 : 128 - 0x80
      11'h1D4: dout <= 8'b10000101; //  468 : 133 - 0x85
      11'h1D5: dout <= 8'b10000110; //  469 : 134 - 0x86
      11'h1D6: dout <= 8'b10000110; //  470 : 134 - 0x86
      11'h1D7: dout <= 8'b10000111; //  471 : 135 - 0x87
      11'h1D8: dout <= 8'b10000100; //  472 : 132 - 0x84
      11'h1D9: dout <= 8'b10000111; //  473 : 135 - 0x87
      11'h1DA: dout <= 8'b10000100; //  474 : 132 - 0x84
      11'h1DB: dout <= 8'b10000111; //  475 : 135 - 0x87
      11'h1DC: dout <= 8'b10000000; //  476 : 128 - 0x80
      11'h1DD: dout <= 8'b10000001; //  477 : 129 - 0x81
      11'h1DE: dout <= 8'b10100111; //  478 : 167 - 0xa7
      11'h1DF: dout <= 8'b10100000; //  479 : 160 - 0xa0
      11'h1E0: dout <= 8'b10100000; //  480 : 160 - 0xa0 -- line 0xf
      11'h1E1: dout <= 8'b10100011; //  481 : 163 - 0xa3
      11'h1E2: dout <= 8'b10010000; //  482 : 144 - 0x90
      11'h1E3: dout <= 8'b10010001; //  483 : 145 - 0x91
      11'h1E4: dout <= 8'b10010111; //  484 : 151 - 0x97
      11'h1E5: dout <= 8'b10010100; //  485 : 148 - 0x94
      11'h1E6: dout <= 8'b10010100; //  486 : 148 - 0x94
      11'h1E7: dout <= 8'b10010101; //  487 : 149 - 0x95
      11'h1E8: dout <= 8'b10010100; //  488 : 148 - 0x94
      11'h1E9: dout <= 8'b10010101; //  489 : 149 - 0x95
      11'h1EA: dout <= 8'b10010110; //  490 : 150 - 0x96
      11'h1EB: dout <= 8'b10010101; //  491 : 149 - 0x95
      11'h1EC: dout <= 8'b10010011; //  492 : 147 - 0x93
      11'h1ED: dout <= 8'b10010010; //  493 : 146 - 0x92
      11'h1EE: dout <= 8'b10010010; //  494 : 146 - 0x92
      11'h1EF: dout <= 8'b10010011; //  495 : 147 - 0x93
      11'h1F0: dout <= 8'b10010010; //  496 : 146 - 0x92
      11'h1F1: dout <= 8'b10010011; //  497 : 147 - 0x93
      11'h1F2: dout <= 8'b10010011; //  498 : 147 - 0x93
      11'h1F3: dout <= 8'b10010010; //  499 : 146 - 0x92
      11'h1F4: dout <= 8'b10010111; //  500 : 151 - 0x97
      11'h1F5: dout <= 8'b10010100; //  501 : 148 - 0x94
      11'h1F6: dout <= 8'b10010110; //  502 : 150 - 0x96
      11'h1F7: dout <= 8'b10010111; //  503 : 151 - 0x97
      11'h1F8: dout <= 8'b10010110; //  504 : 150 - 0x96
      11'h1F9: dout <= 8'b10010101; //  505 : 149 - 0x95
      11'h1FA: dout <= 8'b10010110; //  506 : 150 - 0x96
      11'h1FB: dout <= 8'b10010101; //  507 : 149 - 0x95
      11'h1FC: dout <= 8'b10010000; //  508 : 144 - 0x90
      11'h1FD: dout <= 8'b10010001; //  509 : 145 - 0x91
      11'h1FE: dout <= 8'b10100111; //  510 : 167 - 0xa7
      11'h1FF: dout <= 8'b10100000; //  511 : 160 - 0xa0
      11'h200: dout <= 8'b10100000; //  512 : 160 - 0xa0 -- line 0x10
      11'h201: dout <= 8'b10100011; //  513 : 163 - 0xa3
      11'h202: dout <= 8'b10000010; //  514 : 130 - 0x82
      11'h203: dout <= 8'b10000011; //  515 : 131 - 0x83
      11'h204: dout <= 8'b10000101; //  516 : 133 - 0x85
      11'h205: dout <= 8'b10000110; //  517 : 134 - 0x86
      11'h206: dout <= 8'b10000101; //  518 : 133 - 0x85
      11'h207: dout <= 8'b10000110; //  519 : 134 - 0x86
      11'h208: dout <= 8'b10000101; //  520 : 133 - 0x85
      11'h209: dout <= 8'b10000110; //  521 : 134 - 0x86
      11'h20A: dout <= 8'b10000101; //  522 : 133 - 0x85
      11'h20B: dout <= 8'b10000110; //  523 : 134 - 0x86
      11'h20C: dout <= 8'b10000000; //  524 : 128 - 0x80
      11'h20D: dout <= 8'b10000010; //  525 : 130 - 0x82
      11'h20E: dout <= 8'b10000010; //  526 : 130 - 0x82
      11'h20F: dout <= 8'b10000011; //  527 : 131 - 0x83
      11'h210: dout <= 8'b10000000; //  528 : 128 - 0x80
      11'h211: dout <= 8'b10000001; //  529 : 129 - 0x81
      11'h212: dout <= 8'b10000001; //  530 : 129 - 0x81
      11'h213: dout <= 8'b10000000; //  531 : 128 - 0x80
      11'h214: dout <= 8'b10000101; //  532 : 133 - 0x85
      11'h215: dout <= 8'b10000110; //  533 : 134 - 0x86
      11'h216: dout <= 8'b10000110; //  534 : 134 - 0x86
      11'h217: dout <= 8'b10000111; //  535 : 135 - 0x87
      11'h218: dout <= 8'b10000110; //  536 : 134 - 0x86
      11'h219: dout <= 8'b10000111; //  537 : 135 - 0x87
      11'h21A: dout <= 8'b10000100; //  538 : 132 - 0x84
      11'h21B: dout <= 8'b10000101; //  539 : 133 - 0x85
      11'h21C: dout <= 8'b10000010; //  540 : 130 - 0x82
      11'h21D: dout <= 8'b10000011; //  541 : 131 - 0x83
      11'h21E: dout <= 8'b10100111; //  542 : 167 - 0xa7
      11'h21F: dout <= 8'b10100000; //  543 : 160 - 0xa0
      11'h220: dout <= 8'b10100000; //  544 : 160 - 0xa0 -- line 0x11
      11'h221: dout <= 8'b10100011; //  545 : 163 - 0xa3
      11'h222: dout <= 8'b10010010; //  546 : 146 - 0x92
      11'h223: dout <= 8'b10010011; //  547 : 147 - 0x93
      11'h224: dout <= 8'b10010111; //  548 : 151 - 0x97
      11'h225: dout <= 8'b10010100; //  549 : 148 - 0x94
      11'h226: dout <= 8'b10010111; //  550 : 151 - 0x97
      11'h227: dout <= 8'b10010100; //  551 : 148 - 0x94
      11'h228: dout <= 8'b10010111; //  552 : 151 - 0x97
      11'h229: dout <= 8'b10010100; //  553 : 148 - 0x94
      11'h22A: dout <= 8'b10010111; //  554 : 151 - 0x97
      11'h22B: dout <= 8'b10010100; //  555 : 148 - 0x94
      11'h22C: dout <= 8'b10010010; //  556 : 146 - 0x92
      11'h22D: dout <= 8'b10010001; //  557 : 145 - 0x91
      11'h22E: dout <= 8'b10010010; //  558 : 146 - 0x92
      11'h22F: dout <= 8'b10010011; //  559 : 147 - 0x93
      11'h230: dout <= 8'b10010000; //  560 : 144 - 0x90
      11'h231: dout <= 8'b10010001; //  561 : 145 - 0x91
      11'h232: dout <= 8'b10010011; //  562 : 147 - 0x93
      11'h233: dout <= 8'b10010010; //  563 : 146 - 0x92
      11'h234: dout <= 8'b10010111; //  564 : 151 - 0x97
      11'h235: dout <= 8'b10010100; //  565 : 148 - 0x94
      11'h236: dout <= 8'b10010110; //  566 : 150 - 0x96
      11'h237: dout <= 8'b10010111; //  567 : 151 - 0x97
      11'h238: dout <= 8'b10010110; //  568 : 150 - 0x96
      11'h239: dout <= 8'b10010111; //  569 : 151 - 0x97
      11'h23A: dout <= 8'b10010100; //  570 : 148 - 0x94
      11'h23B: dout <= 8'b10010101; //  571 : 149 - 0x95
      11'h23C: dout <= 8'b10010010; //  572 : 146 - 0x92
      11'h23D: dout <= 8'b10010011; //  573 : 147 - 0x93
      11'h23E: dout <= 8'b10100111; //  574 : 167 - 0xa7
      11'h23F: dout <= 8'b10100000; //  575 : 160 - 0xa0
      11'h240: dout <= 8'b10100000; //  576 : 160 - 0xa0 -- line 0x12
      11'h241: dout <= 8'b10100011; //  577 : 163 - 0xa3
      11'h242: dout <= 8'b10000000; //  578 : 128 - 0x80
      11'h243: dout <= 8'b10000010; //  579 : 130 - 0x82
      11'h244: dout <= 8'b10000100; //  580 : 132 - 0x84
      11'h245: dout <= 8'b10000111; //  581 : 135 - 0x87
      11'h246: dout <= 8'b10000101; //  582 : 133 - 0x85
      11'h247: dout <= 8'b10000110; //  583 : 134 - 0x86
      11'h248: dout <= 8'b10000100; //  584 : 132 - 0x84
      11'h249: dout <= 8'b10000111; //  585 : 135 - 0x87
      11'h24A: dout <= 8'b10000100; //  586 : 132 - 0x84
      11'h24B: dout <= 8'b10000111; //  587 : 135 - 0x87
      11'h24C: dout <= 8'b10000010; //  588 : 130 - 0x82
      11'h24D: dout <= 8'b10000011; //  589 : 131 - 0x83
      11'h24E: dout <= 8'b10000000; //  590 : 128 - 0x80
      11'h24F: dout <= 8'b10000001; //  591 : 129 - 0x81
      11'h250: dout <= 8'b10000000; //  592 : 128 - 0x80
      11'h251: dout <= 8'b10000001; //  593 : 129 - 0x81
      11'h252: dout <= 8'b10000010; //  594 : 130 - 0x82
      11'h253: dout <= 8'b10000011; //  595 : 131 - 0x83
      11'h254: dout <= 8'b10000100; //  596 : 132 - 0x84
      11'h255: dout <= 8'b10000101; //  597 : 133 - 0x85
      11'h256: dout <= 8'b10000101; //  598 : 133 - 0x85
      11'h257: dout <= 8'b10000110; //  599 : 134 - 0x86
      11'h258: dout <= 8'b10000100; //  600 : 132 - 0x84
      11'h259: dout <= 8'b10000111; //  601 : 135 - 0x87
      11'h25A: dout <= 8'b10000100; //  602 : 132 - 0x84
      11'h25B: dout <= 8'b10000111; //  603 : 135 - 0x87
      11'h25C: dout <= 8'b10000000; //  604 : 128 - 0x80
      11'h25D: dout <= 8'b10000001; //  605 : 129 - 0x81
      11'h25E: dout <= 8'b10100111; //  606 : 167 - 0xa7
      11'h25F: dout <= 8'b10100000; //  607 : 160 - 0xa0
      11'h260: dout <= 8'b10100000; //  608 : 160 - 0xa0 -- line 0x13
      11'h261: dout <= 8'b10100011; //  609 : 163 - 0xa3
      11'h262: dout <= 8'b10010010; //  610 : 146 - 0x92
      11'h263: dout <= 8'b10010001; //  611 : 145 - 0x91
      11'h264: dout <= 8'b10010110; //  612 : 150 - 0x96
      11'h265: dout <= 8'b10010101; //  613 : 149 - 0x95
      11'h266: dout <= 8'b10010111; //  614 : 151 - 0x97
      11'h267: dout <= 8'b10010100; //  615 : 148 - 0x94
      11'h268: dout <= 8'b10010110; //  616 : 150 - 0x96
      11'h269: dout <= 8'b10010101; //  617 : 149 - 0x95
      11'h26A: dout <= 8'b10010110; //  618 : 150 - 0x96
      11'h26B: dout <= 8'b10010101; //  619 : 149 - 0x95
      11'h26C: dout <= 8'b10010010; //  620 : 146 - 0x92
      11'h26D: dout <= 8'b10010011; //  621 : 147 - 0x93
      11'h26E: dout <= 8'b10010000; //  622 : 144 - 0x90
      11'h26F: dout <= 8'b10010001; //  623 : 145 - 0x91
      11'h270: dout <= 8'b10010000; //  624 : 144 - 0x90
      11'h271: dout <= 8'b10010001; //  625 : 145 - 0x91
      11'h272: dout <= 8'b10010010; //  626 : 146 - 0x92
      11'h273: dout <= 8'b10010011; //  627 : 147 - 0x93
      11'h274: dout <= 8'b10010100; //  628 : 148 - 0x94
      11'h275: dout <= 8'b10010101; //  629 : 149 - 0x95
      11'h276: dout <= 8'b10010111; //  630 : 151 - 0x97
      11'h277: dout <= 8'b10010100; //  631 : 148 - 0x94
      11'h278: dout <= 8'b10010110; //  632 : 150 - 0x96
      11'h279: dout <= 8'b10010101; //  633 : 149 - 0x95
      11'h27A: dout <= 8'b10010110; //  634 : 150 - 0x96
      11'h27B: dout <= 8'b10010101; //  635 : 149 - 0x95
      11'h27C: dout <= 8'b10010000; //  636 : 144 - 0x90
      11'h27D: dout <= 8'b10010001; //  637 : 145 - 0x91
      11'h27E: dout <= 8'b10100111; //  638 : 167 - 0xa7
      11'h27F: dout <= 8'b10100000; //  639 : 160 - 0xa0
      11'h280: dout <= 8'b10100000; //  640 : 160 - 0xa0 -- line 0x14
      11'h281: dout <= 8'b10100011; //  641 : 163 - 0xa3
      11'h282: dout <= 8'b10000010; //  642 : 130 - 0x82
      11'h283: dout <= 8'b10000011; //  643 : 131 - 0x83
      11'h284: dout <= 8'b10000110; //  644 : 134 - 0x86
      11'h285: dout <= 8'b10000111; //  645 : 135 - 0x87
      11'h286: dout <= 8'b10000100; //  646 : 132 - 0x84
      11'h287: dout <= 8'b10000101; //  647 : 133 - 0x85
      11'h288: dout <= 8'b10000100; //  648 : 132 - 0x84
      11'h289: dout <= 8'b10000111; //  649 : 135 - 0x87
      11'h28A: dout <= 8'b10000100; //  650 : 132 - 0x84
      11'h28B: dout <= 8'b10000111; //  651 : 135 - 0x87
      11'h28C: dout <= 8'b10000110; //  652 : 134 - 0x86
      11'h28D: dout <= 8'b10000111; //  653 : 135 - 0x87
      11'h28E: dout <= 8'b10000100; //  654 : 132 - 0x84
      11'h28F: dout <= 8'b10000111; //  655 : 135 - 0x87
      11'h290: dout <= 8'b10000110; //  656 : 134 - 0x86
      11'h291: dout <= 8'b10000111; //  657 : 135 - 0x87
      11'h292: dout <= 8'b10000110; //  658 : 134 - 0x86
      11'h293: dout <= 8'b10000111; //  659 : 135 - 0x87
      11'h294: dout <= 8'b10000110; //  660 : 134 - 0x86
      11'h295: dout <= 8'b10000111; //  661 : 135 - 0x87
      11'h296: dout <= 8'b10000110; //  662 : 134 - 0x86
      11'h297: dout <= 8'b10000111; //  663 : 135 - 0x87
      11'h298: dout <= 8'b10000101; //  664 : 133 - 0x85
      11'h299: dout <= 8'b10000110; //  665 : 134 - 0x86
      11'h29A: dout <= 8'b10000100; //  666 : 132 - 0x84
      11'h29B: dout <= 8'b10000111; //  667 : 135 - 0x87
      11'h29C: dout <= 8'b10000000; //  668 : 128 - 0x80
      11'h29D: dout <= 8'b10000010; //  669 : 130 - 0x82
      11'h29E: dout <= 8'b10100111; //  670 : 167 - 0xa7
      11'h29F: dout <= 8'b10100000; //  671 : 160 - 0xa0
      11'h2A0: dout <= 8'b10100000; //  672 : 160 - 0xa0 -- line 0x15
      11'h2A1: dout <= 8'b10100011; //  673 : 163 - 0xa3
      11'h2A2: dout <= 8'b10010010; //  674 : 146 - 0x92
      11'h2A3: dout <= 8'b10010011; //  675 : 147 - 0x93
      11'h2A4: dout <= 8'b10010110; //  676 : 150 - 0x96
      11'h2A5: dout <= 8'b10010111; //  677 : 151 - 0x97
      11'h2A6: dout <= 8'b10010100; //  678 : 148 - 0x94
      11'h2A7: dout <= 8'b10010101; //  679 : 149 - 0x95
      11'h2A8: dout <= 8'b10010110; //  680 : 150 - 0x96
      11'h2A9: dout <= 8'b10010101; //  681 : 149 - 0x95
      11'h2AA: dout <= 8'b10010110; //  682 : 150 - 0x96
      11'h2AB: dout <= 8'b10010101; //  683 : 149 - 0x95
      11'h2AC: dout <= 8'b10010110; //  684 : 150 - 0x96
      11'h2AD: dout <= 8'b10010111; //  685 : 151 - 0x97
      11'h2AE: dout <= 8'b10010110; //  686 : 150 - 0x96
      11'h2AF: dout <= 8'b10010101; //  687 : 149 - 0x95
      11'h2B0: dout <= 8'b10010110; //  688 : 150 - 0x96
      11'h2B1: dout <= 8'b10010111; //  689 : 151 - 0x97
      11'h2B2: dout <= 8'b10010110; //  690 : 150 - 0x96
      11'h2B3: dout <= 8'b10010111; //  691 : 151 - 0x97
      11'h2B4: dout <= 8'b10010110; //  692 : 150 - 0x96
      11'h2B5: dout <= 8'b10010111; //  693 : 151 - 0x97
      11'h2B6: dout <= 8'b10010110; //  694 : 150 - 0x96
      11'h2B7: dout <= 8'b10010111; //  695 : 151 - 0x97
      11'h2B8: dout <= 8'b10010111; //  696 : 151 - 0x97
      11'h2B9: dout <= 8'b10010100; //  697 : 148 - 0x94
      11'h2BA: dout <= 8'b10010110; //  698 : 150 - 0x96
      11'h2BB: dout <= 8'b10010101; //  699 : 149 - 0x95
      11'h2BC: dout <= 8'b10010010; //  700 : 146 - 0x92
      11'h2BD: dout <= 8'b10010001; //  701 : 145 - 0x91
      11'h2BE: dout <= 8'b10100111; //  702 : 167 - 0xa7
      11'h2BF: dout <= 8'b10100000; //  703 : 160 - 0xa0
      11'h2C0: dout <= 8'b10100000; //  704 : 160 - 0xa0 -- line 0x16
      11'h2C1: dout <= 8'b10100011; //  705 : 163 - 0xa3
      11'h2C2: dout <= 8'b10000000; //  706 : 128 - 0x80
      11'h2C3: dout <= 8'b10000001; //  707 : 129 - 0x81
      11'h2C4: dout <= 8'b10000101; //  708 : 133 - 0x85
      11'h2C5: dout <= 8'b10000110; //  709 : 134 - 0x86
      11'h2C6: dout <= 8'b10000100; //  710 : 132 - 0x84
      11'h2C7: dout <= 8'b10000101; //  711 : 133 - 0x85
      11'h2C8: dout <= 8'b10000100; //  712 : 132 - 0x84
      11'h2C9: dout <= 8'b10000101; //  713 : 133 - 0x85
      11'h2CA: dout <= 8'b10000100; //  714 : 132 - 0x84
      11'h2CB: dout <= 8'b10000111; //  715 : 135 - 0x87
      11'h2CC: dout <= 8'b10000101; //  716 : 133 - 0x85
      11'h2CD: dout <= 8'b10000110; //  717 : 134 - 0x86
      11'h2CE: dout <= 8'b10000110; //  718 : 134 - 0x86
      11'h2CF: dout <= 8'b10000111; //  719 : 135 - 0x87
      11'h2D0: dout <= 8'b10000110; //  720 : 134 - 0x86
      11'h2D1: dout <= 8'b10000111; //  721 : 135 - 0x87
      11'h2D2: dout <= 8'b10000101; //  722 : 133 - 0x85
      11'h2D3: dout <= 8'b10000110; //  723 : 134 - 0x86
      11'h2D4: dout <= 8'b10000101; //  724 : 133 - 0x85
      11'h2D5: dout <= 8'b10000110; //  725 : 134 - 0x86
      11'h2D6: dout <= 8'b10000110; //  726 : 134 - 0x86
      11'h2D7: dout <= 8'b10000111; //  727 : 135 - 0x87
      11'h2D8: dout <= 8'b10000100; //  728 : 132 - 0x84
      11'h2D9: dout <= 8'b10000111; //  729 : 135 - 0x87
      11'h2DA: dout <= 8'b10000100; //  730 : 132 - 0x84
      11'h2DB: dout <= 8'b10000111; //  731 : 135 - 0x87
      11'h2DC: dout <= 8'b10000000; //  732 : 128 - 0x80
      11'h2DD: dout <= 8'b10000001; //  733 : 129 - 0x81
      11'h2DE: dout <= 8'b10100111; //  734 : 167 - 0xa7
      11'h2DF: dout <= 8'b10100000; //  735 : 160 - 0xa0
      11'h2E0: dout <= 8'b10100000; //  736 : 160 - 0xa0 -- line 0x17
      11'h2E1: dout <= 8'b10100011; //  737 : 163 - 0xa3
      11'h2E2: dout <= 8'b10010000; //  738 : 144 - 0x90
      11'h2E3: dout <= 8'b10010001; //  739 : 145 - 0x91
      11'h2E4: dout <= 8'b10010111; //  740 : 151 - 0x97
      11'h2E5: dout <= 8'b10010100; //  741 : 148 - 0x94
      11'h2E6: dout <= 8'b10010100; //  742 : 148 - 0x94
      11'h2E7: dout <= 8'b10010101; //  743 : 149 - 0x95
      11'h2E8: dout <= 8'b10010100; //  744 : 148 - 0x94
      11'h2E9: dout <= 8'b10010101; //  745 : 149 - 0x95
      11'h2EA: dout <= 8'b10010110; //  746 : 150 - 0x96
      11'h2EB: dout <= 8'b10010101; //  747 : 149 - 0x95
      11'h2EC: dout <= 8'b10010111; //  748 : 151 - 0x97
      11'h2ED: dout <= 8'b10010100; //  749 : 148 - 0x94
      11'h2EE: dout <= 8'b10010110; //  750 : 150 - 0x96
      11'h2EF: dout <= 8'b10010111; //  751 : 151 - 0x97
      11'h2F0: dout <= 8'b10010110; //  752 : 150 - 0x96
      11'h2F1: dout <= 8'b10010111; //  753 : 151 - 0x97
      11'h2F2: dout <= 8'b10010111; //  754 : 151 - 0x97
      11'h2F3: dout <= 8'b10010100; //  755 : 148 - 0x94
      11'h2F4: dout <= 8'b10010111; //  756 : 151 - 0x97
      11'h2F5: dout <= 8'b10010100; //  757 : 148 - 0x94
      11'h2F6: dout <= 8'b10010110; //  758 : 150 - 0x96
      11'h2F7: dout <= 8'b10010111; //  759 : 151 - 0x97
      11'h2F8: dout <= 8'b10010110; //  760 : 150 - 0x96
      11'h2F9: dout <= 8'b10010101; //  761 : 149 - 0x95
      11'h2FA: dout <= 8'b10010110; //  762 : 150 - 0x96
      11'h2FB: dout <= 8'b10010101; //  763 : 149 - 0x95
      11'h2FC: dout <= 8'b10010000; //  764 : 144 - 0x90
      11'h2FD: dout <= 8'b10010001; //  765 : 145 - 0x91
      11'h2FE: dout <= 8'b10100111; //  766 : 167 - 0xa7
      11'h2FF: dout <= 8'b10100000; //  767 : 160 - 0xa0
      11'h300: dout <= 8'b10100000; //  768 : 160 - 0xa0 -- line 0x18
      11'h301: dout <= 8'b10100011; //  769 : 163 - 0xa3
      11'h302: dout <= 8'b10000000; //  770 : 128 - 0x80
      11'h303: dout <= 8'b10000010; //  771 : 130 - 0x82
      11'h304: dout <= 8'b10000100; //  772 : 132 - 0x84
      11'h305: dout <= 8'b10000111; //  773 : 135 - 0x87
      11'h306: dout <= 8'b10000100; //  774 : 132 - 0x84
      11'h307: dout <= 8'b10000111; //  775 : 135 - 0x87
      11'h308: dout <= 8'b10000100; //  776 : 132 - 0x84
      11'h309: dout <= 8'b10000111; //  777 : 135 - 0x87
      11'h30A: dout <= 8'b10000110; //  778 : 134 - 0x86
      11'h30B: dout <= 8'b10000111; //  779 : 135 - 0x87
      11'h30C: dout <= 8'b10000101; //  780 : 133 - 0x85
      11'h30D: dout <= 8'b10000110; //  781 : 134 - 0x86
      11'h30E: dout <= 8'b10000100; //  782 : 132 - 0x84
      11'h30F: dout <= 8'b10000111; //  783 : 135 - 0x87
      11'h310: dout <= 8'b10000100; //  784 : 132 - 0x84
      11'h311: dout <= 8'b10000101; //  785 : 133 - 0x85
      11'h312: dout <= 8'b10000100; //  786 : 132 - 0x84
      11'h313: dout <= 8'b10000111; //  787 : 135 - 0x87
      11'h314: dout <= 8'b10000110; //  788 : 134 - 0x86
      11'h315: dout <= 8'b10000111; //  789 : 135 - 0x87
      11'h316: dout <= 8'b10000110; //  790 : 134 - 0x86
      11'h317: dout <= 8'b10000111; //  791 : 135 - 0x87
      11'h318: dout <= 8'b10000100; //  792 : 132 - 0x84
      11'h319: dout <= 8'b10000111; //  793 : 135 - 0x87
      11'h31A: dout <= 8'b10000101; //  794 : 133 - 0x85
      11'h31B: dout <= 8'b10000110; //  795 : 134 - 0x86
      11'h31C: dout <= 8'b10000000; //  796 : 128 - 0x80
      11'h31D: dout <= 8'b10000010; //  797 : 130 - 0x82
      11'h31E: dout <= 8'b10100111; //  798 : 167 - 0xa7
      11'h31F: dout <= 8'b10100000; //  799 : 160 - 0xa0
      11'h320: dout <= 8'b10100000; //  800 : 160 - 0xa0 -- line 0x19
      11'h321: dout <= 8'b10100011; //  801 : 163 - 0xa3
      11'h322: dout <= 8'b10010010; //  802 : 146 - 0x92
      11'h323: dout <= 8'b10010001; //  803 : 145 - 0x91
      11'h324: dout <= 8'b10010110; //  804 : 150 - 0x96
      11'h325: dout <= 8'b10010101; //  805 : 149 - 0x95
      11'h326: dout <= 8'b10010110; //  806 : 150 - 0x96
      11'h327: dout <= 8'b10010101; //  807 : 149 - 0x95
      11'h328: dout <= 8'b10010110; //  808 : 150 - 0x96
      11'h329: dout <= 8'b10010101; //  809 : 149 - 0x95
      11'h32A: dout <= 8'b10010110; //  810 : 150 - 0x96
      11'h32B: dout <= 8'b10010111; //  811 : 151 - 0x97
      11'h32C: dout <= 8'b10010111; //  812 : 151 - 0x97
      11'h32D: dout <= 8'b10010100; //  813 : 148 - 0x94
      11'h32E: dout <= 8'b10010110; //  814 : 150 - 0x96
      11'h32F: dout <= 8'b10010101; //  815 : 149 - 0x95
      11'h330: dout <= 8'b10010100; //  816 : 148 - 0x94
      11'h331: dout <= 8'b10010101; //  817 : 149 - 0x95
      11'h332: dout <= 8'b10010110; //  818 : 150 - 0x96
      11'h333: dout <= 8'b10010101; //  819 : 149 - 0x95
      11'h334: dout <= 8'b10010110; //  820 : 150 - 0x96
      11'h335: dout <= 8'b10010111; //  821 : 151 - 0x97
      11'h336: dout <= 8'b10010110; //  822 : 150 - 0x96
      11'h337: dout <= 8'b10010111; //  823 : 151 - 0x97
      11'h338: dout <= 8'b10010110; //  824 : 150 - 0x96
      11'h339: dout <= 8'b10010101; //  825 : 149 - 0x95
      11'h33A: dout <= 8'b10010111; //  826 : 151 - 0x97
      11'h33B: dout <= 8'b10010100; //  827 : 148 - 0x94
      11'h33C: dout <= 8'b10010010; //  828 : 146 - 0x92
      11'h33D: dout <= 8'b10010001; //  829 : 145 - 0x91
      11'h33E: dout <= 8'b10100111; //  830 : 167 - 0xa7
      11'h33F: dout <= 8'b10100000; //  831 : 160 - 0xa0
      11'h340: dout <= 8'b10100000; //  832 : 160 - 0xa0 -- line 0x1a
      11'h341: dout <= 8'b10100011; //  833 : 163 - 0xa3
      11'h342: dout <= 8'b10000001; //  834 : 129 - 0x81
      11'h343: dout <= 8'b10000000; //  835 : 128 - 0x80
      11'h344: dout <= 8'b10000000; //  836 : 128 - 0x80
      11'h345: dout <= 8'b10000001; //  837 : 129 - 0x81
      11'h346: dout <= 8'b10000010; //  838 : 130 - 0x82
      11'h347: dout <= 8'b10000011; //  839 : 131 - 0x83
      11'h348: dout <= 8'b10000001; //  840 : 129 - 0x81
      11'h349: dout <= 8'b10000000; //  841 : 128 - 0x80
      11'h34A: dout <= 8'b10000001; //  842 : 129 - 0x81
      11'h34B: dout <= 8'b10000000; //  843 : 128 - 0x80
      11'h34C: dout <= 8'b10000000; //  844 : 128 - 0x80
      11'h34D: dout <= 8'b10000010; //  845 : 130 - 0x82
      11'h34E: dout <= 8'b10000000; //  846 : 128 - 0x80
      11'h34F: dout <= 8'b10000001; //  847 : 129 - 0x81
      11'h350: dout <= 8'b10000001; //  848 : 129 - 0x81
      11'h351: dout <= 8'b10000000; //  849 : 128 - 0x80
      11'h352: dout <= 8'b10000000; //  850 : 128 - 0x80
      11'h353: dout <= 8'b10000010; //  851 : 130 - 0x82
      11'h354: dout <= 8'b10000000; //  852 : 128 - 0x80
      11'h355: dout <= 8'b10000001; //  853 : 129 - 0x81
      11'h356: dout <= 8'b10000010; //  854 : 130 - 0x82
      11'h357: dout <= 8'b10000011; //  855 : 131 - 0x83
      11'h358: dout <= 8'b10000001; //  856 : 129 - 0x81
      11'h359: dout <= 8'b10000000; //  857 : 128 - 0x80
      11'h35A: dout <= 8'b10000000; //  858 : 128 - 0x80
      11'h35B: dout <= 8'b10000001; //  859 : 129 - 0x81
      11'h35C: dout <= 8'b10000000; //  860 : 128 - 0x80
      11'h35D: dout <= 8'b10000001; //  861 : 129 - 0x81
      11'h35E: dout <= 8'b10100111; //  862 : 167 - 0xa7
      11'h35F: dout <= 8'b10100000; //  863 : 160 - 0xa0
      11'h360: dout <= 8'b10100000; //  864 : 160 - 0xa0 -- line 0x1b
      11'h361: dout <= 8'b10100011; //  865 : 163 - 0xa3
      11'h362: dout <= 8'b10010011; //  866 : 147 - 0x93
      11'h363: dout <= 8'b10010010; //  867 : 146 - 0x92
      11'h364: dout <= 8'b10010000; //  868 : 144 - 0x90
      11'h365: dout <= 8'b10010001; //  869 : 145 - 0x91
      11'h366: dout <= 8'b10010010; //  870 : 146 - 0x92
      11'h367: dout <= 8'b10010011; //  871 : 147 - 0x93
      11'h368: dout <= 8'b10010011; //  872 : 147 - 0x93
      11'h369: dout <= 8'b10010010; //  873 : 146 - 0x92
      11'h36A: dout <= 8'b10010011; //  874 : 147 - 0x93
      11'h36B: dout <= 8'b10010010; //  875 : 146 - 0x92
      11'h36C: dout <= 8'b10010010; //  876 : 146 - 0x92
      11'h36D: dout <= 8'b10010001; //  877 : 145 - 0x91
      11'h36E: dout <= 8'b10010000; //  878 : 144 - 0x90
      11'h36F: dout <= 8'b10010001; //  879 : 145 - 0x91
      11'h370: dout <= 8'b10010011; //  880 : 147 - 0x93
      11'h371: dout <= 8'b10010010; //  881 : 146 - 0x92
      11'h372: dout <= 8'b10010010; //  882 : 146 - 0x92
      11'h373: dout <= 8'b10010001; //  883 : 145 - 0x91
      11'h374: dout <= 8'b10010000; //  884 : 144 - 0x90
      11'h375: dout <= 8'b10010001; //  885 : 145 - 0x91
      11'h376: dout <= 8'b10010010; //  886 : 146 - 0x92
      11'h377: dout <= 8'b10010011; //  887 : 147 - 0x93
      11'h378: dout <= 8'b10010011; //  888 : 147 - 0x93
      11'h379: dout <= 8'b10010010; //  889 : 146 - 0x92
      11'h37A: dout <= 8'b10010000; //  890 : 144 - 0x90
      11'h37B: dout <= 8'b10010001; //  891 : 145 - 0x91
      11'h37C: dout <= 8'b10010000; //  892 : 144 - 0x90
      11'h37D: dout <= 8'b10010001; //  893 : 145 - 0x91
      11'h37E: dout <= 8'b10100111; //  894 : 167 - 0xa7
      11'h37F: dout <= 8'b10100000; //  895 : 160 - 0xa0
      11'h380: dout <= 8'b10100000; //  896 : 160 - 0xa0 -- line 0x1c
      11'h381: dout <= 8'b10100100; //  897 : 164 - 0xa4
      11'h382: dout <= 8'b10100101; //  898 : 165 - 0xa5
      11'h383: dout <= 8'b10100101; //  899 : 165 - 0xa5
      11'h384: dout <= 8'b10100101; //  900 : 165 - 0xa5
      11'h385: dout <= 8'b10100101; //  901 : 165 - 0xa5
      11'h386: dout <= 8'b10100101; //  902 : 165 - 0xa5
      11'h387: dout <= 8'b10100101; //  903 : 165 - 0xa5
      11'h388: dout <= 8'b10100101; //  904 : 165 - 0xa5
      11'h389: dout <= 8'b10100101; //  905 : 165 - 0xa5
      11'h38A: dout <= 8'b10100101; //  906 : 165 - 0xa5
      11'h38B: dout <= 8'b10100101; //  907 : 165 - 0xa5
      11'h38C: dout <= 8'b10100101; //  908 : 165 - 0xa5
      11'h38D: dout <= 8'b10100101; //  909 : 165 - 0xa5
      11'h38E: dout <= 8'b10100101; //  910 : 165 - 0xa5
      11'h38F: dout <= 8'b10100101; //  911 : 165 - 0xa5
      11'h390: dout <= 8'b10100101; //  912 : 165 - 0xa5
      11'h391: dout <= 8'b10100101; //  913 : 165 - 0xa5
      11'h392: dout <= 8'b10100101; //  914 : 165 - 0xa5
      11'h393: dout <= 8'b10100101; //  915 : 165 - 0xa5
      11'h394: dout <= 8'b10100101; //  916 : 165 - 0xa5
      11'h395: dout <= 8'b10100101; //  917 : 165 - 0xa5
      11'h396: dout <= 8'b10100101; //  918 : 165 - 0xa5
      11'h397: dout <= 8'b10100101; //  919 : 165 - 0xa5
      11'h398: dout <= 8'b10100101; //  920 : 165 - 0xa5
      11'h399: dout <= 8'b10100101; //  921 : 165 - 0xa5
      11'h39A: dout <= 8'b10100101; //  922 : 165 - 0xa5
      11'h39B: dout <= 8'b10100101; //  923 : 165 - 0xa5
      11'h39C: dout <= 8'b10100101; //  924 : 165 - 0xa5
      11'h39D: dout <= 8'b10100101; //  925 : 165 - 0xa5
      11'h39E: dout <= 8'b10101000; //  926 : 168 - 0xa8
      11'h39F: dout <= 8'b10100000; //  927 : 160 - 0xa0
      11'h3A0: dout <= 8'b10100000; //  928 : 160 - 0xa0 -- line 0x1d
      11'h3A1: dout <= 8'b10100000; //  929 : 160 - 0xa0
      11'h3A2: dout <= 8'b10100000; //  930 : 160 - 0xa0
      11'h3A3: dout <= 8'b10100000; //  931 : 160 - 0xa0
      11'h3A4: dout <= 8'b10100000; //  932 : 160 - 0xa0
      11'h3A5: dout <= 8'b10100000; //  933 : 160 - 0xa0
      11'h3A6: dout <= 8'b10100000; //  934 : 160 - 0xa0
      11'h3A7: dout <= 8'b10100000; //  935 : 160 - 0xa0
      11'h3A8: dout <= 8'b10100000; //  936 : 160 - 0xa0
      11'h3A9: dout <= 8'b10100000; //  937 : 160 - 0xa0
      11'h3AA: dout <= 8'b10100000; //  938 : 160 - 0xa0
      11'h3AB: dout <= 8'b10100000; //  939 : 160 - 0xa0
      11'h3AC: dout <= 8'b10100000; //  940 : 160 - 0xa0
      11'h3AD: dout <= 8'b10100000; //  941 : 160 - 0xa0
      11'h3AE: dout <= 8'b10100000; //  942 : 160 - 0xa0
      11'h3AF: dout <= 8'b10100000; //  943 : 160 - 0xa0
      11'h3B0: dout <= 8'b10100000; //  944 : 160 - 0xa0
      11'h3B1: dout <= 8'b10100000; //  945 : 160 - 0xa0
      11'h3B2: dout <= 8'b10100000; //  946 : 160 - 0xa0
      11'h3B3: dout <= 8'b10100000; //  947 : 160 - 0xa0
      11'h3B4: dout <= 8'b10100000; //  948 : 160 - 0xa0
      11'h3B5: dout <= 8'b10100000; //  949 : 160 - 0xa0
      11'h3B6: dout <= 8'b10100000; //  950 : 160 - 0xa0
      11'h3B7: dout <= 8'b10100000; //  951 : 160 - 0xa0
      11'h3B8: dout <= 8'b10100000; //  952 : 160 - 0xa0
      11'h3B9: dout <= 8'b10100000; //  953 : 160 - 0xa0
      11'h3BA: dout <= 8'b10100000; //  954 : 160 - 0xa0
      11'h3BB: dout <= 8'b10100000; //  955 : 160 - 0xa0
      11'h3BC: dout <= 8'b10100000; //  956 : 160 - 0xa0
      11'h3BD: dout <= 8'b10100000; //  957 : 160 - 0xa0
      11'h3BE: dout <= 8'b10100000; //  958 : 160 - 0xa0
      11'h3BF: dout <= 8'b10100000; //  959 : 160 - 0xa0
        //-- Attribute Table 0----
      11'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0
      11'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout <= 8'b10000000; //  968 : 128 - 0x80
      11'h3C9: dout <= 8'b10100000; //  969 : 160 - 0xa0
      11'h3CA: dout <= 8'b10100000; //  970 : 160 - 0xa0
      11'h3CB: dout <= 8'b10100000; //  971 : 160 - 0xa0
      11'h3CC: dout <= 8'b10100000; //  972 : 160 - 0xa0
      11'h3CD: dout <= 8'b10100000; //  973 : 160 - 0xa0
      11'h3CE: dout <= 8'b10100000; //  974 : 160 - 0xa0
      11'h3CF: dout <= 8'b00100000; //  975 :  32 - 0x20
      11'h3D0: dout <= 8'b10001000; //  976 : 136 - 0x88
      11'h3D1: dout <= 8'b10101010; //  977 : 170 - 0xaa
      11'h3D2: dout <= 8'b10101010; //  978 : 170 - 0xaa
      11'h3D3: dout <= 8'b10101010; //  979 : 170 - 0xaa
      11'h3D4: dout <= 8'b10101010; //  980 : 170 - 0xaa
      11'h3D5: dout <= 8'b10101010; //  981 : 170 - 0xaa
      11'h3D6: dout <= 8'b10101010; //  982 : 170 - 0xaa
      11'h3D7: dout <= 8'b00100010; //  983 :  34 - 0x22
      11'h3D8: dout <= 8'b10001000; //  984 : 136 - 0x88
      11'h3D9: dout <= 8'b10101010; //  985 : 170 - 0xaa
      11'h3DA: dout <= 8'b10101010; //  986 : 170 - 0xaa
      11'h3DB: dout <= 8'b10101010; //  987 : 170 - 0xaa
      11'h3DC: dout <= 8'b10101010; //  988 : 170 - 0xaa
      11'h3DD: dout <= 8'b10101010; //  989 : 170 - 0xaa
      11'h3DE: dout <= 8'b10101010; //  990 : 170 - 0xaa
      11'h3DF: dout <= 8'b00100010; //  991 :  34 - 0x22
      11'h3E0: dout <= 8'b10001000; //  992 : 136 - 0x88
      11'h3E1: dout <= 8'b10101010; //  993 : 170 - 0xaa
      11'h3E2: dout <= 8'b10101010; //  994 : 170 - 0xaa
      11'h3E3: dout <= 8'b10101010; //  995 : 170 - 0xaa
      11'h3E4: dout <= 8'b10101010; //  996 : 170 - 0xaa
      11'h3E5: dout <= 8'b10101010; //  997 : 170 - 0xaa
      11'h3E6: dout <= 8'b10101010; //  998 : 170 - 0xaa
      11'h3E7: dout <= 8'b00100010; //  999 :  34 - 0x22
      11'h3E8: dout <= 8'b10001000; // 1000 : 136 - 0x88
      11'h3E9: dout <= 8'b10101010; // 1001 : 170 - 0xaa
      11'h3EA: dout <= 8'b10101010; // 1002 : 170 - 0xaa
      11'h3EB: dout <= 8'b10101010; // 1003 : 170 - 0xaa
      11'h3EC: dout <= 8'b10101010; // 1004 : 170 - 0xaa
      11'h3ED: dout <= 8'b10101010; // 1005 : 170 - 0xaa
      11'h3EE: dout <= 8'b10101010; // 1006 : 170 - 0xaa
      11'h3EF: dout <= 8'b00100010; // 1007 :  34 - 0x22
      11'h3F0: dout <= 8'b10001000; // 1008 : 136 - 0x88
      11'h3F1: dout <= 8'b10101010; // 1009 : 170 - 0xaa
      11'h3F2: dout <= 8'b10101010; // 1010 : 170 - 0xaa
      11'h3F3: dout <= 8'b10101010; // 1011 : 170 - 0xaa
      11'h3F4: dout <= 8'b10101010; // 1012 : 170 - 0xaa
      11'h3F5: dout <= 8'b10101010; // 1013 : 170 - 0xaa
      11'h3F6: dout <= 8'b10101010; // 1014 : 170 - 0xaa
      11'h3F7: dout <= 8'b00100010; // 1015 :  34 - 0x22
      11'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0
      11'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      11'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      11'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      11'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      11'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      11'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      11'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
     //----- Name Table 1---------
      11'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- line 0x0
      11'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      11'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      11'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      11'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      11'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      11'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      11'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      11'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0
      11'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      11'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      11'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      11'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      11'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0
      11'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      11'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      11'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      11'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      11'h415: dout <= 8'b00000000; // 1045 :   0 - 0x0
      11'h416: dout <= 8'b00000000; // 1046 :   0 - 0x0
      11'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      11'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0
      11'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      11'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      11'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- line 0x1
      11'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      11'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      11'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      11'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      11'h425: dout <= 8'b00000000; // 1061 :   0 - 0x0
      11'h426: dout <= 8'b00000000; // 1062 :   0 - 0x0
      11'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      11'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0
      11'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      11'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      11'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      11'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      11'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      11'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      11'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0
      11'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      11'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      11'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      11'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      11'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      11'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      11'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0
      11'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      11'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      11'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      11'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      11'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      11'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      11'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- line 0x2
      11'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      11'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      11'h443: dout <= 8'b00000000; // 1091 :   0 - 0x0
      11'h444: dout <= 8'b00000000; // 1092 :   0 - 0x0
      11'h445: dout <= 8'b00000000; // 1093 :   0 - 0x0
      11'h446: dout <= 8'b00000000; // 1094 :   0 - 0x0
      11'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      11'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0
      11'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      11'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      11'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      11'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      11'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      11'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      11'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0
      11'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      11'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      11'h453: dout <= 8'b00000000; // 1107 :   0 - 0x0
      11'h454: dout <= 8'b00000000; // 1108 :   0 - 0x0
      11'h455: dout <= 8'b00000000; // 1109 :   0 - 0x0
      11'h456: dout <= 8'b00000000; // 1110 :   0 - 0x0
      11'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      11'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0
      11'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      11'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      11'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      11'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      11'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      11'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      11'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- line 0x3
      11'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      11'h464: dout <= 8'b00000000; // 1124 :   0 - 0x0
      11'h465: dout <= 8'b00000000; // 1125 :   0 - 0x0
      11'h466: dout <= 8'b00000000; // 1126 :   0 - 0x0
      11'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      11'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0
      11'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      11'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      11'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      11'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      11'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      11'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      11'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      11'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0
      11'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      11'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      11'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      11'h474: dout <= 8'b00000000; // 1140 :   0 - 0x0
      11'h475: dout <= 8'b00000000; // 1141 :   0 - 0x0
      11'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      11'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      11'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0
      11'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      11'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      11'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      11'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      11'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- line 0x4
      11'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout <= 8'b00000000; // 1156 :   0 - 0x0
      11'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      11'h486: dout <= 8'b00000000; // 1158 :   0 - 0x0
      11'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      11'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0
      11'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      11'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      11'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      11'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      11'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      11'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      11'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0
      11'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      11'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      11'h493: dout <= 8'b00000000; // 1171 :   0 - 0x0
      11'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      11'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      11'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      11'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      11'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0
      11'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      11'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      11'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      11'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      11'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      11'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      11'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- line 0x5
      11'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      11'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      11'h4A4: dout <= 8'b00000000; // 1188 :   0 - 0x0
      11'h4A5: dout <= 8'b00000000; // 1189 :   0 - 0x0
      11'h4A6: dout <= 8'b00000000; // 1190 :   0 - 0x0
      11'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      11'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0
      11'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      11'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      11'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      11'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      11'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      11'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      11'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0
      11'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      11'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      11'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      11'h4B4: dout <= 8'b00000000; // 1204 :   0 - 0x0
      11'h4B5: dout <= 8'b00000000; // 1205 :   0 - 0x0
      11'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      11'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      11'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0
      11'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      11'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      11'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      11'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      11'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      11'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      11'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      11'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- line 0x6
      11'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      11'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout <= 8'b00000000; // 1219 :   0 - 0x0
      11'h4C4: dout <= 8'b00000000; // 1220 :   0 - 0x0
      11'h4C5: dout <= 8'b00000000; // 1221 :   0 - 0x0
      11'h4C6: dout <= 8'b00000000; // 1222 :   0 - 0x0
      11'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      11'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0
      11'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      11'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      11'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      11'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      11'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      11'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      11'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0
      11'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      11'h4D3: dout <= 8'b00000000; // 1235 :   0 - 0x0
      11'h4D4: dout <= 8'b00000000; // 1236 :   0 - 0x0
      11'h4D5: dout <= 8'b00000000; // 1237 :   0 - 0x0
      11'h4D6: dout <= 8'b00000000; // 1238 :   0 - 0x0
      11'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      11'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0
      11'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      11'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      11'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      11'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      11'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      11'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      11'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- line 0x7
      11'h4E1: dout <= 8'b00000000; // 1249 :   0 - 0x0
      11'h4E2: dout <= 8'b00000000; // 1250 :   0 - 0x0
      11'h4E3: dout <= 8'b00000000; // 1251 :   0 - 0x0
      11'h4E4: dout <= 8'b00000000; // 1252 :   0 - 0x0
      11'h4E5: dout <= 8'b00000000; // 1253 :   0 - 0x0
      11'h4E6: dout <= 8'b00000000; // 1254 :   0 - 0x0
      11'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      11'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0
      11'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      11'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      11'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      11'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      11'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      11'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      11'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout <= 8'b00000000; // 1264 :   0 - 0x0
      11'h4F1: dout <= 8'b00000000; // 1265 :   0 - 0x0
      11'h4F2: dout <= 8'b00000000; // 1266 :   0 - 0x0
      11'h4F3: dout <= 8'b00000000; // 1267 :   0 - 0x0
      11'h4F4: dout <= 8'b00000000; // 1268 :   0 - 0x0
      11'h4F5: dout <= 8'b00000000; // 1269 :   0 - 0x0
      11'h4F6: dout <= 8'b00000000; // 1270 :   0 - 0x0
      11'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      11'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0
      11'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      11'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout <= 8'b00000000; // 1280 :   0 - 0x0 -- line 0x8
      11'h501: dout <= 8'b00000000; // 1281 :   0 - 0x0
      11'h502: dout <= 8'b00000000; // 1282 :   0 - 0x0
      11'h503: dout <= 8'b00000000; // 1283 :   0 - 0x0
      11'h504: dout <= 8'b00000000; // 1284 :   0 - 0x0
      11'h505: dout <= 8'b00000000; // 1285 :   0 - 0x0
      11'h506: dout <= 8'b00000000; // 1286 :   0 - 0x0
      11'h507: dout <= 8'b00000000; // 1287 :   0 - 0x0
      11'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0
      11'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      11'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      11'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      11'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      11'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      11'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      11'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      11'h510: dout <= 8'b00000000; // 1296 :   0 - 0x0
      11'h511: dout <= 8'b00000000; // 1297 :   0 - 0x0
      11'h512: dout <= 8'b00000000; // 1298 :   0 - 0x0
      11'h513: dout <= 8'b00000000; // 1299 :   0 - 0x0
      11'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      11'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      11'h516: dout <= 8'b00000000; // 1302 :   0 - 0x0
      11'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0
      11'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      11'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      11'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      11'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      11'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      11'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      11'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      11'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- line 0x9
      11'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      11'h522: dout <= 8'b00000000; // 1314 :   0 - 0x0
      11'h523: dout <= 8'b00000000; // 1315 :   0 - 0x0
      11'h524: dout <= 8'b00000000; // 1316 :   0 - 0x0
      11'h525: dout <= 8'b00000000; // 1317 :   0 - 0x0
      11'h526: dout <= 8'b00000000; // 1318 :   0 - 0x0
      11'h527: dout <= 8'b00000000; // 1319 :   0 - 0x0
      11'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0
      11'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      11'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      11'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      11'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      11'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      11'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      11'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0
      11'h531: dout <= 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout <= 8'b00000000; // 1330 :   0 - 0x0
      11'h533: dout <= 8'b00000000; // 1331 :   0 - 0x0
      11'h534: dout <= 8'b00000000; // 1332 :   0 - 0x0
      11'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      11'h536: dout <= 8'b00000000; // 1334 :   0 - 0x0
      11'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      11'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0
      11'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      11'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      11'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      11'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      11'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      11'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      11'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      11'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- line 0xa
      11'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      11'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      11'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      11'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      11'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      11'h546: dout <= 8'b00000000; // 1350 :   0 - 0x0
      11'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      11'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0
      11'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      11'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      11'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      11'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      11'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      11'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      11'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      11'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0
      11'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      11'h554: dout <= 8'b00000000; // 1364 :   0 - 0x0
      11'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      11'h556: dout <= 8'b00000000; // 1366 :   0 - 0x0
      11'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0
      11'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      11'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- line 0xb
      11'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      11'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      11'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      11'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      11'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0
      11'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      11'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      11'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      11'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      11'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      11'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      11'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      11'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0
      11'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      11'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      11'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      11'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      11'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      11'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0
      11'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      11'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      11'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      11'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      11'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      11'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      11'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- line 0xc
      11'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      11'h582: dout <= 8'b00000000; // 1410 :   0 - 0x0
      11'h583: dout <= 8'b00000000; // 1411 :   0 - 0x0
      11'h584: dout <= 8'b00000000; // 1412 :   0 - 0x0
      11'h585: dout <= 8'b00000000; // 1413 :   0 - 0x0
      11'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      11'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      11'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0
      11'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      11'h58A: dout <= 8'b00000000; // 1418 :   0 - 0x0
      11'h58B: dout <= 8'b00000000; // 1419 :   0 - 0x0
      11'h58C: dout <= 8'b00000000; // 1420 :   0 - 0x0
      11'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      11'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      11'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      11'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0
      11'h591: dout <= 8'b00000000; // 1425 :   0 - 0x0
      11'h592: dout <= 8'b00000000; // 1426 :   0 - 0x0
      11'h593: dout <= 8'b00000000; // 1427 :   0 - 0x0
      11'h594: dout <= 8'b00000000; // 1428 :   0 - 0x0
      11'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      11'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      11'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0
      11'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      11'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      11'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      11'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      11'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      11'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      11'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- line 0xd
      11'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      11'h5A2: dout <= 8'b00000000; // 1442 :   0 - 0x0
      11'h5A3: dout <= 8'b00000000; // 1443 :   0 - 0x0
      11'h5A4: dout <= 8'b00000000; // 1444 :   0 - 0x0
      11'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      11'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      11'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0
      11'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      11'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      11'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      11'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      11'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      11'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      11'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0
      11'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      11'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      11'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      11'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      11'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      11'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      11'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0
      11'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      11'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      11'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      11'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      11'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      11'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      11'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- line 0xe
      11'h5C1: dout <= 8'b00000000; // 1473 :   0 - 0x0
      11'h5C2: dout <= 8'b00000000; // 1474 :   0 - 0x0
      11'h5C3: dout <= 8'b00000000; // 1475 :   0 - 0x0
      11'h5C4: dout <= 8'b00000000; // 1476 :   0 - 0x0
      11'h5C5: dout <= 8'b00000000; // 1477 :   0 - 0x0
      11'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      11'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0
      11'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      11'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      11'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      11'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      11'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      11'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      11'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0
      11'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      11'h5D2: dout <= 8'b00000000; // 1490 :   0 - 0x0
      11'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      11'h5D4: dout <= 8'b00000000; // 1492 :   0 - 0x0
      11'h5D5: dout <= 8'b00000000; // 1493 :   0 - 0x0
      11'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      11'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0
      11'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      11'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      11'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      11'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      11'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- line 0xf
      11'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      11'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      11'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      11'h5E4: dout <= 8'b00000000; // 1508 :   0 - 0x0
      11'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      11'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      11'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0
      11'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      11'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      11'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      11'h5EC: dout <= 8'b00000000; // 1516 :   0 - 0x0
      11'h5ED: dout <= 8'b00000000; // 1517 :   0 - 0x0
      11'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0
      11'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      11'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      11'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      11'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      11'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      11'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      11'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0
      11'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- line 0x10
      11'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      11'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      11'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout <= 8'b00000000; // 1542 :   0 - 0x0
      11'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0
      11'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      11'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0
      11'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      11'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      11'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0
      11'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      11'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      11'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      11'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      11'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      11'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- line 0x11
      11'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0
      11'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      11'h62A: dout <= 8'b00000000; // 1578 :   0 - 0x0
      11'h62B: dout <= 8'b00000000; // 1579 :   0 - 0x0
      11'h62C: dout <= 8'b00000000; // 1580 :   0 - 0x0
      11'h62D: dout <= 8'b00000000; // 1581 :   0 - 0x0
      11'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      11'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0
      11'h631: dout <= 8'b00000000; // 1585 :   0 - 0x0
      11'h632: dout <= 8'b00000000; // 1586 :   0 - 0x0
      11'h633: dout <= 8'b00000000; // 1587 :   0 - 0x0
      11'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      11'h635: dout <= 8'b00000000; // 1589 :   0 - 0x0
      11'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      11'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout <= 8'b00000000; // 1592 :   0 - 0x0
      11'h639: dout <= 8'b00000000; // 1593 :   0 - 0x0
      11'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      11'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      11'h63C: dout <= 8'b00000000; // 1596 :   0 - 0x0
      11'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      11'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      11'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- line 0x12
      11'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0
      11'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      11'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      11'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      11'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      11'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0
      11'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      11'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      11'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      11'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      11'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      11'h656: dout <= 8'b00000000; // 1622 :   0 - 0x0
      11'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      11'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0
      11'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      11'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      11'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      11'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      11'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      11'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- line 0x13
      11'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      11'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      11'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      11'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      11'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0
      11'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      11'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      11'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      11'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      11'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      11'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0
      11'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout <= 8'b00000000; // 1653 :   0 - 0x0
      11'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      11'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      11'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0
      11'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      11'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- line 0x14
      11'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      11'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      11'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      11'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0
      11'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      11'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      11'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      11'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      11'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      11'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0
      11'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      11'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      11'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      11'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      11'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      11'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0
      11'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      11'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      11'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      11'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      11'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      11'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      11'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      11'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- line 0x15
      11'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      11'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      11'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      11'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      11'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0
      11'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      11'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      11'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      11'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      11'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      11'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      11'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      11'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0
      11'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout <= 8'b00000000; // 1715 :   0 - 0x0
      11'h6B4: dout <= 8'b00000000; // 1716 :   0 - 0x0
      11'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      11'h6B6: dout <= 8'b00000000; // 1718 :   0 - 0x0
      11'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      11'h6B8: dout <= 8'b00000000; // 1720 :   0 - 0x0
      11'h6B9: dout <= 8'b00000000; // 1721 :   0 - 0x0
      11'h6BA: dout <= 8'b00000000; // 1722 :   0 - 0x0
      11'h6BB: dout <= 8'b00000000; // 1723 :   0 - 0x0
      11'h6BC: dout <= 8'b00000000; // 1724 :   0 - 0x0
      11'h6BD: dout <= 8'b00000000; // 1725 :   0 - 0x0
      11'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      11'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- line 0x16
      11'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      11'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      11'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      11'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      11'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      11'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0
      11'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      11'h6CA: dout <= 8'b00000000; // 1738 :   0 - 0x0
      11'h6CB: dout <= 8'b00000000; // 1739 :   0 - 0x0
      11'h6CC: dout <= 8'b00000000; // 1740 :   0 - 0x0
      11'h6CD: dout <= 8'b00000000; // 1741 :   0 - 0x0
      11'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      11'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      11'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0
      11'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      11'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      11'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      11'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      11'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      11'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0
      11'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      11'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      11'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      11'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      11'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      11'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      11'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      11'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- line 0x17
      11'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      11'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      11'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      11'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      11'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      11'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0
      11'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      11'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      11'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      11'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      11'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      11'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      11'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout <= 8'b00000000; // 1776 :   0 - 0x0
      11'h6F1: dout <= 8'b00000000; // 1777 :   0 - 0x0
      11'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      11'h6F3: dout <= 8'b00000000; // 1779 :   0 - 0x0
      11'h6F4: dout <= 8'b00000000; // 1780 :   0 - 0x0
      11'h6F5: dout <= 8'b00000000; // 1781 :   0 - 0x0
      11'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      11'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      11'h6F8: dout <= 8'b00000000; // 1784 :   0 - 0x0
      11'h6F9: dout <= 8'b00000000; // 1785 :   0 - 0x0
      11'h6FA: dout <= 8'b00000000; // 1786 :   0 - 0x0
      11'h6FB: dout <= 8'b00000000; // 1787 :   0 - 0x0
      11'h6FC: dout <= 8'b00000000; // 1788 :   0 - 0x0
      11'h6FD: dout <= 8'b00000000; // 1789 :   0 - 0x0
      11'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      11'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      11'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- line 0x18
      11'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      11'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      11'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      11'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      11'h705: dout <= 8'b00000000; // 1797 :   0 - 0x0
      11'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      11'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0
      11'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      11'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      11'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      11'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0
      11'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      11'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      11'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      11'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout <= 8'b00000000; // 1813 :   0 - 0x0
      11'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0
      11'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      11'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      11'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      11'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      11'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      11'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      11'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      11'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- line 0x19
      11'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      11'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      11'h723: dout <= 8'b00000000; // 1827 :   0 - 0x0
      11'h724: dout <= 8'b00000000; // 1828 :   0 - 0x0
      11'h725: dout <= 8'b00000000; // 1829 :   0 - 0x0
      11'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      11'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      11'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0
      11'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      11'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      11'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      11'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      11'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      11'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      11'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      11'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0
      11'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      11'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      11'h735: dout <= 8'b00000000; // 1845 :   0 - 0x0
      11'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      11'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0
      11'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      11'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      11'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      11'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      11'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      11'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      11'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      11'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- line 0x1a
      11'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      11'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0
      11'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      11'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      11'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      11'h74C: dout <= 8'b00000000; // 1868 :   0 - 0x0
      11'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0
      11'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      11'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      11'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0
      11'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      11'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      11'h75B: dout <= 8'b00000000; // 1883 :   0 - 0x0
      11'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      11'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      11'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      11'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- line 0x1b
      11'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      11'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0
      11'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      11'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      11'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      11'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0
      11'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      11'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      11'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0
      11'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      11'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout <= 8'b10100101; // 1920 : 165 - 0xa5 -- line 0x1c
      11'h781: dout <= 8'b10100101; // 1921 : 165 - 0xa5
      11'h782: dout <= 8'b10100101; // 1922 : 165 - 0xa5
      11'h783: dout <= 8'b10100101; // 1923 : 165 - 0xa5
      11'h784: dout <= 8'b10100101; // 1924 : 165 - 0xa5
      11'h785: dout <= 8'b10100101; // 1925 : 165 - 0xa5
      11'h786: dout <= 8'b10100101; // 1926 : 165 - 0xa5
      11'h787: dout <= 8'b10100101; // 1927 : 165 - 0xa5
      11'h788: dout <= 8'b10100101; // 1928 : 165 - 0xa5
      11'h789: dout <= 8'b10100101; // 1929 : 165 - 0xa5
      11'h78A: dout <= 8'b10100101; // 1930 : 165 - 0xa5
      11'h78B: dout <= 8'b10100101; // 1931 : 165 - 0xa5
      11'h78C: dout <= 8'b10100101; // 1932 : 165 - 0xa5
      11'h78D: dout <= 8'b10100101; // 1933 : 165 - 0xa5
      11'h78E: dout <= 8'b10100101; // 1934 : 165 - 0xa5
      11'h78F: dout <= 8'b10100101; // 1935 : 165 - 0xa5
      11'h790: dout <= 8'b10100101; // 1936 : 165 - 0xa5
      11'h791: dout <= 8'b10100101; // 1937 : 165 - 0xa5
      11'h792: dout <= 8'b10100101; // 1938 : 165 - 0xa5
      11'h793: dout <= 8'b10100101; // 1939 : 165 - 0xa5
      11'h794: dout <= 8'b10100101; // 1940 : 165 - 0xa5
      11'h795: dout <= 8'b10100101; // 1941 : 165 - 0xa5
      11'h796: dout <= 8'b10100101; // 1942 : 165 - 0xa5
      11'h797: dout <= 8'b10100101; // 1943 : 165 - 0xa5
      11'h798: dout <= 8'b10100101; // 1944 : 165 - 0xa5
      11'h799: dout <= 8'b10100101; // 1945 : 165 - 0xa5
      11'h79A: dout <= 8'b10100101; // 1946 : 165 - 0xa5
      11'h79B: dout <= 8'b10100101; // 1947 : 165 - 0xa5
      11'h79C: dout <= 8'b10100101; // 1948 : 165 - 0xa5
      11'h79D: dout <= 8'b10100101; // 1949 : 165 - 0xa5
      11'h79E: dout <= 8'b10100101; // 1950 : 165 - 0xa5
      11'h79F: dout <= 8'b10100101; // 1951 : 165 - 0xa5
      11'h7A0: dout <= 8'b10100000; // 1952 : 160 - 0xa0 -- line 0x1d
      11'h7A1: dout <= 8'b10100000; // 1953 : 160 - 0xa0
      11'h7A2: dout <= 8'b10100000; // 1954 : 160 - 0xa0
      11'h7A3: dout <= 8'b10100000; // 1955 : 160 - 0xa0
      11'h7A4: dout <= 8'b10100000; // 1956 : 160 - 0xa0
      11'h7A5: dout <= 8'b10100000; // 1957 : 160 - 0xa0
      11'h7A6: dout <= 8'b10100000; // 1958 : 160 - 0xa0
      11'h7A7: dout <= 8'b10100000; // 1959 : 160 - 0xa0
      11'h7A8: dout <= 8'b10100000; // 1960 : 160 - 0xa0
      11'h7A9: dout <= 8'b10100000; // 1961 : 160 - 0xa0
      11'h7AA: dout <= 8'b10100000; // 1962 : 160 - 0xa0
      11'h7AB: dout <= 8'b10100000; // 1963 : 160 - 0xa0
      11'h7AC: dout <= 8'b10100000; // 1964 : 160 - 0xa0
      11'h7AD: dout <= 8'b10100000; // 1965 : 160 - 0xa0
      11'h7AE: dout <= 8'b10100000; // 1966 : 160 - 0xa0
      11'h7AF: dout <= 8'b10100000; // 1967 : 160 - 0xa0
      11'h7B0: dout <= 8'b10100000; // 1968 : 160 - 0xa0
      11'h7B1: dout <= 8'b10100000; // 1969 : 160 - 0xa0
      11'h7B2: dout <= 8'b10100000; // 1970 : 160 - 0xa0
      11'h7B3: dout <= 8'b10100000; // 1971 : 160 - 0xa0
      11'h7B4: dout <= 8'b10100000; // 1972 : 160 - 0xa0
      11'h7B5: dout <= 8'b10100000; // 1973 : 160 - 0xa0
      11'h7B6: dout <= 8'b10100000; // 1974 : 160 - 0xa0
      11'h7B7: dout <= 8'b10100000; // 1975 : 160 - 0xa0
      11'h7B8: dout <= 8'b10100000; // 1976 : 160 - 0xa0
      11'h7B9: dout <= 8'b10100000; // 1977 : 160 - 0xa0
      11'h7BA: dout <= 8'b10100000; // 1978 : 160 - 0xa0
      11'h7BB: dout <= 8'b10100000; // 1979 : 160 - 0xa0
      11'h7BC: dout <= 8'b10100000; // 1980 : 160 - 0xa0
      11'h7BD: dout <= 8'b10100000; // 1981 : 160 - 0xa0
      11'h7BE: dout <= 8'b10100000; // 1982 : 160 - 0xa0
      11'h7BF: dout <= 8'b10100000; // 1983 : 160 - 0xa0
        //-- Attribute Table 1----
      11'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0
      11'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0
      11'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0
      11'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0
      11'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0
      11'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout <= 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0
      11'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0
      11'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0
      11'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout <= 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout <= 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
