//-   Background Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_PACMAN_BG_PLN0
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 0
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      11'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      11'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      11'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      11'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Background 0x1
      11'h9: dout  = 8'b00111000; //    9 :  56 - 0x38
      11'hA: dout  = 8'b01111100; //   10 : 124 - 0x7c
      11'hB: dout  = 8'b11111110; //   11 : 254 - 0xfe
      11'hC: dout  = 8'b11111110; //   12 : 254 - 0xfe
      11'hD: dout  = 8'b11111110; //   13 : 254 - 0xfe
      11'hE: dout  = 8'b01111100; //   14 : 124 - 0x7c
      11'hF: dout  = 8'b00111000; //   15 :  56 - 0x38
      11'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Background 0x2
      11'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      11'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      11'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      11'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      11'h15: dout  = 8'b00000000; //   21 :   0 - 0x0
      11'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- Background 0x3
      11'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      11'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      11'h1B: dout  = 8'b00011000; //   27 :  24 - 0x18
      11'h1C: dout  = 8'b00011000; //   28 :  24 - 0x18
      11'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      11'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      11'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Background 0x4
      11'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      11'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      11'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      11'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      11'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      11'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout  = 8'b00000000; //   40 :   0 - 0x0 -- Background 0x5
      11'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      11'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      11'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      11'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      11'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Background 0x6
      11'h31: dout  = 8'b00000000; //   49 :   0 - 0x0
      11'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      11'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      11'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      11'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      11'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      11'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout  = 8'b00000000; //   56 :   0 - 0x0 -- Background 0x7
      11'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      11'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      11'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      11'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      11'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Background 0x8
      11'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      11'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      11'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      11'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      11'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Background 0x9
      11'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      11'h4B: dout  = 8'b00011000; //   75 :  24 - 0x18
      11'h4C: dout  = 8'b00011000; //   76 :  24 - 0x18
      11'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      11'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Background 0xa
      11'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      11'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      11'h53: dout  = 8'b00000000; //   83 :   0 - 0x0
      11'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      11'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      11'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- Background 0xb
      11'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      11'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      11'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      11'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      11'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      11'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Background 0xc
      11'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      11'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      11'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      11'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      11'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout  = 8'b00000000; //  104 :   0 - 0x0 -- Background 0xd
      11'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      11'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      11'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      11'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      11'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      11'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Background 0xe
      11'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      11'h72: dout  = 8'b00000000; //  114 :   0 - 0x0
      11'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      11'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      11'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      11'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Background 0xf
      11'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      11'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      11'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      11'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      11'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      11'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      11'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Background 0x10
      11'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      11'h82: dout  = 8'b11111111; //  130 : 255 - 0xff
      11'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      11'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      11'h85: dout  = 8'b11111111; //  133 : 255 - 0xff
      11'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      11'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout  = 8'b00100100; //  136 :  36 - 0x24 -- Background 0x11
      11'h89: dout  = 8'b00100100; //  137 :  36 - 0x24
      11'h8A: dout  = 8'b00100100; //  138 :  36 - 0x24
      11'h8B: dout  = 8'b00100100; //  139 :  36 - 0x24
      11'h8C: dout  = 8'b00100100; //  140 :  36 - 0x24
      11'h8D: dout  = 8'b00100100; //  141 :  36 - 0x24
      11'h8E: dout  = 8'b00100100; //  142 :  36 - 0x24
      11'h8F: dout  = 8'b00100100; //  143 :  36 - 0x24
      11'h90: dout  = 8'b00100100; //  144 :  36 - 0x24 -- Background 0x12
      11'h91: dout  = 8'b00100100; //  145 :  36 - 0x24
      11'h92: dout  = 8'b11000011; //  146 : 195 - 0xc3
      11'h93: dout  = 8'b00000000; //  147 :   0 - 0x0
      11'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      11'h95: dout  = 8'b11111111; //  149 : 255 - 0xff
      11'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- Background 0x13
      11'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      11'h9A: dout  = 8'b11111111; //  154 : 255 - 0xff
      11'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      11'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      11'h9D: dout  = 8'b11000011; //  157 : 195 - 0xc3
      11'h9E: dout  = 8'b00100100; //  158 :  36 - 0x24
      11'h9F: dout  = 8'b00100100; //  159 :  36 - 0x24
      11'hA0: dout  = 8'b00100100; //  160 :  36 - 0x24 -- Background 0x14
      11'hA1: dout  = 8'b00100100; //  161 :  36 - 0x24
      11'hA2: dout  = 8'b11000100; //  162 : 196 - 0xc4
      11'hA3: dout  = 8'b00000100; //  163 :   4 - 0x4
      11'hA4: dout  = 8'b00000100; //  164 :   4 - 0x4
      11'hA5: dout  = 8'b11000100; //  165 : 196 - 0xc4
      11'hA6: dout  = 8'b00100100; //  166 :  36 - 0x24
      11'hA7: dout  = 8'b00100100; //  167 :  36 - 0x24
      11'hA8: dout  = 8'b00100100; //  168 :  36 - 0x24 -- Background 0x15
      11'hA9: dout  = 8'b00100100; //  169 :  36 - 0x24
      11'hAA: dout  = 8'b00100011; //  170 :  35 - 0x23
      11'hAB: dout  = 8'b00100000; //  171 :  32 - 0x20
      11'hAC: dout  = 8'b00100000; //  172 :  32 - 0x20
      11'hAD: dout  = 8'b00100011; //  173 :  35 - 0x23
      11'hAE: dout  = 8'b00100100; //  174 :  36 - 0x24
      11'hAF: dout  = 8'b00100100; //  175 :  36 - 0x24
      11'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Background 0x16
      11'hB1: dout  = 8'b00000000; //  177 :   0 - 0x0
      11'hB2: dout  = 8'b00001111; //  178 :  15 - 0xf
      11'hB3: dout  = 8'b00010000; //  179 :  16 - 0x10
      11'hB4: dout  = 8'b11110000; //  180 : 240 - 0xf0
      11'hB5: dout  = 8'b00001111; //  181 :  15 - 0xf
      11'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      11'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout  = 8'b00000000; //  184 :   0 - 0x0 -- Background 0x17
      11'hB9: dout  = 8'b00000000; //  185 :   0 - 0x0
      11'hBA: dout  = 8'b11110000; //  186 : 240 - 0xf0
      11'hBB: dout  = 8'b00001000; //  187 :   8 - 0x8
      11'hBC: dout  = 8'b00001111; //  188 :  15 - 0xf
      11'hBD: dout  = 8'b11110000; //  189 : 240 - 0xf0
      11'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Background 0x18
      11'hC1: dout  = 8'b00000000; //  193 :   0 - 0x0
      11'hC2: dout  = 8'b11110000; //  194 : 240 - 0xf0
      11'hC3: dout  = 8'b00001000; //  195 :   8 - 0x8
      11'hC4: dout  = 8'b00001000; //  196 :   8 - 0x8
      11'hC5: dout  = 8'b11110000; //  197 : 240 - 0xf0
      11'hC6: dout  = 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- Background 0x19
      11'hC9: dout  = 8'b00000000; //  201 :   0 - 0x0
      11'hCA: dout  = 8'b00001111; //  202 :  15 - 0xf
      11'hCB: dout  = 8'b00010000; //  203 :  16 - 0x10
      11'hCC: dout  = 8'b00010000; //  204 :  16 - 0x10
      11'hCD: dout  = 8'b00001111; //  205 :  15 - 0xf
      11'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout  = 8'b00100100; //  208 :  36 - 0x24 -- Background 0x1a
      11'hD1: dout  = 8'b00100100; //  209 :  36 - 0x24
      11'hD2: dout  = 8'b00100100; //  210 :  36 - 0x24
      11'hD3: dout  = 8'b00100100; //  211 :  36 - 0x24
      11'hD4: dout  = 8'b00011000; //  212 :  24 - 0x18
      11'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      11'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- Background 0x1b
      11'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      11'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      11'hDB: dout  = 8'b00011000; //  219 :  24 - 0x18
      11'hDC: dout  = 8'b00100100; //  220 :  36 - 0x24
      11'hDD: dout  = 8'b00100100; //  221 :  36 - 0x24
      11'hDE: dout  = 8'b00100100; //  222 :  36 - 0x24
      11'hDF: dout  = 8'b00100100; //  223 :  36 - 0x24
      11'hE0: dout  = 8'b00100100; //  224 :  36 - 0x24 -- Background 0x1c
      11'hE1: dout  = 8'b00100100; //  225 :  36 - 0x24
      11'hE2: dout  = 8'b11000100; //  226 : 196 - 0xc4
      11'hE3: dout  = 8'b00000100; //  227 :   4 - 0x4
      11'hE4: dout  = 8'b00001000; //  228 :   8 - 0x8
      11'hE5: dout  = 8'b11110000; //  229 : 240 - 0xf0
      11'hE6: dout  = 8'b00000000; //  230 :   0 - 0x0
      11'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0 -- Background 0x1d
      11'hE9: dout  = 8'b00000000; //  233 :   0 - 0x0
      11'hEA: dout  = 8'b11110000; //  234 : 240 - 0xf0
      11'hEB: dout  = 8'b00001000; //  235 :   8 - 0x8
      11'hEC: dout  = 8'b00000100; //  236 :   4 - 0x4
      11'hED: dout  = 8'b11000100; //  237 : 196 - 0xc4
      11'hEE: dout  = 8'b00100100; //  238 :  36 - 0x24
      11'hEF: dout  = 8'b00100100; //  239 :  36 - 0x24
      11'hF0: dout  = 8'b00100100; //  240 :  36 - 0x24 -- Background 0x1e
      11'hF1: dout  = 8'b00100100; //  241 :  36 - 0x24
      11'hF2: dout  = 8'b00100011; //  242 :  35 - 0x23
      11'hF3: dout  = 8'b00100000; //  243 :  32 - 0x20
      11'hF4: dout  = 8'b00010000; //  244 :  16 - 0x10
      11'hF5: dout  = 8'b00001111; //  245 :  15 - 0xf
      11'hF6: dout  = 8'b00000000; //  246 :   0 - 0x0
      11'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- Background 0x1f
      11'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout  = 8'b00001111; //  250 :  15 - 0xf
      11'hFB: dout  = 8'b00010000; //  251 :  16 - 0x10
      11'hFC: dout  = 8'b00100000; //  252 :  32 - 0x20
      11'hFD: dout  = 8'b00100011; //  253 :  35 - 0x23
      11'hFE: dout  = 8'b00100100; //  254 :  36 - 0x24
      11'hFF: dout  = 8'b00100100; //  255 :  36 - 0x24
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Background 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Background 0x21
      11'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout  = 8'b11110000; //  266 : 240 - 0xf0
      11'h10B: dout  = 8'b00001000; //  267 :   8 - 0x8
      11'h10C: dout  = 8'b00001000; //  268 :   8 - 0x8
      11'h10D: dout  = 8'b11110000; //  269 : 240 - 0xf0
      11'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Background 0x22
      11'h111: dout  = 8'b00000000; //  273 :   0 - 0x0
      11'h112: dout  = 8'b00001111; //  274 :  15 - 0xf
      11'h113: dout  = 8'b00010000; //  275 :  16 - 0x10
      11'h114: dout  = 8'b00010000; //  276 :  16 - 0x10
      11'h115: dout  = 8'b00001111; //  277 :  15 - 0xf
      11'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b11111111; //  280 : 255 - 0xff -- Background 0x23
      11'h119: dout  = 8'b11111111; //  281 : 255 - 0xff
      11'h11A: dout  = 8'b11100001; //  282 : 225 - 0xe1
      11'h11B: dout  = 8'b11100001; //  283 : 225 - 0xe1
      11'h11C: dout  = 8'b11100001; //  284 : 225 - 0xe1
      11'h11D: dout  = 8'b11100001; //  285 : 225 - 0xe1
      11'h11E: dout  = 8'b11100001; //  286 : 225 - 0xe1
      11'h11F: dout  = 8'b11100001; //  287 : 225 - 0xe1
      11'h120: dout  = 8'b10000111; //  288 : 135 - 0x87 -- Background 0x24
      11'h121: dout  = 8'b11000111; //  289 : 199 - 0xc7
      11'h122: dout  = 8'b11000000; //  290 : 192 - 0xc0
      11'h123: dout  = 8'b11000111; //  291 : 199 - 0xc7
      11'h124: dout  = 8'b11001111; //  292 : 207 - 0xcf
      11'h125: dout  = 8'b11001110; //  293 : 206 - 0xce
      11'h126: dout  = 8'b11001111; //  294 : 207 - 0xcf
      11'h127: dout  = 8'b11000111; //  295 : 199 - 0xc7
      11'h128: dout  = 8'b11111000; //  296 : 248 - 0xf8 -- Background 0x25
      11'h129: dout  = 8'b11111100; //  297 : 252 - 0xfc
      11'h12A: dout  = 8'b00011100; //  298 :  28 - 0x1c
      11'h12B: dout  = 8'b11111100; //  299 : 252 - 0xfc
      11'h12C: dout  = 8'b11111100; //  300 : 252 - 0xfc
      11'h12D: dout  = 8'b00011100; //  301 :  28 - 0x1c
      11'h12E: dout  = 8'b11111100; //  302 : 252 - 0xfc
      11'h12F: dout  = 8'b11111100; //  303 : 252 - 0xfc
      11'h130: dout  = 8'b11111111; //  304 : 255 - 0xff -- Background 0x26
      11'h131: dout  = 8'b11111111; //  305 : 255 - 0xff
      11'h132: dout  = 8'b11100111; //  306 : 231 - 0xe7
      11'h133: dout  = 8'b11100111; //  307 : 231 - 0xe7
      11'h134: dout  = 8'b11100111; //  308 : 231 - 0xe7
      11'h135: dout  = 8'b11100111; //  309 : 231 - 0xe7
      11'h136: dout  = 8'b11100111; //  310 : 231 - 0xe7
      11'h137: dout  = 8'b11100111; //  311 : 231 - 0xe7
      11'h138: dout  = 8'b11110000; //  312 : 240 - 0xf0 -- Background 0x27
      11'h139: dout  = 8'b11111001; //  313 : 249 - 0xf9
      11'h13A: dout  = 8'b00111001; //  314 :  57 - 0x39
      11'h13B: dout  = 8'b00111001; //  315 :  57 - 0x39
      11'h13C: dout  = 8'b00111001; //  316 :  57 - 0x39
      11'h13D: dout  = 8'b00111001; //  317 :  57 - 0x39
      11'h13E: dout  = 8'b00111001; //  318 :  57 - 0x39
      11'h13F: dout  = 8'b00111000; //  319 :  56 - 0x38
      11'h140: dout  = 8'b11111111; //  320 : 255 - 0xff -- Background 0x28
      11'h141: dout  = 8'b11111111; //  321 : 255 - 0xff
      11'h142: dout  = 8'b11000000; //  322 : 192 - 0xc0
      11'h143: dout  = 8'b11000000; //  323 : 192 - 0xc0
      11'h144: dout  = 8'b11000000; //  324 : 192 - 0xc0
      11'h145: dout  = 8'b11000000; //  325 : 192 - 0xc0
      11'h146: dout  = 8'b11111111; //  326 : 255 - 0xff
      11'h147: dout  = 8'b11111111; //  327 : 255 - 0xff
      11'h148: dout  = 8'b00011111; //  328 :  31 - 0x1f -- Background 0x29
      11'h149: dout  = 8'b00111111; //  329 :  63 - 0x3f
      11'h14A: dout  = 8'b00110000; //  330 :  48 - 0x30
      11'h14B: dout  = 8'b00110000; //  331 :  48 - 0x30
      11'h14C: dout  = 8'b00110000; //  332 :  48 - 0x30
      11'h14D: dout  = 8'b00110000; //  333 :  48 - 0x30
      11'h14E: dout  = 8'b00111111; //  334 :  63 - 0x3f
      11'h14F: dout  = 8'b00011111; //  335 :  31 - 0x1f
      11'h150: dout  = 8'b11100011; //  336 : 227 - 0xe3 -- Background 0x2a
      11'h151: dout  = 8'b11110011; //  337 : 243 - 0xf3
      11'h152: dout  = 8'b01110000; //  338 : 112 - 0x70
      11'h153: dout  = 8'b01110000; //  339 : 112 - 0x70
      11'h154: dout  = 8'b01110000; //  340 : 112 - 0x70
      11'h155: dout  = 8'b01110000; //  341 : 112 - 0x70
      11'h156: dout  = 8'b11110000; //  342 : 240 - 0xf0
      11'h157: dout  = 8'b11100000; //  343 : 224 - 0xe0
      11'h158: dout  = 8'b11111110; //  344 : 254 - 0xfe -- Background 0x2b
      11'h159: dout  = 8'b11111110; //  345 : 254 - 0xfe
      11'h15A: dout  = 8'b01110000; //  346 : 112 - 0x70
      11'h15B: dout  = 8'b01110000; //  347 : 112 - 0x70
      11'h15C: dout  = 8'b01110000; //  348 : 112 - 0x70
      11'h15D: dout  = 8'b01110000; //  349 : 112 - 0x70
      11'h15E: dout  = 8'b01110000; //  350 : 112 - 0x70
      11'h15F: dout  = 8'b01110000; //  351 : 112 - 0x70
      11'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Background 0x2c
      11'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout  = 8'b11111111; //  356 : 255 - 0xff
      11'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Background 0x2d
      11'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout  = 8'b00000000; //  362 :   0 - 0x0
      11'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      11'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      11'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Background 0x2e
      11'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout  = 8'b00011000; //  371 :  24 - 0x18
      11'h174: dout  = 8'b00011000; //  372 :  24 - 0x18
      11'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b00000000; //  376 :   0 - 0x0 -- Background 0x2f
      11'h179: dout  = 8'b00000000; //  377 :   0 - 0x0
      11'h17A: dout  = 8'b00000000; //  378 :   0 - 0x0
      11'h17B: dout  = 8'b00000000; //  379 :   0 - 0x0
      11'h17C: dout  = 8'b00000000; //  380 :   0 - 0x0
      11'h17D: dout  = 8'b00000000; //  381 :   0 - 0x0
      11'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      11'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout  = 8'b00011100; //  384 :  28 - 0x1c -- Background 0x30
      11'h181: dout  = 8'b00100110; //  385 :  38 - 0x26
      11'h182: dout  = 8'b01100011; //  386 :  99 - 0x63
      11'h183: dout  = 8'b01100011; //  387 :  99 - 0x63
      11'h184: dout  = 8'b01100011; //  388 :  99 - 0x63
      11'h185: dout  = 8'b00110010; //  389 :  50 - 0x32
      11'h186: dout  = 8'b00011100; //  390 :  28 - 0x1c
      11'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout  = 8'b00001100; //  392 :  12 - 0xc -- Background 0x31
      11'h189: dout  = 8'b00011100; //  393 :  28 - 0x1c
      11'h18A: dout  = 8'b00001100; //  394 :  12 - 0xc
      11'h18B: dout  = 8'b00001100; //  395 :  12 - 0xc
      11'h18C: dout  = 8'b00001100; //  396 :  12 - 0xc
      11'h18D: dout  = 8'b00001100; //  397 :  12 - 0xc
      11'h18E: dout  = 8'b00111111; //  398 :  63 - 0x3f
      11'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout  = 8'b00111110; //  400 :  62 - 0x3e -- Background 0x32
      11'h191: dout  = 8'b01100011; //  401 :  99 - 0x63
      11'h192: dout  = 8'b00000111; //  402 :   7 - 0x7
      11'h193: dout  = 8'b00011110; //  403 :  30 - 0x1e
      11'h194: dout  = 8'b00111100; //  404 :  60 - 0x3c
      11'h195: dout  = 8'b01110000; //  405 : 112 - 0x70
      11'h196: dout  = 8'b01111111; //  406 : 127 - 0x7f
      11'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      11'h198: dout  = 8'b00111111; //  408 :  63 - 0x3f -- Background 0x33
      11'h199: dout  = 8'b00000110; //  409 :   6 - 0x6
      11'h19A: dout  = 8'b00001100; //  410 :  12 - 0xc
      11'h19B: dout  = 8'b00011110; //  411 :  30 - 0x1e
      11'h19C: dout  = 8'b00000011; //  412 :   3 - 0x3
      11'h19D: dout  = 8'b01100011; //  413 :  99 - 0x63
      11'h19E: dout  = 8'b00111110; //  414 :  62 - 0x3e
      11'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout  = 8'b00001110; //  416 :  14 - 0xe -- Background 0x34
      11'h1A1: dout  = 8'b00011110; //  417 :  30 - 0x1e
      11'h1A2: dout  = 8'b00110110; //  418 :  54 - 0x36
      11'h1A3: dout  = 8'b01100110; //  419 : 102 - 0x66
      11'h1A4: dout  = 8'b01111111; //  420 : 127 - 0x7f
      11'h1A5: dout  = 8'b00000110; //  421 :   6 - 0x6
      11'h1A6: dout  = 8'b00000110; //  422 :   6 - 0x6
      11'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      11'h1A8: dout  = 8'b01111110; //  424 : 126 - 0x7e -- Background 0x35
      11'h1A9: dout  = 8'b01100000; //  425 :  96 - 0x60
      11'h1AA: dout  = 8'b01111110; //  426 : 126 - 0x7e
      11'h1AB: dout  = 8'b00000011; //  427 :   3 - 0x3
      11'h1AC: dout  = 8'b00000011; //  428 :   3 - 0x3
      11'h1AD: dout  = 8'b01100011; //  429 :  99 - 0x63
      11'h1AE: dout  = 8'b00111110; //  430 :  62 - 0x3e
      11'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout  = 8'b00011110; //  432 :  30 - 0x1e -- Background 0x36
      11'h1B1: dout  = 8'b00110000; //  433 :  48 - 0x30
      11'h1B2: dout  = 8'b01100000; //  434 :  96 - 0x60
      11'h1B3: dout  = 8'b01111110; //  435 : 126 - 0x7e
      11'h1B4: dout  = 8'b01100011; //  436 :  99 - 0x63
      11'h1B5: dout  = 8'b01100011; //  437 :  99 - 0x63
      11'h1B6: dout  = 8'b00111110; //  438 :  62 - 0x3e
      11'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout  = 8'b01111111; //  440 : 127 - 0x7f -- Background 0x37
      11'h1B9: dout  = 8'b01100011; //  441 :  99 - 0x63
      11'h1BA: dout  = 8'b00000110; //  442 :   6 - 0x6
      11'h1BB: dout  = 8'b00001100; //  443 :  12 - 0xc
      11'h1BC: dout  = 8'b00011000; //  444 :  24 - 0x18
      11'h1BD: dout  = 8'b00011000; //  445 :  24 - 0x18
      11'h1BE: dout  = 8'b00011000; //  446 :  24 - 0x18
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b00111100; //  448 :  60 - 0x3c -- Background 0x38
      11'h1C1: dout  = 8'b01100010; //  449 :  98 - 0x62
      11'h1C2: dout  = 8'b01110010; //  450 : 114 - 0x72
      11'h1C3: dout  = 8'b00111100; //  451 :  60 - 0x3c
      11'h1C4: dout  = 8'b01001111; //  452 :  79 - 0x4f
      11'h1C5: dout  = 8'b01000011; //  453 :  67 - 0x43
      11'h1C6: dout  = 8'b00111110; //  454 :  62 - 0x3e
      11'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout  = 8'b00111110; //  456 :  62 - 0x3e -- Background 0x39
      11'h1C9: dout  = 8'b01100011; //  457 :  99 - 0x63
      11'h1CA: dout  = 8'b01100011; //  458 :  99 - 0x63
      11'h1CB: dout  = 8'b00111111; //  459 :  63 - 0x3f
      11'h1CC: dout  = 8'b00000011; //  460 :   3 - 0x3
      11'h1CD: dout  = 8'b00000110; //  461 :   6 - 0x6
      11'h1CE: dout  = 8'b00111100; //  462 :  60 - 0x3c
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout  = 8'b01111110; //  467 : 126 - 0x7e
      11'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Background 0x3b
      11'h1D9: dout  = 8'b00000010; //  473 :   2 - 0x2
      11'h1DA: dout  = 8'b00000100; //  474 :   4 - 0x4
      11'h1DB: dout  = 8'b00001000; //  475 :   8 - 0x8
      11'h1DC: dout  = 8'b00010000; //  476 :  16 - 0x10
      11'h1DD: dout  = 8'b00100000; //  477 :  32 - 0x20
      11'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Background 0x3c
      11'h1E1: dout  = 8'b00000111; //  481 :   7 - 0x7
      11'h1E2: dout  = 8'b00011111; //  482 :  31 - 0x1f
      11'h1E3: dout  = 8'b00111111; //  483 :  63 - 0x3f
      11'h1E4: dout  = 8'b00111111; //  484 :  63 - 0x3f
      11'h1E5: dout  = 8'b00001111; //  485 :  15 - 0xf
      11'h1E6: dout  = 8'b00000011; //  486 :   3 - 0x3
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Background 0x3d
      11'h1E9: dout  = 8'b11000000; //  489 : 192 - 0xc0
      11'h1EA: dout  = 8'b11110000; //  490 : 240 - 0xf0
      11'h1EB: dout  = 8'b11111000; //  491 : 248 - 0xf8
      11'h1EC: dout  = 8'b11111000; //  492 : 248 - 0xf8
      11'h1ED: dout  = 8'b11111100; //  493 : 252 - 0xfc
      11'h1EE: dout  = 8'b11111100; //  494 : 252 - 0xfc
      11'h1EF: dout  = 8'b11111100; //  495 : 252 - 0xfc
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout  = 8'b00000011; //  497 :   3 - 0x3
      11'h1F2: dout  = 8'b00001111; //  498 :  15 - 0xf
      11'h1F3: dout  = 8'b00111111; //  499 :  63 - 0x3f
      11'h1F4: dout  = 8'b00111111; //  500 :  63 - 0x3f
      11'h1F5: dout  = 8'b00011111; //  501 :  31 - 0x1f
      11'h1F6: dout  = 8'b00000111; //  502 :   7 - 0x7
      11'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout  = 8'b11111100; //  504 : 252 - 0xfc -- Background 0x3f
      11'h1F9: dout  = 8'b11111100; //  505 : 252 - 0xfc
      11'h1FA: dout  = 8'b11111100; //  506 : 252 - 0xfc
      11'h1FB: dout  = 8'b11111000; //  507 : 248 - 0xf8
      11'h1FC: dout  = 8'b11111000; //  508 : 248 - 0xf8
      11'h1FD: dout  = 8'b11110000; //  509 : 240 - 0xf0
      11'h1FE: dout  = 8'b11000000; //  510 : 192 - 0xc0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Background 0x40
      11'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      11'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      11'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00011100; //  520 :  28 - 0x1c -- Background 0x41
      11'h209: dout  = 8'b00110110; //  521 :  54 - 0x36
      11'h20A: dout  = 8'b01100011; //  522 :  99 - 0x63
      11'h20B: dout  = 8'b01100011; //  523 :  99 - 0x63
      11'h20C: dout  = 8'b01111111; //  524 : 127 - 0x7f
      11'h20D: dout  = 8'b01100011; //  525 :  99 - 0x63
      11'h20E: dout  = 8'b01100011; //  526 :  99 - 0x63
      11'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout  = 8'b01111110; //  528 : 126 - 0x7e -- Background 0x42
      11'h211: dout  = 8'b01100011; //  529 :  99 - 0x63
      11'h212: dout  = 8'b01100011; //  530 :  99 - 0x63
      11'h213: dout  = 8'b01111110; //  531 : 126 - 0x7e
      11'h214: dout  = 8'b01100011; //  532 :  99 - 0x63
      11'h215: dout  = 8'b01100011; //  533 :  99 - 0x63
      11'h216: dout  = 8'b01111110; //  534 : 126 - 0x7e
      11'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout  = 8'b00011110; //  536 :  30 - 0x1e -- Background 0x43
      11'h219: dout  = 8'b00110011; //  537 :  51 - 0x33
      11'h21A: dout  = 8'b01100000; //  538 :  96 - 0x60
      11'h21B: dout  = 8'b01100000; //  539 :  96 - 0x60
      11'h21C: dout  = 8'b01100000; //  540 :  96 - 0x60
      11'h21D: dout  = 8'b00110011; //  541 :  51 - 0x33
      11'h21E: dout  = 8'b00011110; //  542 :  30 - 0x1e
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b01111100; //  544 : 124 - 0x7c -- Background 0x44
      11'h221: dout  = 8'b01100110; //  545 : 102 - 0x66
      11'h222: dout  = 8'b01100011; //  546 :  99 - 0x63
      11'h223: dout  = 8'b01100011; //  547 :  99 - 0x63
      11'h224: dout  = 8'b01100011; //  548 :  99 - 0x63
      11'h225: dout  = 8'b01100110; //  549 : 102 - 0x66
      11'h226: dout  = 8'b01111100; //  550 : 124 - 0x7c
      11'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout  = 8'b01111111; //  552 : 127 - 0x7f -- Background 0x45
      11'h229: dout  = 8'b01100000; //  553 :  96 - 0x60
      11'h22A: dout  = 8'b01100000; //  554 :  96 - 0x60
      11'h22B: dout  = 8'b01111110; //  555 : 126 - 0x7e
      11'h22C: dout  = 8'b01100000; //  556 :  96 - 0x60
      11'h22D: dout  = 8'b01100000; //  557 :  96 - 0x60
      11'h22E: dout  = 8'b01111111; //  558 : 127 - 0x7f
      11'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout  = 8'b01111111; //  560 : 127 - 0x7f -- Background 0x46
      11'h231: dout  = 8'b01100000; //  561 :  96 - 0x60
      11'h232: dout  = 8'b01100000; //  562 :  96 - 0x60
      11'h233: dout  = 8'b01111110; //  563 : 126 - 0x7e
      11'h234: dout  = 8'b01100000; //  564 :  96 - 0x60
      11'h235: dout  = 8'b01100000; //  565 :  96 - 0x60
      11'h236: dout  = 8'b01100000; //  566 :  96 - 0x60
      11'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout  = 8'b00011111; //  568 :  31 - 0x1f -- Background 0x47
      11'h239: dout  = 8'b00110000; //  569 :  48 - 0x30
      11'h23A: dout  = 8'b01100000; //  570 :  96 - 0x60
      11'h23B: dout  = 8'b01100111; //  571 : 103 - 0x67
      11'h23C: dout  = 8'b01100011; //  572 :  99 - 0x63
      11'h23D: dout  = 8'b00110011; //  573 :  51 - 0x33
      11'h23E: dout  = 8'b00011111; //  574 :  31 - 0x1f
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b01100011; //  576 :  99 - 0x63 -- Background 0x48
      11'h241: dout  = 8'b01100011; //  577 :  99 - 0x63
      11'h242: dout  = 8'b01100011; //  578 :  99 - 0x63
      11'h243: dout  = 8'b01111111; //  579 : 127 - 0x7f
      11'h244: dout  = 8'b01100011; //  580 :  99 - 0x63
      11'h245: dout  = 8'b01100011; //  581 :  99 - 0x63
      11'h246: dout  = 8'b01100011; //  582 :  99 - 0x63
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b00111111; //  584 :  63 - 0x3f -- Background 0x49
      11'h249: dout  = 8'b00001100; //  585 :  12 - 0xc
      11'h24A: dout  = 8'b00001100; //  586 :  12 - 0xc
      11'h24B: dout  = 8'b00001100; //  587 :  12 - 0xc
      11'h24C: dout  = 8'b00001100; //  588 :  12 - 0xc
      11'h24D: dout  = 8'b00001100; //  589 :  12 - 0xc
      11'h24E: dout  = 8'b00111111; //  590 :  63 - 0x3f
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b00000011; //  592 :   3 - 0x3 -- Background 0x4a
      11'h251: dout  = 8'b00000011; //  593 :   3 - 0x3
      11'h252: dout  = 8'b00000011; //  594 :   3 - 0x3
      11'h253: dout  = 8'b00000011; //  595 :   3 - 0x3
      11'h254: dout  = 8'b00000011; //  596 :   3 - 0x3
      11'h255: dout  = 8'b01100011; //  597 :  99 - 0x63
      11'h256: dout  = 8'b00111110; //  598 :  62 - 0x3e
      11'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout  = 8'b01100011; //  600 :  99 - 0x63 -- Background 0x4b
      11'h259: dout  = 8'b01100110; //  601 : 102 - 0x66
      11'h25A: dout  = 8'b01101100; //  602 : 108 - 0x6c
      11'h25B: dout  = 8'b01111000; //  603 : 120 - 0x78
      11'h25C: dout  = 8'b01111100; //  604 : 124 - 0x7c
      11'h25D: dout  = 8'b01100110; //  605 : 102 - 0x66
      11'h25E: dout  = 8'b01100011; //  606 :  99 - 0x63
      11'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout  = 8'b01100000; //  608 :  96 - 0x60 -- Background 0x4c
      11'h261: dout  = 8'b01100000; //  609 :  96 - 0x60
      11'h262: dout  = 8'b01100000; //  610 :  96 - 0x60
      11'h263: dout  = 8'b01100000; //  611 :  96 - 0x60
      11'h264: dout  = 8'b01100000; //  612 :  96 - 0x60
      11'h265: dout  = 8'b01100000; //  613 :  96 - 0x60
      11'h266: dout  = 8'b01111111; //  614 : 127 - 0x7f
      11'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      11'h268: dout  = 8'b01100011; //  616 :  99 - 0x63 -- Background 0x4d
      11'h269: dout  = 8'b01110111; //  617 : 119 - 0x77
      11'h26A: dout  = 8'b01111111; //  618 : 127 - 0x7f
      11'h26B: dout  = 8'b01111111; //  619 : 127 - 0x7f
      11'h26C: dout  = 8'b01101011; //  620 : 107 - 0x6b
      11'h26D: dout  = 8'b01100011; //  621 :  99 - 0x63
      11'h26E: dout  = 8'b01100011; //  622 :  99 - 0x63
      11'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout  = 8'b01100011; //  624 :  99 - 0x63 -- Background 0x4e
      11'h271: dout  = 8'b01110011; //  625 : 115 - 0x73
      11'h272: dout  = 8'b01111011; //  626 : 123 - 0x7b
      11'h273: dout  = 8'b01111111; //  627 : 127 - 0x7f
      11'h274: dout  = 8'b01101111; //  628 : 111 - 0x6f
      11'h275: dout  = 8'b01100111; //  629 : 103 - 0x67
      11'h276: dout  = 8'b01100011; //  630 :  99 - 0x63
      11'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      11'h278: dout  = 8'b00111110; //  632 :  62 - 0x3e -- Background 0x4f
      11'h279: dout  = 8'b01100011; //  633 :  99 - 0x63
      11'h27A: dout  = 8'b01100011; //  634 :  99 - 0x63
      11'h27B: dout  = 8'b01100011; //  635 :  99 - 0x63
      11'h27C: dout  = 8'b01100011; //  636 :  99 - 0x63
      11'h27D: dout  = 8'b01100011; //  637 :  99 - 0x63
      11'h27E: dout  = 8'b00111110; //  638 :  62 - 0x3e
      11'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      11'h280: dout  = 8'b01111110; //  640 : 126 - 0x7e -- Background 0x50
      11'h281: dout  = 8'b01100011; //  641 :  99 - 0x63
      11'h282: dout  = 8'b01100011; //  642 :  99 - 0x63
      11'h283: dout  = 8'b01100011; //  643 :  99 - 0x63
      11'h284: dout  = 8'b01111110; //  644 : 126 - 0x7e
      11'h285: dout  = 8'b01100000; //  645 :  96 - 0x60
      11'h286: dout  = 8'b01100000; //  646 :  96 - 0x60
      11'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      11'h288: dout  = 8'b00111110; //  648 :  62 - 0x3e -- Background 0x51
      11'h289: dout  = 8'b01100011; //  649 :  99 - 0x63
      11'h28A: dout  = 8'b01100011; //  650 :  99 - 0x63
      11'h28B: dout  = 8'b01100011; //  651 :  99 - 0x63
      11'h28C: dout  = 8'b01101111; //  652 : 111 - 0x6f
      11'h28D: dout  = 8'b01100110; //  653 : 102 - 0x66
      11'h28E: dout  = 8'b00111101; //  654 :  61 - 0x3d
      11'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      11'h290: dout  = 8'b01111110; //  656 : 126 - 0x7e -- Background 0x52
      11'h291: dout  = 8'b01100011; //  657 :  99 - 0x63
      11'h292: dout  = 8'b01100011; //  658 :  99 - 0x63
      11'h293: dout  = 8'b01100111; //  659 : 103 - 0x67
      11'h294: dout  = 8'b01111100; //  660 : 124 - 0x7c
      11'h295: dout  = 8'b01101110; //  661 : 110 - 0x6e
      11'h296: dout  = 8'b01100111; //  662 : 103 - 0x67
      11'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      11'h298: dout  = 8'b00111100; //  664 :  60 - 0x3c -- Background 0x53
      11'h299: dout  = 8'b01100110; //  665 : 102 - 0x66
      11'h29A: dout  = 8'b01100000; //  666 :  96 - 0x60
      11'h29B: dout  = 8'b00111110; //  667 :  62 - 0x3e
      11'h29C: dout  = 8'b00000011; //  668 :   3 - 0x3
      11'h29D: dout  = 8'b01100011; //  669 :  99 - 0x63
      11'h29E: dout  = 8'b00111110; //  670 :  62 - 0x3e
      11'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout  = 8'b00111111; //  672 :  63 - 0x3f -- Background 0x54
      11'h2A1: dout  = 8'b00001100; //  673 :  12 - 0xc
      11'h2A2: dout  = 8'b00001100; //  674 :  12 - 0xc
      11'h2A3: dout  = 8'b00001100; //  675 :  12 - 0xc
      11'h2A4: dout  = 8'b00001100; //  676 :  12 - 0xc
      11'h2A5: dout  = 8'b00001100; //  677 :  12 - 0xc
      11'h2A6: dout  = 8'b00001100; //  678 :  12 - 0xc
      11'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      11'h2A8: dout  = 8'b01100011; //  680 :  99 - 0x63 -- Background 0x55
      11'h2A9: dout  = 8'b01100011; //  681 :  99 - 0x63
      11'h2AA: dout  = 8'b01100011; //  682 :  99 - 0x63
      11'h2AB: dout  = 8'b01100011; //  683 :  99 - 0x63
      11'h2AC: dout  = 8'b01100011; //  684 :  99 - 0x63
      11'h2AD: dout  = 8'b01100011; //  685 :  99 - 0x63
      11'h2AE: dout  = 8'b00111110; //  686 :  62 - 0x3e
      11'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      11'h2B0: dout  = 8'b01100011; //  688 :  99 - 0x63 -- Background 0x56
      11'h2B1: dout  = 8'b01100011; //  689 :  99 - 0x63
      11'h2B2: dout  = 8'b01100011; //  690 :  99 - 0x63
      11'h2B3: dout  = 8'b01110111; //  691 : 119 - 0x77
      11'h2B4: dout  = 8'b00111110; //  692 :  62 - 0x3e
      11'h2B5: dout  = 8'b00011100; //  693 :  28 - 0x1c
      11'h2B6: dout  = 8'b00001000; //  694 :   8 - 0x8
      11'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout  = 8'b01100011; //  696 :  99 - 0x63 -- Background 0x57
      11'h2B9: dout  = 8'b01100011; //  697 :  99 - 0x63
      11'h2BA: dout  = 8'b01101011; //  698 : 107 - 0x6b
      11'h2BB: dout  = 8'b01111111; //  699 : 127 - 0x7f
      11'h2BC: dout  = 8'b01111111; //  700 : 127 - 0x7f
      11'h2BD: dout  = 8'b01110111; //  701 : 119 - 0x77
      11'h2BE: dout  = 8'b01100011; //  702 :  99 - 0x63
      11'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout  = 8'b01100011; //  704 :  99 - 0x63 -- Background 0x58
      11'h2C1: dout  = 8'b01110111; //  705 : 119 - 0x77
      11'h2C2: dout  = 8'b00111110; //  706 :  62 - 0x3e
      11'h2C3: dout  = 8'b00011100; //  707 :  28 - 0x1c
      11'h2C4: dout  = 8'b00111110; //  708 :  62 - 0x3e
      11'h2C5: dout  = 8'b01110111; //  709 : 119 - 0x77
      11'h2C6: dout  = 8'b01100011; //  710 :  99 - 0x63
      11'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      11'h2C8: dout  = 8'b00110011; //  712 :  51 - 0x33 -- Background 0x59
      11'h2C9: dout  = 8'b00110011; //  713 :  51 - 0x33
      11'h2CA: dout  = 8'b00110011; //  714 :  51 - 0x33
      11'h2CB: dout  = 8'b00011110; //  715 :  30 - 0x1e
      11'h2CC: dout  = 8'b00001100; //  716 :  12 - 0xc
      11'h2CD: dout  = 8'b00001100; //  717 :  12 - 0xc
      11'h2CE: dout  = 8'b00001100; //  718 :  12 - 0xc
      11'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      11'h2D0: dout  = 8'b01111111; //  720 : 127 - 0x7f -- Background 0x5a
      11'h2D1: dout  = 8'b00000111; //  721 :   7 - 0x7
      11'h2D2: dout  = 8'b00001110; //  722 :  14 - 0xe
      11'h2D3: dout  = 8'b00011100; //  723 :  28 - 0x1c
      11'h2D4: dout  = 8'b00111000; //  724 :  56 - 0x38
      11'h2D5: dout  = 8'b01110000; //  725 : 112 - 0x70
      11'h2D6: dout  = 8'b01111111; //  726 : 127 - 0x7f
      11'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Background 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      11'h2DD: dout  = 8'b00110000; //  733 :  48 - 0x30
      11'h2DE: dout  = 8'b00110000; //  734 :  48 - 0x30
      11'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      11'h2E0: dout  = 8'b11000000; //  736 : 192 - 0xc0 -- Background 0x5c
      11'h2E1: dout  = 8'b11110000; //  737 : 240 - 0xf0
      11'h2E2: dout  = 8'b11111100; //  738 : 252 - 0xfc
      11'h2E3: dout  = 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout  = 8'b11111100; //  740 : 252 - 0xfc
      11'h2E5: dout  = 8'b11110000; //  741 : 240 - 0xf0
      11'h2E6: dout  = 8'b11000000; //  742 : 192 - 0xc0
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b00111100; //  744 :  60 - 0x3c -- Background 0x5d
      11'h2E9: dout  = 8'b01000010; //  745 :  66 - 0x42
      11'h2EA: dout  = 8'b10011001; //  746 : 153 - 0x99
      11'h2EB: dout  = 8'b10100001; //  747 : 161 - 0xa1
      11'h2EC: dout  = 8'b10100001; //  748 : 161 - 0xa1
      11'h2ED: dout  = 8'b10011001; //  749 : 153 - 0x99
      11'h2EE: dout  = 8'b01000010; //  750 :  66 - 0x42
      11'h2EF: dout  = 8'b00111100; //  751 :  60 - 0x3c
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Background 0x5e
      11'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      11'h2F2: dout  = 8'b00010000; //  754 :  16 - 0x10
      11'h2F3: dout  = 8'b00010000; //  755 :  16 - 0x10
      11'h2F4: dout  = 8'b00010000; //  756 :  16 - 0x10
      11'h2F5: dout  = 8'b00010000; //  757 :  16 - 0x10
      11'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b00110110; //  760 :  54 - 0x36 -- Background 0x5f
      11'h2F9: dout  = 8'b00110110; //  761 :  54 - 0x36
      11'h2FA: dout  = 8'b00010010; //  762 :  18 - 0x12
      11'h2FB: dout  = 8'b00000000; //  763 :   0 - 0x0
      11'h2FC: dout  = 8'b00000000; //  764 :   0 - 0x0
      11'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      11'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      11'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      11'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Background 0x60
      11'h301: dout  = 8'b00000000; //  769 :   0 - 0x0
      11'h302: dout  = 8'b00000000; //  770 :   0 - 0x0
      11'h303: dout  = 8'b00000000; //  771 :   0 - 0x0
      11'h304: dout  = 8'b00000000; //  772 :   0 - 0x0
      11'h305: dout  = 8'b00000001; //  773 :   1 - 0x1
      11'h306: dout  = 8'b00011110; //  774 :  30 - 0x1e
      11'h307: dout  = 8'b00111011; //  775 :  59 - 0x3b
      11'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Background 0x61
      11'h309: dout  = 8'b00000000; //  777 :   0 - 0x0
      11'h30A: dout  = 8'b00001100; //  778 :  12 - 0xc
      11'h30B: dout  = 8'b00111100; //  779 :  60 - 0x3c
      11'h30C: dout  = 8'b11010000; //  780 : 208 - 0xd0
      11'h30D: dout  = 8'b00010000; //  781 :  16 - 0x10
      11'h30E: dout  = 8'b00100000; //  782 :  32 - 0x20
      11'h30F: dout  = 8'b01000000; //  783 :  64 - 0x40
      11'h310: dout  = 8'b00111110; //  784 :  62 - 0x3e -- Background 0x62
      11'h311: dout  = 8'b00101101; //  785 :  45 - 0x2d
      11'h312: dout  = 8'b00110101; //  786 :  53 - 0x35
      11'h313: dout  = 8'b00011101; //  787 :  29 - 0x1d
      11'h314: dout  = 8'b00000001; //  788 :   1 - 0x1
      11'h315: dout  = 8'b00000000; //  789 :   0 - 0x0
      11'h316: dout  = 8'b00000000; //  790 :   0 - 0x0
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b10110000; //  792 : 176 - 0xb0 -- Background 0x63
      11'h319: dout  = 8'b10111000; //  793 : 184 - 0xb8
      11'h31A: dout  = 8'b11111000; //  794 : 248 - 0xf8
      11'h31B: dout  = 8'b01111000; //  795 : 120 - 0x78
      11'h31C: dout  = 8'b10011000; //  796 : 152 - 0x98
      11'h31D: dout  = 8'b11110000; //  797 : 240 - 0xf0
      11'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      11'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Background 0x64
      11'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      11'h322: dout  = 8'b00000111; //  802 :   7 - 0x7
      11'h323: dout  = 8'b00000011; //  803 :   3 - 0x3
      11'h324: dout  = 8'b00001101; //  804 :  13 - 0xd
      11'h325: dout  = 8'b00011110; //  805 :  30 - 0x1e
      11'h326: dout  = 8'b00010111; //  806 :  23 - 0x17
      11'h327: dout  = 8'b00011101; //  807 :  29 - 0x1d
      11'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Background 0x65
      11'h329: dout  = 8'b10000000; //  809 : 128 - 0x80
      11'h32A: dout  = 8'b01110000; //  810 : 112 - 0x70
      11'h32B: dout  = 8'b11100000; //  811 : 224 - 0xe0
      11'h32C: dout  = 8'b11011000; //  812 : 216 - 0xd8
      11'h32D: dout  = 8'b10111100; //  813 : 188 - 0xbc
      11'h32E: dout  = 8'b01110100; //  814 : 116 - 0x74
      11'h32F: dout  = 8'b11011100; //  815 : 220 - 0xdc
      11'h330: dout  = 8'b00011111; //  816 :  31 - 0x1f -- Background 0x66
      11'h331: dout  = 8'b00001011; //  817 :  11 - 0xb
      11'h332: dout  = 8'b00001111; //  818 :  15 - 0xf
      11'h333: dout  = 8'b00000101; //  819 :   5 - 0x5
      11'h334: dout  = 8'b00000011; //  820 :   3 - 0x3
      11'h335: dout  = 8'b00000001; //  821 :   1 - 0x1
      11'h336: dout  = 8'b00000000; //  822 :   0 - 0x0
      11'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      11'h338: dout  = 8'b11111100; //  824 : 252 - 0xfc -- Background 0x67
      11'h339: dout  = 8'b01101000; //  825 : 104 - 0x68
      11'h33A: dout  = 8'b11111000; //  826 : 248 - 0xf8
      11'h33B: dout  = 8'b10110000; //  827 : 176 - 0xb0
      11'h33C: dout  = 8'b11100000; //  828 : 224 - 0xe0
      11'h33D: dout  = 8'b10000000; //  829 : 128 - 0x80
      11'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Background 0x68
      11'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Background 0x69
      11'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      11'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      11'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      11'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      11'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      11'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Background 0x6a
      11'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Background 0x6b
      11'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      11'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      11'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      11'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Background 0x6c
      11'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      11'h362: dout  = 8'b00000001; //  866 :   1 - 0x1
      11'h363: dout  = 8'b00011101; //  867 :  29 - 0x1d
      11'h364: dout  = 8'b00111110; //  868 :  62 - 0x3e
      11'h365: dout  = 8'b00111111; //  869 :  63 - 0x3f
      11'h366: dout  = 8'b00111111; //  870 :  63 - 0x3f
      11'h367: dout  = 8'b00111111; //  871 :  63 - 0x3f
      11'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Background 0x6d
      11'h369: dout  = 8'b10000000; //  873 : 128 - 0x80
      11'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout  = 8'b01110000; //  875 : 112 - 0x70
      11'h36C: dout  = 8'b11111000; //  876 : 248 - 0xf8
      11'h36D: dout  = 8'b11111100; //  877 : 252 - 0xfc
      11'h36E: dout  = 8'b11111100; //  878 : 252 - 0xfc
      11'h36F: dout  = 8'b11111100; //  879 : 252 - 0xfc
      11'h370: dout  = 8'b00111111; //  880 :  63 - 0x3f -- Background 0x6e
      11'h371: dout  = 8'b00111111; //  881 :  63 - 0x3f
      11'h372: dout  = 8'b00011111; //  882 :  31 - 0x1f
      11'h373: dout  = 8'b00011111; //  883 :  31 - 0x1f
      11'h374: dout  = 8'b00001111; //  884 :  15 - 0xf
      11'h375: dout  = 8'b00000110; //  885 :   6 - 0x6
      11'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout  = 8'b11101100; //  888 : 236 - 0xec -- Background 0x6f
      11'h379: dout  = 8'b11101100; //  889 : 236 - 0xec
      11'h37A: dout  = 8'b11011000; //  890 : 216 - 0xd8
      11'h37B: dout  = 8'b11111000; //  891 : 248 - 0xf8
      11'h37C: dout  = 8'b11110000; //  892 : 240 - 0xf0
      11'h37D: dout  = 8'b11100000; //  893 : 224 - 0xe0
      11'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Background 0x70
      11'h381: dout  = 8'b00000100; //  897 :   4 - 0x4
      11'h382: dout  = 8'b00000011; //  898 :   3 - 0x3
      11'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      11'h384: dout  = 8'b00000001; //  900 :   1 - 0x1
      11'h385: dout  = 8'b00000111; //  901 :   7 - 0x7
      11'h386: dout  = 8'b00001111; //  902 :  15 - 0xf
      11'h387: dout  = 8'b00001100; //  903 :  12 - 0xc
      11'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- Background 0x71
      11'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      11'h38A: dout  = 8'b11100000; //  906 : 224 - 0xe0
      11'h38B: dout  = 8'b10000000; //  907 : 128 - 0x80
      11'h38C: dout  = 8'b01000000; //  908 :  64 - 0x40
      11'h38D: dout  = 8'b11110000; //  909 : 240 - 0xf0
      11'h38E: dout  = 8'b10011000; //  910 : 152 - 0x98
      11'h38F: dout  = 8'b11111000; //  911 : 248 - 0xf8
      11'h390: dout  = 8'b00011111; //  912 :  31 - 0x1f -- Background 0x72
      11'h391: dout  = 8'b00010011; //  913 :  19 - 0x13
      11'h392: dout  = 8'b00011111; //  914 :  31 - 0x1f
      11'h393: dout  = 8'b00001111; //  915 :  15 - 0xf
      11'h394: dout  = 8'b00001001; //  916 :   9 - 0x9
      11'h395: dout  = 8'b00000111; //  917 :   7 - 0x7
      11'h396: dout  = 8'b00000001; //  918 :   1 - 0x1
      11'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      11'h398: dout  = 8'b11100100; //  920 : 228 - 0xe4 -- Background 0x73
      11'h399: dout  = 8'b00111100; //  921 :  60 - 0x3c
      11'h39A: dout  = 8'b11100100; //  922 : 228 - 0xe4
      11'h39B: dout  = 8'b00111000; //  923 :  56 - 0x38
      11'h39C: dout  = 8'b11111000; //  924 : 248 - 0xf8
      11'h39D: dout  = 8'b11110000; //  925 : 240 - 0xf0
      11'h39E: dout  = 8'b11000000; //  926 : 192 - 0xc0
      11'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Background 0x74
      11'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      11'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      11'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      11'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      11'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      11'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      11'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Background 0x75
      11'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      11'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      11'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      11'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      11'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      11'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      11'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      11'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Background 0x76
      11'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      11'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      11'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      11'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      11'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      11'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      11'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      11'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Background 0x77
      11'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      11'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      11'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      11'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      11'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      11'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      11'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- Background 0x79
      11'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Background 0x7a
      11'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      11'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Background 0x7b
      11'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Background 0x7c
      11'h3E1: dout  = 8'b00000001; //  993 :   1 - 0x1
      11'h3E2: dout  = 8'b00000110; //  994 :   6 - 0x6
      11'h3E3: dout  = 8'b00000111; //  995 :   7 - 0x7
      11'h3E4: dout  = 8'b00000111; //  996 :   7 - 0x7
      11'h3E5: dout  = 8'b00000111; //  997 :   7 - 0x7
      11'h3E6: dout  = 8'b00000001; //  998 :   1 - 0x1
      11'h3E7: dout  = 8'b00000011; //  999 :   3 - 0x3
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Background 0x7d
      11'h3E9: dout  = 8'b11000000; // 1001 : 192 - 0xc0
      11'h3EA: dout  = 8'b00110000; // 1002 :  48 - 0x30
      11'h3EB: dout  = 8'b11110000; // 1003 : 240 - 0xf0
      11'h3EC: dout  = 8'b11110000; // 1004 : 240 - 0xf0
      11'h3ED: dout  = 8'b11110000; // 1005 : 240 - 0xf0
      11'h3EE: dout  = 8'b01000000; // 1006 :  64 - 0x40
      11'h3EF: dout  = 8'b01000000; // 1007 :  64 - 0x40
      11'h3F0: dout  = 8'b00000001; // 1008 :   1 - 0x1 -- Background 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b00000001; // 1010 :   1 - 0x1
      11'h3F3: dout  = 8'b00000011; // 1011 :   3 - 0x3
      11'h3F4: dout  = 8'b00000001; // 1012 :   1 - 0x1
      11'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout  = 8'b01000000; // 1016 :  64 - 0x40 -- Background 0x7f
      11'h3F9: dout  = 8'b01000000; // 1017 :  64 - 0x40
      11'h3FA: dout  = 8'b01000000; // 1018 :  64 - 0x40
      11'h3FB: dout  = 8'b01000000; // 1019 :  64 - 0x40
      11'h3FC: dout  = 8'b01000000; // 1020 :  64 - 0x40
      11'h3FD: dout  = 8'b10000000; // 1021 : 128 - 0x80
      11'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      11'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      11'h400: dout  = 8'b11111111; // 1024 : 255 - 0xff -- Background 0x80
      11'h401: dout  = 8'b11111111; // 1025 : 255 - 0xff
      11'h402: dout  = 8'b11111111; // 1026 : 255 - 0xff
      11'h403: dout  = 8'b11111111; // 1027 : 255 - 0xff
      11'h404: dout  = 8'b11000000; // 1028 : 192 - 0xc0
      11'h405: dout  = 8'b11000000; // 1029 : 192 - 0xc0
      11'h406: dout  = 8'b11000000; // 1030 : 192 - 0xc0
      11'h407: dout  = 8'b11000111; // 1031 : 199 - 0xc7
      11'h408: dout  = 8'b11111111; // 1032 : 255 - 0xff -- Background 0x81
      11'h409: dout  = 8'b11111111; // 1033 : 255 - 0xff
      11'h40A: dout  = 8'b11111111; // 1034 : 255 - 0xff
      11'h40B: dout  = 8'b11111111; // 1035 : 255 - 0xff
      11'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      11'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      11'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      11'h40F: dout  = 8'b11111111; // 1039 : 255 - 0xff
      11'h410: dout  = 8'b11111111; // 1040 : 255 - 0xff -- Background 0x82
      11'h411: dout  = 8'b11111111; // 1041 : 255 - 0xff
      11'h412: dout  = 8'b11111111; // 1042 : 255 - 0xff
      11'h413: dout  = 8'b11111111; // 1043 : 255 - 0xff
      11'h414: dout  = 8'b01111111; // 1044 : 127 - 0x7f
      11'h415: dout  = 8'b00111111; // 1045 :  63 - 0x3f
      11'h416: dout  = 8'b00011111; // 1046 :  31 - 0x1f
      11'h417: dout  = 8'b11001111; // 1047 : 207 - 0xcf
      11'h418: dout  = 8'b11111111; // 1048 : 255 - 0xff -- Background 0x83
      11'h419: dout  = 8'b11111111; // 1049 : 255 - 0xff
      11'h41A: dout  = 8'b11111111; // 1050 : 255 - 0xff
      11'h41B: dout  = 8'b11110111; // 1051 : 247 - 0xf7
      11'h41C: dout  = 8'b11110111; // 1052 : 247 - 0xf7
      11'h41D: dout  = 8'b11100010; // 1053 : 226 - 0xe2
      11'h41E: dout  = 8'b11100000; // 1054 : 224 - 0xe0
      11'h41F: dout  = 8'b11000110; // 1055 : 198 - 0xc6
      11'h420: dout  = 8'b11111111; // 1056 : 255 - 0xff -- Background 0x84
      11'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout  = 8'b11111111; // 1058 : 255 - 0xff
      11'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout  = 8'b10111111; // 1060 : 191 - 0xbf
      11'h425: dout  = 8'b10111111; // 1061 : 191 - 0xbf
      11'h426: dout  = 8'b00011111; // 1062 :  31 - 0x1f
      11'h427: dout  = 8'b00011111; // 1063 :  31 - 0x1f
      11'h428: dout  = 8'b11111111; // 1064 : 255 - 0xff -- Background 0x85
      11'h429: dout  = 8'b11111111; // 1065 : 255 - 0xff
      11'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      11'h42B: dout  = 8'b11111111; // 1067 : 255 - 0xff
      11'h42C: dout  = 8'b11111110; // 1068 : 254 - 0xfe
      11'h42D: dout  = 8'b11111000; // 1069 : 248 - 0xf8
      11'h42E: dout  = 8'b11100000; // 1070 : 224 - 0xe0
      11'h42F: dout  = 8'b11000000; // 1071 : 192 - 0xc0
      11'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Background 0x86
      11'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      11'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      11'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      11'h434: dout  = 8'b00000111; // 1076 :   7 - 0x7
      11'h435: dout  = 8'b00000000; // 1077 :   0 - 0x0
      11'h436: dout  = 8'b00111111; // 1078 :  63 - 0x3f
      11'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      11'h438: dout  = 8'b11111111; // 1080 : 255 - 0xff -- Background 0x87
      11'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout  = 8'b11111111; // 1085 : 255 - 0xff
      11'h43E: dout  = 8'b00111111; // 1086 :  63 - 0x3f
      11'h43F: dout  = 8'b11001111; // 1087 : 207 - 0xcf
      11'h440: dout  = 8'b11111111; // 1088 : 255 - 0xff -- Background 0x88
      11'h441: dout  = 8'b11111111; // 1089 : 255 - 0xff
      11'h442: dout  = 8'b11111111; // 1090 : 255 - 0xff
      11'h443: dout  = 8'b11111111; // 1091 : 255 - 0xff
      11'h444: dout  = 8'b11111111; // 1092 : 255 - 0xff
      11'h445: dout  = 8'b11111111; // 1093 : 255 - 0xff
      11'h446: dout  = 8'b11111111; // 1094 : 255 - 0xff
      11'h447: dout  = 8'b11111111; // 1095 : 255 - 0xff
      11'h448: dout  = 8'b11111111; // 1096 : 255 - 0xff -- Background 0x89
      11'h449: dout  = 8'b11111111; // 1097 : 255 - 0xff
      11'h44A: dout  = 8'b11111111; // 1098 : 255 - 0xff
      11'h44B: dout  = 8'b01110111; // 1099 : 119 - 0x77
      11'h44C: dout  = 8'b00010011; // 1100 :  19 - 0x13
      11'h44D: dout  = 8'b00000001; // 1101 :   1 - 0x1
      11'h44E: dout  = 8'b00010000; // 1102 :  16 - 0x10
      11'h44F: dout  = 8'b00011000; // 1103 :  24 - 0x18
      11'h450: dout  = 8'b11111111; // 1104 : 255 - 0xff -- Background 0x8a
      11'h451: dout  = 8'b11111111; // 1105 : 255 - 0xff
      11'h452: dout  = 8'b11111111; // 1106 : 255 - 0xff
      11'h453: dout  = 8'b11111111; // 1107 : 255 - 0xff
      11'h454: dout  = 8'b11111111; // 1108 : 255 - 0xff
      11'h455: dout  = 8'b11111111; // 1109 : 255 - 0xff
      11'h456: dout  = 8'b11111111; // 1110 : 255 - 0xff
      11'h457: dout  = 8'b01111111; // 1111 : 127 - 0x7f
      11'h458: dout  = 8'b11111111; // 1112 : 255 - 0xff -- Background 0x8b
      11'h459: dout  = 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout  = 8'b11111111; // 1114 : 255 - 0xff
      11'h45B: dout  = 8'b11110111; // 1115 : 247 - 0xf7
      11'h45C: dout  = 8'b11100101; // 1116 : 229 - 0xe5
      11'h45D: dout  = 8'b11000001; // 1117 : 193 - 0xc1
      11'h45E: dout  = 8'b10000100; // 1118 : 132 - 0x84
      11'h45F: dout  = 8'b00001100; // 1119 :  12 - 0xc
      11'h460: dout  = 8'b11111111; // 1120 : 255 - 0xff -- Background 0x8c
      11'h461: dout  = 8'b11111111; // 1121 : 255 - 0xff
      11'h462: dout  = 8'b11111111; // 1122 : 255 - 0xff
      11'h463: dout  = 8'b11111111; // 1123 : 255 - 0xff
      11'h464: dout  = 8'b11111111; // 1124 : 255 - 0xff
      11'h465: dout  = 8'b01111111; // 1125 : 127 - 0x7f
      11'h466: dout  = 8'b01111110; // 1126 : 126 - 0x7e
      11'h467: dout  = 8'b01111110; // 1127 : 126 - 0x7e
      11'h468: dout  = 8'b11111111; // 1128 : 255 - 0xff -- Background 0x8d
      11'h469: dout  = 8'b11111111; // 1129 : 255 - 0xff
      11'h46A: dout  = 8'b10111111; // 1130 : 191 - 0xbf
      11'h46B: dout  = 8'b10110111; // 1131 : 183 - 0xb7
      11'h46C: dout  = 8'b00010111; // 1132 :  23 - 0x17
      11'h46D: dout  = 8'b00000011; // 1133 :   3 - 0x3
      11'h46E: dout  = 8'b00100011; // 1134 :  35 - 0x23
      11'h46F: dout  = 8'b00100001; // 1135 :  33 - 0x21
      11'h470: dout  = 8'b11111111; // 1136 : 255 - 0xff -- Background 0x8e
      11'h471: dout  = 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout  = 8'b11111011; // 1138 : 251 - 0xfb
      11'h473: dout  = 8'b11111001; // 1139 : 249 - 0xf9
      11'h474: dout  = 8'b11111000; // 1140 : 248 - 0xf8
      11'h475: dout  = 8'b11111000; // 1141 : 248 - 0xf8
      11'h476: dout  = 8'b11111000; // 1142 : 248 - 0xf8
      11'h477: dout  = 8'b11111000; // 1143 : 248 - 0xf8
      11'h478: dout  = 8'b11111111; // 1144 : 255 - 0xff -- Background 0x8f
      11'h479: dout  = 8'b11111111; // 1145 : 255 - 0xff
      11'h47A: dout  = 8'b01111000; // 1146 : 120 - 0x78
      11'h47B: dout  = 8'b00111000; // 1147 :  56 - 0x38
      11'h47C: dout  = 8'b00011000; // 1148 :  24 - 0x18
      11'h47D: dout  = 8'b00001000; // 1149 :   8 - 0x8
      11'h47E: dout  = 8'b10000000; // 1150 : 128 - 0x80
      11'h47F: dout  = 8'b11000000; // 1151 : 192 - 0xc0
      11'h480: dout  = 8'b11111111; // 1152 : 255 - 0xff -- Background 0x90
      11'h481: dout  = 8'b11111111; // 1153 : 255 - 0xff
      11'h482: dout  = 8'b00000001; // 1154 :   1 - 0x1
      11'h483: dout  = 8'b00000001; // 1155 :   1 - 0x1
      11'h484: dout  = 8'b00000001; // 1156 :   1 - 0x1
      11'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      11'h486: dout  = 8'b11111111; // 1158 : 255 - 0xff
      11'h487: dout  = 8'b11111111; // 1159 : 255 - 0xff
      11'h488: dout  = 8'b11111111; // 1160 : 255 - 0xff -- Background 0x91
      11'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout  = 8'b11111111; // 1162 : 255 - 0xff
      11'h48B: dout  = 8'b11111111; // 1163 : 255 - 0xff
      11'h48C: dout  = 8'b11111111; // 1164 : 255 - 0xff
      11'h48D: dout  = 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout  = 8'b01111111; // 1166 : 127 - 0x7f
      11'h48F: dout  = 8'b00111111; // 1167 :  63 - 0x3f
      11'h490: dout  = 8'b11000111; // 1168 : 199 - 0xc7 -- Background 0x92
      11'h491: dout  = 8'b11000111; // 1169 : 199 - 0xc7
      11'h492: dout  = 8'b11000111; // 1170 : 199 - 0xc7
      11'h493: dout  = 8'b11000111; // 1171 : 199 - 0xc7
      11'h494: dout  = 8'b11000111; // 1172 : 199 - 0xc7
      11'h495: dout  = 8'b11000111; // 1173 : 199 - 0xc7
      11'h496: dout  = 8'b11000111; // 1174 : 199 - 0xc7
      11'h497: dout  = 8'b11000111; // 1175 : 199 - 0xc7
      11'h498: dout  = 8'b11111111; // 1176 : 255 - 0xff -- Background 0x93
      11'h499: dout  = 8'b11111111; // 1177 : 255 - 0xff
      11'h49A: dout  = 8'b11111111; // 1178 : 255 - 0xff
      11'h49B: dout  = 8'b11111111; // 1179 : 255 - 0xff
      11'h49C: dout  = 8'b11111001; // 1180 : 249 - 0xf9
      11'h49D: dout  = 8'b11111001; // 1181 : 249 - 0xf9
      11'h49E: dout  = 8'b11111111; // 1182 : 255 - 0xff
      11'h49F: dout  = 8'b11111111; // 1183 : 255 - 0xff
      11'h4A0: dout  = 8'b11110111; // 1184 : 247 - 0xf7 -- Background 0x94
      11'h4A1: dout  = 8'b11111011; // 1185 : 251 - 0xfb
      11'h4A2: dout  = 8'b11111011; // 1186 : 251 - 0xfb
      11'h4A3: dout  = 8'b11111101; // 1187 : 253 - 0xfd
      11'h4A4: dout  = 8'b11111100; // 1188 : 252 - 0xfc
      11'h4A5: dout  = 8'b11111100; // 1189 : 252 - 0xfc
      11'h4A6: dout  = 8'b01111100; // 1190 : 124 - 0x7c
      11'h4A7: dout  = 8'b01111100; // 1191 : 124 - 0x7c
      11'h4A8: dout  = 8'b11000111; // 1192 : 199 - 0xc7 -- Background 0x95
      11'h4A9: dout  = 8'b10001111; // 1193 : 143 - 0x8f
      11'h4AA: dout  = 8'b10001111; // 1194 : 143 - 0x8f
      11'h4AB: dout  = 8'b00011111; // 1195 :  31 - 0x1f
      11'h4AC: dout  = 8'b00011111; // 1196 :  31 - 0x1f
      11'h4AD: dout  = 8'b00111111; // 1197 :  63 - 0x3f
      11'h4AE: dout  = 8'b00111111; // 1198 :  63 - 0x3f
      11'h4AF: dout  = 8'b01111111; // 1199 : 127 - 0x7f
      11'h4B0: dout  = 8'b00001111; // 1200 :  15 - 0xf -- Background 0x96
      11'h4B1: dout  = 8'b00001111; // 1201 :  15 - 0xf
      11'h4B2: dout  = 8'b10000111; // 1202 : 135 - 0x87
      11'h4B3: dout  = 8'b10000111; // 1203 : 135 - 0x87
      11'h4B4: dout  = 8'b11000010; // 1204 : 194 - 0xc2
      11'h4B5: dout  = 8'b11000010; // 1205 : 194 - 0xc2
      11'h4B6: dout  = 8'b11100000; // 1206 : 224 - 0xe0
      11'h4B7: dout  = 8'b11100000; // 1207 : 224 - 0xe0
      11'h4B8: dout  = 8'b10000011; // 1208 : 131 - 0x83 -- Background 0x97
      11'h4B9: dout  = 8'b10001111; // 1209 : 143 - 0x8f
      11'h4BA: dout  = 8'b00001111; // 1210 :  15 - 0xf
      11'h4BB: dout  = 8'b00011111; // 1211 :  31 - 0x1f
      11'h4BC: dout  = 8'b00011111; // 1212 :  31 - 0x1f
      11'h4BD: dout  = 8'b00111111; // 1213 :  63 - 0x3f
      11'h4BE: dout  = 8'b00111111; // 1214 :  63 - 0x3f
      11'h4BF: dout  = 8'b00111111; // 1215 :  63 - 0x3f
      11'h4C0: dout  = 8'b11111111; // 1216 : 255 - 0xff -- Background 0x98
      11'h4C1: dout  = 8'b11111111; // 1217 : 255 - 0xff
      11'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      11'h4C3: dout  = 8'b11111110; // 1219 : 254 - 0xfe
      11'h4C4: dout  = 8'b11111001; // 1220 : 249 - 0xf9
      11'h4C5: dout  = 8'b11100111; // 1221 : 231 - 0xe7
      11'h4C6: dout  = 8'b11111100; // 1222 : 252 - 0xfc
      11'h4C7: dout  = 8'b11110000; // 1223 : 240 - 0xf0
      11'h4C8: dout  = 8'b11110111; // 1224 : 247 - 0xf7 -- Background 0x99
      11'h4C9: dout  = 8'b11111011; // 1225 : 251 - 0xfb
      11'h4CA: dout  = 8'b11111011; // 1226 : 251 - 0xfb
      11'h4CB: dout  = 8'b01110011; // 1227 : 115 - 0x73
      11'h4CC: dout  = 8'b11000001; // 1228 : 193 - 0xc1
      11'h4CD: dout  = 8'b00000011; // 1229 :   3 - 0x3
      11'h4CE: dout  = 8'b00001111; // 1230 :  15 - 0xf
      11'h4CF: dout  = 8'b00111111; // 1231 :  63 - 0x3f
      11'h4D0: dout  = 8'b11111111; // 1232 : 255 - 0xff -- Background 0x9a
      11'h4D1: dout  = 8'b11111111; // 1233 : 255 - 0xff
      11'h4D2: dout  = 8'b11111111; // 1234 : 255 - 0xff
      11'h4D3: dout  = 8'b10000000; // 1235 : 128 - 0x80
      11'h4D4: dout  = 8'b10000000; // 1236 : 128 - 0x80
      11'h4D5: dout  = 8'b10000000; // 1237 : 128 - 0x80
      11'h4D6: dout  = 8'b10001111; // 1238 : 143 - 0x8f
      11'h4D7: dout  = 8'b10001111; // 1239 : 143 - 0x8f
      11'h4D8: dout  = 8'b11111111; // 1240 : 255 - 0xff -- Background 0x9b
      11'h4D9: dout  = 8'b11111111; // 1241 : 255 - 0xff
      11'h4DA: dout  = 8'b11111111; // 1242 : 255 - 0xff
      11'h4DB: dout  = 8'b00001111; // 1243 :  15 - 0xf
      11'h4DC: dout  = 8'b00001111; // 1244 :  15 - 0xf
      11'h4DD: dout  = 8'b00000111; // 1245 :   7 - 0x7
      11'h4DE: dout  = 8'b11110111; // 1246 : 247 - 0xf7
      11'h4DF: dout  = 8'b11110001; // 1247 : 241 - 0xf1
      11'h4E0: dout  = 8'b00011100; // 1248 :  28 - 0x1c -- Background 0x9c
      11'h4E1: dout  = 8'b00011110; // 1249 :  30 - 0x1e
      11'h4E2: dout  = 8'b00011111; // 1250 :  31 - 0x1f
      11'h4E3: dout  = 8'b00011111; // 1251 :  31 - 0x1f
      11'h4E4: dout  = 8'b00011111; // 1252 :  31 - 0x1f
      11'h4E5: dout  = 8'b00011111; // 1253 :  31 - 0x1f
      11'h4E6: dout  = 8'b00011111; // 1254 :  31 - 0x1f
      11'h4E7: dout  = 8'b00011111; // 1255 :  31 - 0x1f
      11'h4E8: dout  = 8'b00111110; // 1256 :  62 - 0x3e -- Background 0x9d
      11'h4E9: dout  = 8'b00011100; // 1257 :  28 - 0x1c
      11'h4EA: dout  = 8'b00001000; // 1258 :   8 - 0x8
      11'h4EB: dout  = 8'b10000000; // 1259 : 128 - 0x80
      11'h4EC: dout  = 8'b11000001; // 1260 : 193 - 0xc1
      11'h4ED: dout  = 8'b11100011; // 1261 : 227 - 0xe3
      11'h4EE: dout  = 8'b11110111; // 1262 : 247 - 0xf7
      11'h4EF: dout  = 8'b11111111; // 1263 : 255 - 0xff
      11'h4F0: dout  = 8'b00011100; // 1264 :  28 - 0x1c -- Background 0x9e
      11'h4F1: dout  = 8'b00111100; // 1265 :  60 - 0x3c
      11'h4F2: dout  = 8'b01111100; // 1266 : 124 - 0x7c
      11'h4F3: dout  = 8'b11111100; // 1267 : 252 - 0xfc
      11'h4F4: dout  = 8'b11111100; // 1268 : 252 - 0xfc
      11'h4F5: dout  = 8'b11111100; // 1269 : 252 - 0xfc
      11'h4F6: dout  = 8'b11111100; // 1270 : 252 - 0xfc
      11'h4F7: dout  = 8'b11111100; // 1271 : 252 - 0xfc
      11'h4F8: dout  = 8'b01111100; // 1272 : 124 - 0x7c -- Background 0x9f
      11'h4F9: dout  = 8'b01111100; // 1273 : 124 - 0x7c
      11'h4FA: dout  = 8'b01111000; // 1274 : 120 - 0x78
      11'h4FB: dout  = 8'b01111000; // 1275 : 120 - 0x78
      11'h4FC: dout  = 8'b01110001; // 1276 : 113 - 0x71
      11'h4FD: dout  = 8'b01110001; // 1277 : 113 - 0x71
      11'h4FE: dout  = 8'b01100011; // 1278 :  99 - 0x63
      11'h4FF: dout  = 8'b01100011; // 1279 :  99 - 0x63
      11'h500: dout  = 8'b01110001; // 1280 : 113 - 0x71 -- Background 0xa0
      11'h501: dout  = 8'b01110000; // 1281 : 112 - 0x70
      11'h502: dout  = 8'b11111000; // 1282 : 248 - 0xf8
      11'h503: dout  = 8'b11111000; // 1283 : 248 - 0xf8
      11'h504: dout  = 8'b11111100; // 1284 : 252 - 0xfc
      11'h505: dout  = 8'b11111100; // 1285 : 252 - 0xfc
      11'h506: dout  = 8'b11111110; // 1286 : 254 - 0xfe
      11'h507: dout  = 8'b11111110; // 1287 : 254 - 0xfe
      11'h508: dout  = 8'b11111000; // 1288 : 248 - 0xf8 -- Background 0xa1
      11'h509: dout  = 8'b11111000; // 1289 : 248 - 0xf8
      11'h50A: dout  = 8'b11111000; // 1290 : 248 - 0xf8
      11'h50B: dout  = 8'b01111000; // 1291 : 120 - 0x78
      11'h50C: dout  = 8'b01111000; // 1292 : 120 - 0x78
      11'h50D: dout  = 8'b00111000; // 1293 :  56 - 0x38
      11'h50E: dout  = 8'b00111000; // 1294 :  56 - 0x38
      11'h50F: dout  = 8'b00011000; // 1295 :  24 - 0x18
      11'h510: dout  = 8'b11100000; // 1296 : 224 - 0xe0 -- Background 0xa2
      11'h511: dout  = 8'b11110000; // 1297 : 240 - 0xf0
      11'h512: dout  = 8'b11111000; // 1298 : 248 - 0xf8
      11'h513: dout  = 8'b11111000; // 1299 : 248 - 0xf8
      11'h514: dout  = 8'b11111100; // 1300 : 252 - 0xfc
      11'h515: dout  = 8'b11111100; // 1301 : 252 - 0xfc
      11'h516: dout  = 8'b11111110; // 1302 : 254 - 0xfe
      11'h517: dout  = 8'b11111111; // 1303 : 255 - 0xff
      11'h518: dout  = 8'b11111111; // 1304 : 255 - 0xff -- Background 0xa3
      11'h519: dout  = 8'b11111111; // 1305 : 255 - 0xff
      11'h51A: dout  = 8'b11111111; // 1306 : 255 - 0xff
      11'h51B: dout  = 8'b11111111; // 1307 : 255 - 0xff
      11'h51C: dout  = 8'b11111111; // 1308 : 255 - 0xff
      11'h51D: dout  = 8'b11111111; // 1309 : 255 - 0xff
      11'h51E: dout  = 8'b11111111; // 1310 : 255 - 0xff
      11'h51F: dout  = 8'b11111111; // 1311 : 255 - 0xff
      11'h520: dout  = 8'b00011111; // 1312 :  31 - 0x1f -- Background 0xa4
      11'h521: dout  = 8'b00011111; // 1313 :  31 - 0x1f
      11'h522: dout  = 8'b00011111; // 1314 :  31 - 0x1f
      11'h523: dout  = 8'b00011111; // 1315 :  31 - 0x1f
      11'h524: dout  = 8'b00011111; // 1316 :  31 - 0x1f
      11'h525: dout  = 8'b00011111; // 1317 :  31 - 0x1f
      11'h526: dout  = 8'b00011111; // 1318 :  31 - 0x1f
      11'h527: dout  = 8'b00011111; // 1319 :  31 - 0x1f
      11'h528: dout  = 8'b11111000; // 1320 : 248 - 0xf8 -- Background 0xa5
      11'h529: dout  = 8'b11111111; // 1321 : 255 - 0xff
      11'h52A: dout  = 8'b11111111; // 1322 : 255 - 0xff
      11'h52B: dout  = 8'b11111000; // 1323 : 248 - 0xf8
      11'h52C: dout  = 8'b11111000; // 1324 : 248 - 0xf8
      11'h52D: dout  = 8'b11111000; // 1325 : 248 - 0xf8
      11'h52E: dout  = 8'b11111000; // 1326 : 248 - 0xf8
      11'h52F: dout  = 8'b11111000; // 1327 : 248 - 0xf8
      11'h530: dout  = 8'b11111100; // 1328 : 252 - 0xfc -- Background 0xa6
      11'h531: dout  = 8'b11111000; // 1329 : 248 - 0xf8
      11'h532: dout  = 8'b11110000; // 1330 : 240 - 0xf0
      11'h533: dout  = 8'b00000001; // 1331 :   1 - 0x1
      11'h534: dout  = 8'b00000001; // 1332 :   1 - 0x1
      11'h535: dout  = 8'b00000011; // 1333 :   3 - 0x3
      11'h536: dout  = 8'b11000011; // 1334 : 195 - 0xc3
      11'h537: dout  = 8'b10000111; // 1335 : 135 - 0x87
      11'h538: dout  = 8'b01111111; // 1336 : 127 - 0x7f -- Background 0xa7
      11'h539: dout  = 8'b11111001; // 1337 : 249 - 0xf9
      11'h53A: dout  = 8'b11111001; // 1338 : 249 - 0xf9
      11'h53B: dout  = 8'b11111111; // 1339 : 255 - 0xff
      11'h53C: dout  = 8'b11111110; // 1340 : 254 - 0xfe
      11'h53D: dout  = 8'b11111100; // 1341 : 252 - 0xfc
      11'h53E: dout  = 8'b11111111; // 1342 : 255 - 0xff
      11'h53F: dout  = 8'b11111111; // 1343 : 255 - 0xff
      11'h540: dout  = 8'b11110000; // 1344 : 240 - 0xf0 -- Background 0xa8
      11'h541: dout  = 8'b11110000; // 1345 : 240 - 0xf0
      11'h542: dout  = 8'b11111000; // 1346 : 248 - 0xf8
      11'h543: dout  = 8'b01111000; // 1347 : 120 - 0x78
      11'h544: dout  = 8'b11111100; // 1348 : 252 - 0xfc
      11'h545: dout  = 8'b11110100; // 1349 : 244 - 0xf4
      11'h546: dout  = 8'b11110110; // 1350 : 246 - 0xf6
      11'h547: dout  = 8'b11111010; // 1351 : 250 - 0xfa
      11'h548: dout  = 8'b00111111; // 1352 :  63 - 0x3f -- Background 0xa9
      11'h549: dout  = 8'b00111111; // 1353 :  63 - 0x3f
      11'h54A: dout  = 8'b00111111; // 1354 :  63 - 0x3f
      11'h54B: dout  = 8'b00111111; // 1355 :  63 - 0x3f
      11'h54C: dout  = 8'b00111111; // 1356 :  63 - 0x3f
      11'h54D: dout  = 8'b00011111; // 1357 :  31 - 0x1f
      11'h54E: dout  = 8'b00001111; // 1358 :  15 - 0xf
      11'h54F: dout  = 8'b00000111; // 1359 :   7 - 0x7
      11'h550: dout  = 8'b11100000; // 1360 : 224 - 0xe0 -- Background 0xaa
      11'h551: dout  = 8'b11111000; // 1361 : 248 - 0xf8
      11'h552: dout  = 8'b11111111; // 1362 : 255 - 0xff
      11'h553: dout  = 8'b11110011; // 1363 : 243 - 0xf3
      11'h554: dout  = 8'b11111100; // 1364 : 252 - 0xfc
      11'h555: dout  = 8'b11111111; // 1365 : 255 - 0xff
      11'h556: dout  = 8'b11111111; // 1366 : 255 - 0xff
      11'h557: dout  = 8'b11111111; // 1367 : 255 - 0xff
      11'h558: dout  = 8'b11111111; // 1368 : 255 - 0xff -- Background 0xab
      11'h559: dout  = 8'b11111111; // 1369 : 255 - 0xff
      11'h55A: dout  = 8'b00111111; // 1370 :  63 - 0x3f
      11'h55B: dout  = 8'b11001111; // 1371 : 207 - 0xcf
      11'h55C: dout  = 8'b11110011; // 1372 : 243 - 0xf3
      11'h55D: dout  = 8'b00111101; // 1373 :  61 - 0x3d
      11'h55E: dout  = 8'b11011000; // 1374 : 216 - 0xd8
      11'h55F: dout  = 8'b10110000; // 1375 : 176 - 0xb0
      11'h560: dout  = 8'b10001111; // 1376 : 143 - 0x8f -- Background 0xac
      11'h561: dout  = 8'b11101111; // 1377 : 239 - 0xef
      11'h562: dout  = 8'b11100000; // 1378 : 224 - 0xe0
      11'h563: dout  = 8'b11111000; // 1379 : 248 - 0xf8
      11'h564: dout  = 8'b11111000; // 1380 : 248 - 0xf8
      11'h565: dout  = 8'b11111111; // 1381 : 255 - 0xff
      11'h566: dout  = 8'b11111111; // 1382 : 255 - 0xff
      11'h567: dout  = 8'b11111111; // 1383 : 255 - 0xff
      11'h568: dout  = 8'b11110001; // 1384 : 241 - 0xf1 -- Background 0xad
      11'h569: dout  = 8'b11110001; // 1385 : 241 - 0xf1
      11'h56A: dout  = 8'b00000001; // 1386 :   1 - 0x1
      11'h56B: dout  = 8'b00000001; // 1387 :   1 - 0x1
      11'h56C: dout  = 8'b00000001; // 1388 :   1 - 0x1
      11'h56D: dout  = 8'b11111111; // 1389 : 255 - 0xff
      11'h56E: dout  = 8'b11111111; // 1390 : 255 - 0xff
      11'h56F: dout  = 8'b11111111; // 1391 : 255 - 0xff
      11'h570: dout  = 8'b00011111; // 1392 :  31 - 0x1f -- Background 0xae
      11'h571: dout  = 8'b00011111; // 1393 :  31 - 0x1f
      11'h572: dout  = 8'b00011111; // 1394 :  31 - 0x1f
      11'h573: dout  = 8'b00011111; // 1395 :  31 - 0x1f
      11'h574: dout  = 8'b00011111; // 1396 :  31 - 0x1f
      11'h575: dout  = 8'b00011111; // 1397 :  31 - 0x1f
      11'h576: dout  = 8'b00011111; // 1398 :  31 - 0x1f
      11'h577: dout  = 8'b00011111; // 1399 :  31 - 0x1f
      11'h578: dout  = 8'b11111100; // 1400 : 252 - 0xfc -- Background 0xaf
      11'h579: dout  = 8'b11111100; // 1401 : 252 - 0xfc
      11'h57A: dout  = 8'b11111100; // 1402 : 252 - 0xfc
      11'h57B: dout  = 8'b11111100; // 1403 : 252 - 0xfc
      11'h57C: dout  = 8'b11110100; // 1404 : 244 - 0xf4
      11'h57D: dout  = 8'b11110100; // 1405 : 244 - 0xf4
      11'h57E: dout  = 8'b11110100; // 1406 : 244 - 0xf4
      11'h57F: dout  = 8'b11110100; // 1407 : 244 - 0xf4
      11'h580: dout  = 8'b00001100; // 1408 :  12 - 0xc -- Background 0xb0
      11'h581: dout  = 8'b00011100; // 1409 :  28 - 0x1c
      11'h582: dout  = 8'b00001100; // 1410 :  12 - 0xc
      11'h583: dout  = 8'b00001100; // 1411 :  12 - 0xc
      11'h584: dout  = 8'b00001100; // 1412 :  12 - 0xc
      11'h585: dout  = 8'b00001100; // 1413 :  12 - 0xc
      11'h586: dout  = 8'b00111111; // 1414 :  63 - 0x3f
      11'h587: dout  = 8'b00000000; // 1415 :   0 - 0x0
      11'h588: dout  = 8'b00111110; // 1416 :  62 - 0x3e -- Background 0xb1
      11'h589: dout  = 8'b01100011; // 1417 :  99 - 0x63
      11'h58A: dout  = 8'b00000111; // 1418 :   7 - 0x7
      11'h58B: dout  = 8'b00011110; // 1419 :  30 - 0x1e
      11'h58C: dout  = 8'b00111100; // 1420 :  60 - 0x3c
      11'h58D: dout  = 8'b01110000; // 1421 : 112 - 0x70
      11'h58E: dout  = 8'b01111111; // 1422 : 127 - 0x7f
      11'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      11'h590: dout  = 8'b01111110; // 1424 : 126 - 0x7e -- Background 0xb2
      11'h591: dout  = 8'b01100011; // 1425 :  99 - 0x63
      11'h592: dout  = 8'b01100011; // 1426 :  99 - 0x63
      11'h593: dout  = 8'b01100011; // 1427 :  99 - 0x63
      11'h594: dout  = 8'b01111110; // 1428 : 126 - 0x7e
      11'h595: dout  = 8'b01100000; // 1429 :  96 - 0x60
      11'h596: dout  = 8'b01100000; // 1430 :  96 - 0x60
      11'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout  = 8'b01100011; // 1432 :  99 - 0x63 -- Background 0xb3
      11'h599: dout  = 8'b01100011; // 1433 :  99 - 0x63
      11'h59A: dout  = 8'b01100011; // 1434 :  99 - 0x63
      11'h59B: dout  = 8'b01100011; // 1435 :  99 - 0x63
      11'h59C: dout  = 8'b01100011; // 1436 :  99 - 0x63
      11'h59D: dout  = 8'b01100011; // 1437 :  99 - 0x63
      11'h59E: dout  = 8'b00111110; // 1438 :  62 - 0x3e
      11'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout  = 8'b01100011; // 1440 :  99 - 0x63 -- Background 0xb4
      11'h5A1: dout  = 8'b01100011; // 1441 :  99 - 0x63
      11'h5A2: dout  = 8'b01100011; // 1442 :  99 - 0x63
      11'h5A3: dout  = 8'b01111111; // 1443 : 127 - 0x7f
      11'h5A4: dout  = 8'b01100011; // 1444 :  99 - 0x63
      11'h5A5: dout  = 8'b01100011; // 1445 :  99 - 0x63
      11'h5A6: dout  = 8'b01100011; // 1446 :  99 - 0x63
      11'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout  = 8'b00111111; // 1448 :  63 - 0x3f -- Background 0xb5
      11'h5A9: dout  = 8'b00001100; // 1449 :  12 - 0xc
      11'h5AA: dout  = 8'b00001100; // 1450 :  12 - 0xc
      11'h5AB: dout  = 8'b00001100; // 1451 :  12 - 0xc
      11'h5AC: dout  = 8'b00001100; // 1452 :  12 - 0xc
      11'h5AD: dout  = 8'b00001100; // 1453 :  12 - 0xc
      11'h5AE: dout  = 8'b00111111; // 1454 :  63 - 0x3f
      11'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Background 0xb6
      11'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      11'h5B2: dout  = 8'b00000000; // 1458 :   0 - 0x0
      11'h5B3: dout  = 8'b01111110; // 1459 : 126 - 0x7e
      11'h5B4: dout  = 8'b00000000; // 1460 :   0 - 0x0
      11'h5B5: dout  = 8'b00000000; // 1461 :   0 - 0x0
      11'h5B6: dout  = 8'b00000000; // 1462 :   0 - 0x0
      11'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout  = 8'b00111100; // 1464 :  60 - 0x3c -- Background 0xb7
      11'h5B9: dout  = 8'b01100110; // 1465 : 102 - 0x66
      11'h5BA: dout  = 8'b01100000; // 1466 :  96 - 0x60
      11'h5BB: dout  = 8'b00111110; // 1467 :  62 - 0x3e
      11'h5BC: dout  = 8'b00000011; // 1468 :   3 - 0x3
      11'h5BD: dout  = 8'b01100011; // 1469 :  99 - 0x63
      11'h5BE: dout  = 8'b00111110; // 1470 :  62 - 0x3e
      11'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout  = 8'b00011110; // 1472 :  30 - 0x1e -- Background 0xb8
      11'h5C1: dout  = 8'b00110011; // 1473 :  51 - 0x33
      11'h5C2: dout  = 8'b01100000; // 1474 :  96 - 0x60
      11'h5C3: dout  = 8'b01100000; // 1475 :  96 - 0x60
      11'h5C4: dout  = 8'b01100000; // 1476 :  96 - 0x60
      11'h5C5: dout  = 8'b00110011; // 1477 :  51 - 0x33
      11'h5C6: dout  = 8'b00011110; // 1478 :  30 - 0x1e
      11'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout  = 8'b00111110; // 1480 :  62 - 0x3e -- Background 0xb9
      11'h5C9: dout  = 8'b01100011; // 1481 :  99 - 0x63
      11'h5CA: dout  = 8'b01100011; // 1482 :  99 - 0x63
      11'h5CB: dout  = 8'b01100011; // 1483 :  99 - 0x63
      11'h5CC: dout  = 8'b01100011; // 1484 :  99 - 0x63
      11'h5CD: dout  = 8'b01100011; // 1485 :  99 - 0x63
      11'h5CE: dout  = 8'b00111110; // 1486 :  62 - 0x3e
      11'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout  = 8'b01111110; // 1488 : 126 - 0x7e -- Background 0xba
      11'h5D1: dout  = 8'b01100011; // 1489 :  99 - 0x63
      11'h5D2: dout  = 8'b01100011; // 1490 :  99 - 0x63
      11'h5D3: dout  = 8'b01100111; // 1491 : 103 - 0x67
      11'h5D4: dout  = 8'b01111100; // 1492 : 124 - 0x7c
      11'h5D5: dout  = 8'b01101110; // 1493 : 110 - 0x6e
      11'h5D6: dout  = 8'b01100111; // 1494 : 103 - 0x67
      11'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout  = 8'b01111111; // 1496 : 127 - 0x7f -- Background 0xbb
      11'h5D9: dout  = 8'b01100000; // 1497 :  96 - 0x60
      11'h5DA: dout  = 8'b01100000; // 1498 :  96 - 0x60
      11'h5DB: dout  = 8'b01111110; // 1499 : 126 - 0x7e
      11'h5DC: dout  = 8'b01100000; // 1500 :  96 - 0x60
      11'h5DD: dout  = 8'b01100000; // 1501 :  96 - 0x60
      11'h5DE: dout  = 8'b01111111; // 1502 : 127 - 0x7f
      11'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Background 0xbc
      11'h5E1: dout  = 8'b00100010; // 1505 :  34 - 0x22
      11'h5E2: dout  = 8'b01100101; // 1506 : 101 - 0x65
      11'h5E3: dout  = 8'b00100101; // 1507 :  37 - 0x25
      11'h5E4: dout  = 8'b00100101; // 1508 :  37 - 0x25
      11'h5E5: dout  = 8'b01110010; // 1509 : 114 - 0x72
      11'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      11'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- Background 0xbd
      11'h5E9: dout  = 8'b01110010; // 1513 : 114 - 0x72
      11'h5EA: dout  = 8'b01000101; // 1514 :  69 - 0x45
      11'h5EB: dout  = 8'b01100101; // 1515 : 101 - 0x65
      11'h5EC: dout  = 8'b00010101; // 1516 :  21 - 0x15
      11'h5ED: dout  = 8'b01100010; // 1517 :  98 - 0x62
      11'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Background 0xbe
      11'h5F1: dout  = 8'b01100111; // 1521 : 103 - 0x67
      11'h5F2: dout  = 8'b01010010; // 1522 :  82 - 0x52
      11'h5F3: dout  = 8'b01100010; // 1523 :  98 - 0x62
      11'h5F4: dout  = 8'b01000010; // 1524 :  66 - 0x42
      11'h5F5: dout  = 8'b01000010; // 1525 :  66 - 0x42
      11'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      11'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Background 0xbf
      11'h5F9: dout  = 8'b01100000; // 1529 :  96 - 0x60
      11'h5FA: dout  = 8'b10000000; // 1530 : 128 - 0x80
      11'h5FB: dout  = 8'b01000000; // 1531 :  64 - 0x40
      11'h5FC: dout  = 8'b00100000; // 1532 :  32 - 0x20
      11'h5FD: dout  = 8'b11000110; // 1533 : 198 - 0xc6
      11'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout  = 8'b01100011; // 1536 :  99 - 0x63 -- Background 0xc0
      11'h601: dout  = 8'b01100110; // 1537 : 102 - 0x66
      11'h602: dout  = 8'b01101100; // 1538 : 108 - 0x6c
      11'h603: dout  = 8'b01111000; // 1539 : 120 - 0x78
      11'h604: dout  = 8'b01111100; // 1540 : 124 - 0x7c
      11'h605: dout  = 8'b01100110; // 1541 : 102 - 0x66
      11'h606: dout  = 8'b01100011; // 1542 :  99 - 0x63
      11'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout  = 8'b00111111; // 1544 :  63 - 0x3f -- Background 0xc1
      11'h609: dout  = 8'b00001100; // 1545 :  12 - 0xc
      11'h60A: dout  = 8'b00001100; // 1546 :  12 - 0xc
      11'h60B: dout  = 8'b00001100; // 1547 :  12 - 0xc
      11'h60C: dout  = 8'b00001100; // 1548 :  12 - 0xc
      11'h60D: dout  = 8'b00001100; // 1549 :  12 - 0xc
      11'h60E: dout  = 8'b00111111; // 1550 :  63 - 0x3f
      11'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout  = 8'b01100011; // 1552 :  99 - 0x63 -- Background 0xc2
      11'h611: dout  = 8'b01110111; // 1553 : 119 - 0x77
      11'h612: dout  = 8'b01111111; // 1554 : 127 - 0x7f
      11'h613: dout  = 8'b01111111; // 1555 : 127 - 0x7f
      11'h614: dout  = 8'b01101011; // 1556 : 107 - 0x6b
      11'h615: dout  = 8'b01100011; // 1557 :  99 - 0x63
      11'h616: dout  = 8'b01100011; // 1558 :  99 - 0x63
      11'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout  = 8'b00011100; // 1560 :  28 - 0x1c -- Background 0xc3
      11'h619: dout  = 8'b00110110; // 1561 :  54 - 0x36
      11'h61A: dout  = 8'b01100011; // 1562 :  99 - 0x63
      11'h61B: dout  = 8'b01100011; // 1563 :  99 - 0x63
      11'h61C: dout  = 8'b01111111; // 1564 : 127 - 0x7f
      11'h61D: dout  = 8'b01100011; // 1565 :  99 - 0x63
      11'h61E: dout  = 8'b01100011; // 1566 :  99 - 0x63
      11'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout  = 8'b00011111; // 1568 :  31 - 0x1f -- Background 0xc4
      11'h621: dout  = 8'b00110000; // 1569 :  48 - 0x30
      11'h622: dout  = 8'b01100000; // 1570 :  96 - 0x60
      11'h623: dout  = 8'b01100111; // 1571 : 103 - 0x67
      11'h624: dout  = 8'b01100011; // 1572 :  99 - 0x63
      11'h625: dout  = 8'b00110011; // 1573 :  51 - 0x33
      11'h626: dout  = 8'b00011111; // 1574 :  31 - 0x1f
      11'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout  = 8'b01100011; // 1576 :  99 - 0x63 -- Background 0xc5
      11'h629: dout  = 8'b01100011; // 1577 :  99 - 0x63
      11'h62A: dout  = 8'b01100011; // 1578 :  99 - 0x63
      11'h62B: dout  = 8'b01100011; // 1579 :  99 - 0x63
      11'h62C: dout  = 8'b01100011; // 1580 :  99 - 0x63
      11'h62D: dout  = 8'b01100011; // 1581 :  99 - 0x63
      11'h62E: dout  = 8'b00111110; // 1582 :  62 - 0x3e
      11'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout  = 8'b01111110; // 1584 : 126 - 0x7e -- Background 0xc6
      11'h631: dout  = 8'b01100011; // 1585 :  99 - 0x63
      11'h632: dout  = 8'b01100011; // 1586 :  99 - 0x63
      11'h633: dout  = 8'b01100111; // 1587 : 103 - 0x67
      11'h634: dout  = 8'b01111100; // 1588 : 124 - 0x7c
      11'h635: dout  = 8'b01101110; // 1589 : 110 - 0x6e
      11'h636: dout  = 8'b01100111; // 1590 : 103 - 0x67
      11'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout  = 8'b01111111; // 1592 : 127 - 0x7f -- Background 0xc7
      11'h639: dout  = 8'b01100000; // 1593 :  96 - 0x60
      11'h63A: dout  = 8'b01100000; // 1594 :  96 - 0x60
      11'h63B: dout  = 8'b01111110; // 1595 : 126 - 0x7e
      11'h63C: dout  = 8'b01100000; // 1596 :  96 - 0x60
      11'h63D: dout  = 8'b01100000; // 1597 :  96 - 0x60
      11'h63E: dout  = 8'b01111111; // 1598 : 127 - 0x7f
      11'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout  = 8'b00110110; // 1600 :  54 - 0x36 -- Background 0xc8
      11'h641: dout  = 8'b00110110; // 1601 :  54 - 0x36
      11'h642: dout  = 8'b00010010; // 1602 :  18 - 0x12
      11'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout  = 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout  = 8'b00111110; // 1608 :  62 - 0x3e -- Background 0xc9
      11'h649: dout  = 8'b01100011; // 1609 :  99 - 0x63
      11'h64A: dout  = 8'b01100011; // 1610 :  99 - 0x63
      11'h64B: dout  = 8'b01100011; // 1611 :  99 - 0x63
      11'h64C: dout  = 8'b01100011; // 1612 :  99 - 0x63
      11'h64D: dout  = 8'b01100011; // 1613 :  99 - 0x63
      11'h64E: dout  = 8'b00111110; // 1614 :  62 - 0x3e
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b00111100; // 1616 :  60 - 0x3c -- Background 0xca
      11'h651: dout  = 8'b01100110; // 1617 : 102 - 0x66
      11'h652: dout  = 8'b01100000; // 1618 :  96 - 0x60
      11'h653: dout  = 8'b00111110; // 1619 :  62 - 0x3e
      11'h654: dout  = 8'b00000011; // 1620 :   3 - 0x3
      11'h655: dout  = 8'b01100011; // 1621 :  99 - 0x63
      11'h656: dout  = 8'b00111110; // 1622 :  62 - 0x3e
      11'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      11'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- Background 0xcb
      11'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      11'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      11'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      11'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      11'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      11'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Background 0xcc
      11'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      11'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      11'h665: dout  = 8'b00000000; // 1637 :   0 - 0x0
      11'h666: dout  = 8'b00000000; // 1638 :   0 - 0x0
      11'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Background 0xcd
      11'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout  = 8'b00000000; // 1643 :   0 - 0x0
      11'h66C: dout  = 8'b00000000; // 1644 :   0 - 0x0
      11'h66D: dout  = 8'b00000000; // 1645 :   0 - 0x0
      11'h66E: dout  = 8'b00000000; // 1646 :   0 - 0x0
      11'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      11'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Background 0xce
      11'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      11'h676: dout  = 8'b00000000; // 1654 :   0 - 0x0
      11'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      11'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- Background 0xcf
      11'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      11'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout  = 8'b01000111; // 1664 :  71 - 0x47 -- Background 0xd0
      11'h681: dout  = 8'b01000111; // 1665 :  71 - 0x47
      11'h682: dout  = 8'b00001111; // 1666 :  15 - 0xf
      11'h683: dout  = 8'b00001111; // 1667 :  15 - 0xf
      11'h684: dout  = 8'b00011111; // 1668 :  31 - 0x1f
      11'h685: dout  = 8'b00011111; // 1669 :  31 - 0x1f
      11'h686: dout  = 8'b00111111; // 1670 :  63 - 0x3f
      11'h687: dout  = 8'b00111111; // 1671 :  63 - 0x3f
      11'h688: dout  = 8'b11111111; // 1672 : 255 - 0xff -- Background 0xd1
      11'h689: dout  = 8'b11001111; // 1673 : 207 - 0xcf
      11'h68A: dout  = 8'b11001111; // 1674 : 207 - 0xcf
      11'h68B: dout  = 8'b11111011; // 1675 : 251 - 0xfb
      11'h68C: dout  = 8'b11110111; // 1676 : 247 - 0xf7
      11'h68D: dout  = 8'b11100111; // 1677 : 231 - 0xe7
      11'h68E: dout  = 8'b11111111; // 1678 : 255 - 0xff
      11'h68F: dout  = 8'b11111111; // 1679 : 255 - 0xff
      11'h690: dout  = 8'b00011000; // 1680 :  24 - 0x18 -- Background 0xd2
      11'h691: dout  = 8'b00001000; // 1681 :   8 - 0x8
      11'h692: dout  = 8'b10001000; // 1682 : 136 - 0x88
      11'h693: dout  = 8'b10000000; // 1683 : 128 - 0x80
      11'h694: dout  = 8'b01000000; // 1684 :  64 - 0x40
      11'h695: dout  = 8'b01000000; // 1685 :  64 - 0x40
      11'h696: dout  = 8'b10100000; // 1686 : 160 - 0xa0
      11'h697: dout  = 8'b10100000; // 1687 : 160 - 0xa0
      11'h698: dout  = 8'b11111111; // 1688 : 255 - 0xff -- Background 0xd3
      11'h699: dout  = 8'b11111111; // 1689 : 255 - 0xff
      11'h69A: dout  = 8'b11111111; // 1690 : 255 - 0xff
      11'h69B: dout  = 8'b11111111; // 1691 : 255 - 0xff
      11'h69C: dout  = 8'b11111101; // 1692 : 253 - 0xfd
      11'h69D: dout  = 8'b11111101; // 1693 : 253 - 0xfd
      11'h69E: dout  = 8'b11111101; // 1694 : 253 - 0xfd
      11'h69F: dout  = 8'b11111101; // 1695 : 253 - 0xfd
      11'h6A0: dout  = 8'b11000111; // 1696 : 199 - 0xc7 -- Background 0xd4
      11'h6A1: dout  = 8'b11110111; // 1697 : 247 - 0xf7
      11'h6A2: dout  = 8'b11110000; // 1698 : 240 - 0xf0
      11'h6A3: dout  = 8'b11111000; // 1699 : 248 - 0xf8
      11'h6A4: dout  = 8'b11111000; // 1700 : 248 - 0xf8
      11'h6A5: dout  = 8'b11111111; // 1701 : 255 - 0xff
      11'h6A6: dout  = 8'b11111111; // 1702 : 255 - 0xff
      11'h6A7: dout  = 8'b11111111; // 1703 : 255 - 0xff
      11'h6A8: dout  = 8'b11111000; // 1704 : 248 - 0xf8 -- Background 0xd5
      11'h6A9: dout  = 8'b11111000; // 1705 : 248 - 0xf8
      11'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      11'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      11'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      11'h6AD: dout  = 8'b11111111; // 1709 : 255 - 0xff
      11'h6AE: dout  = 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout  = 8'b11111111; // 1711 : 255 - 0xff
      11'h6B0: dout  = 8'b10001111; // 1712 : 143 - 0x8f -- Background 0xd6
      11'h6B1: dout  = 8'b11101111; // 1713 : 239 - 0xef
      11'h6B2: dout  = 8'b11000000; // 1714 : 192 - 0xc0
      11'h6B3: dout  = 8'b11110000; // 1715 : 240 - 0xf0
      11'h6B4: dout  = 8'b11100000; // 1716 : 224 - 0xe0
      11'h6B5: dout  = 8'b11111111; // 1717 : 255 - 0xff
      11'h6B6: dout  = 8'b11111111; // 1718 : 255 - 0xff
      11'h6B7: dout  = 8'b11111111; // 1719 : 255 - 0xff
      11'h6B8: dout  = 8'b11111111; // 1720 : 255 - 0xff -- Background 0xd7
      11'h6B9: dout  = 8'b11111111; // 1721 : 255 - 0xff
      11'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      11'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      11'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      11'h6BD: dout  = 8'b11111111; // 1725 : 255 - 0xff
      11'h6BE: dout  = 8'b11111111; // 1726 : 255 - 0xff
      11'h6BF: dout  = 8'b11111111; // 1727 : 255 - 0xff
      11'h6C0: dout  = 8'b11000011; // 1728 : 195 - 0xc3 -- Background 0xd8
      11'h6C1: dout  = 8'b11111111; // 1729 : 255 - 0xff
      11'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      11'h6C4: dout  = 8'b00000000; // 1732 :   0 - 0x0
      11'h6C5: dout  = 8'b11111111; // 1733 : 255 - 0xff
      11'h6C6: dout  = 8'b11111111; // 1734 : 255 - 0xff
      11'h6C7: dout  = 8'b11111111; // 1735 : 255 - 0xff
      11'h6C8: dout  = 8'b00000011; // 1736 :   3 - 0x3 -- Background 0xd9
      11'h6C9: dout  = 8'b10000001; // 1737 : 129 - 0x81
      11'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      11'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      11'h6CC: dout  = 8'b00000011; // 1740 :   3 - 0x3
      11'h6CD: dout  = 8'b11111111; // 1741 : 255 - 0xff
      11'h6CE: dout  = 8'b11111111; // 1742 : 255 - 0xff
      11'h6CF: dout  = 8'b11111111; // 1743 : 255 - 0xff
      11'h6D0: dout  = 8'b11111111; // 1744 : 255 - 0xff -- Background 0xda
      11'h6D1: dout  = 8'b11111111; // 1745 : 255 - 0xff
      11'h6D2: dout  = 8'b01111110; // 1746 : 126 - 0x7e
      11'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      11'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout  = 8'b11100000; // 1749 : 224 - 0xe0
      11'h6D6: dout  = 8'b11111111; // 1750 : 255 - 0xff
      11'h6D7: dout  = 8'b11111111; // 1751 : 255 - 0xff
      11'h6D8: dout  = 8'b01100001; // 1752 :  97 - 0x61 -- Background 0xdb
      11'h6D9: dout  = 8'b11000011; // 1753 : 195 - 0xc3
      11'h6DA: dout  = 8'b00000111; // 1754 :   7 - 0x7
      11'h6DB: dout  = 8'b00001111; // 1755 :  15 - 0xf
      11'h6DC: dout  = 8'b00011111; // 1756 :  31 - 0x1f
      11'h6DD: dout  = 8'b01111111; // 1757 : 127 - 0x7f
      11'h6DE: dout  = 8'b11111111; // 1758 : 255 - 0xff
      11'h6DF: dout  = 8'b11111111; // 1759 : 255 - 0xff
      11'h6E0: dout  = 8'b00011111; // 1760 :  31 - 0x1f -- Background 0xdc
      11'h6E1: dout  = 8'b11011111; // 1761 : 223 - 0xdf
      11'h6E2: dout  = 8'b11000000; // 1762 : 192 - 0xc0
      11'h6E3: dout  = 8'b11110000; // 1763 : 240 - 0xf0
      11'h6E4: dout  = 8'b11110000; // 1764 : 240 - 0xf0
      11'h6E5: dout  = 8'b11111111; // 1765 : 255 - 0xff
      11'h6E6: dout  = 8'b11111111; // 1766 : 255 - 0xff
      11'h6E7: dout  = 8'b11111111; // 1767 : 255 - 0xff
      11'h6E8: dout  = 8'b10000100; // 1768 : 132 - 0x84 -- Background 0xdd
      11'h6E9: dout  = 8'b11111100; // 1769 : 252 - 0xfc
      11'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      11'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      11'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      11'h6ED: dout  = 8'b11111111; // 1773 : 255 - 0xff
      11'h6EE: dout  = 8'b11111111; // 1774 : 255 - 0xff
      11'h6EF: dout  = 8'b11111111; // 1775 : 255 - 0xff
      11'h6F0: dout  = 8'b01111111; // 1776 : 127 - 0x7f -- Background 0xde
      11'h6F1: dout  = 8'b01111111; // 1777 : 127 - 0x7f
      11'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      11'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      11'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      11'h6F5: dout  = 8'b11111111; // 1781 : 255 - 0xff
      11'h6F6: dout  = 8'b11111111; // 1782 : 255 - 0xff
      11'h6F7: dout  = 8'b11111111; // 1783 : 255 - 0xff
      11'h6F8: dout  = 8'b11111100; // 1784 : 252 - 0xfc -- Background 0xdf
      11'h6F9: dout  = 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      11'h6FB: dout  = 8'b00000000; // 1787 :   0 - 0x0
      11'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      11'h6FD: dout  = 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout  = 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout  = 8'b11111111; // 1791 : 255 - 0xff
      11'h700: dout  = 8'b00110000; // 1792 :  48 - 0x30 -- Background 0xe0
      11'h701: dout  = 8'b11110000; // 1793 : 240 - 0xf0
      11'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      11'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      11'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      11'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout  = 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout  = 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Background 0xe1
      11'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      11'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout  = 8'b11111111; // 1805 : 255 - 0xff
      11'h70E: dout  = 8'b11111111; // 1806 : 255 - 0xff
      11'h70F: dout  = 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout  = 8'b11100001; // 1808 : 225 - 0xe1 -- Background 0xe2
      11'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      11'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      11'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout  = 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout  = 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout  = 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout  = 8'b00011111; // 1816 :  31 - 0x1f -- Background 0xe3
      11'h719: dout  = 8'b00011111; // 1817 :  31 - 0x1f
      11'h71A: dout  = 8'b00011111; // 1818 :  31 - 0x1f
      11'h71B: dout  = 8'b00011111; // 1819 :  31 - 0x1f
      11'h71C: dout  = 8'b00011111; // 1820 :  31 - 0x1f
      11'h71D: dout  = 8'b11111111; // 1821 : 255 - 0xff
      11'h71E: dout  = 8'b11111111; // 1822 : 255 - 0xff
      11'h71F: dout  = 8'b11111111; // 1823 : 255 - 0xff
      11'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Background 0xe4
      11'h721: dout  = 8'b00011111; // 1825 :  31 - 0x1f
      11'h722: dout  = 8'b00111111; // 1826 :  63 - 0x3f
      11'h723: dout  = 8'b01111000; // 1827 : 120 - 0x78
      11'h724: dout  = 8'b01110111; // 1828 : 119 - 0x77
      11'h725: dout  = 8'b01101111; // 1829 : 111 - 0x6f
      11'h726: dout  = 8'b01101111; // 1830 : 111 - 0x6f
      11'h727: dout  = 8'b01101111; // 1831 : 111 - 0x6f
      11'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Background 0xe5
      11'h729: dout  = 8'b11111000; // 1833 : 248 - 0xf8
      11'h72A: dout  = 8'b11111100; // 1834 : 252 - 0xfc
      11'h72B: dout  = 8'b00011110; // 1835 :  30 - 0x1e
      11'h72C: dout  = 8'b11101110; // 1836 : 238 - 0xee
      11'h72D: dout  = 8'b11110110; // 1837 : 246 - 0xf6
      11'h72E: dout  = 8'b11110110; // 1838 : 246 - 0xf6
      11'h72F: dout  = 8'b11110110; // 1839 : 246 - 0xf6
      11'h730: dout  = 8'b11110110; // 1840 : 246 - 0xf6 -- Background 0xe6
      11'h731: dout  = 8'b11110110; // 1841 : 246 - 0xf6
      11'h732: dout  = 8'b11110110; // 1842 : 246 - 0xf6
      11'h733: dout  = 8'b11101110; // 1843 : 238 - 0xee
      11'h734: dout  = 8'b00011110; // 1844 :  30 - 0x1e
      11'h735: dout  = 8'b11111100; // 1845 : 252 - 0xfc
      11'h736: dout  = 8'b11111000; // 1846 : 248 - 0xf8
      11'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout  = 8'b01101111; // 1848 : 111 - 0x6f -- Background 0xe7
      11'h739: dout  = 8'b01101111; // 1849 : 111 - 0x6f
      11'h73A: dout  = 8'b01101111; // 1850 : 111 - 0x6f
      11'h73B: dout  = 8'b01110111; // 1851 : 119 - 0x77
      11'h73C: dout  = 8'b01111000; // 1852 : 120 - 0x78
      11'h73D: dout  = 8'b00111111; // 1853 :  63 - 0x3f
      11'h73E: dout  = 8'b00011111; // 1854 :  31 - 0x1f
      11'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Background 0xe8
      11'h741: dout  = 8'b11111111; // 1857 : 255 - 0xff
      11'h742: dout  = 8'b11111111; // 1858 : 255 - 0xff
      11'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout  = 8'b11111111; // 1860 : 255 - 0xff
      11'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout  = 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout  = 8'b11110110; // 1864 : 246 - 0xf6 -- Background 0xe9
      11'h749: dout  = 8'b11110110; // 1865 : 246 - 0xf6
      11'h74A: dout  = 8'b11110110; // 1866 : 246 - 0xf6
      11'h74B: dout  = 8'b11110110; // 1867 : 246 - 0xf6
      11'h74C: dout  = 8'b11110110; // 1868 : 246 - 0xf6
      11'h74D: dout  = 8'b11110110; // 1869 : 246 - 0xf6
      11'h74E: dout  = 8'b11110110; // 1870 : 246 - 0xf6
      11'h74F: dout  = 8'b11110110; // 1871 : 246 - 0xf6
      11'h750: dout  = 8'b11111111; // 1872 : 255 - 0xff -- Background 0xea
      11'h751: dout  = 8'b11111111; // 1873 : 255 - 0xff
      11'h752: dout  = 8'b11111111; // 1874 : 255 - 0xff
      11'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      11'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout  = 8'b11111111; // 1877 : 255 - 0xff
      11'h756: dout  = 8'b11111111; // 1878 : 255 - 0xff
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b01101111; // 1880 : 111 - 0x6f -- Background 0xeb
      11'h759: dout  = 8'b01101111; // 1881 : 111 - 0x6f
      11'h75A: dout  = 8'b01101111; // 1882 : 111 - 0x6f
      11'h75B: dout  = 8'b01101111; // 1883 : 111 - 0x6f
      11'h75C: dout  = 8'b01101111; // 1884 : 111 - 0x6f
      11'h75D: dout  = 8'b01101111; // 1885 : 111 - 0x6f
      11'h75E: dout  = 8'b01101111; // 1886 : 111 - 0x6f
      11'h75F: dout  = 8'b01101111; // 1887 : 111 - 0x6f
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Background 0xec
      11'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      11'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0 -- Background 0xed
      11'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      11'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      11'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      11'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Background 0xee
      11'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      11'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      11'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- Background 0xef
      11'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      11'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Background 0xf0
      11'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      11'h782: dout  = 8'b11111111; // 1922 : 255 - 0xff
      11'h783: dout  = 8'b11111111; // 1923 : 255 - 0xff
      11'h784: dout  = 8'b11111111; // 1924 : 255 - 0xff
      11'h785: dout  = 8'b11111111; // 1925 : 255 - 0xff
      11'h786: dout  = 8'b11111111; // 1926 : 255 - 0xff
      11'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      11'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- Background 0xf1
      11'h789: dout  = 8'b11111111; // 1929 : 255 - 0xff
      11'h78A: dout  = 8'b11111111; // 1930 : 255 - 0xff
      11'h78B: dout  = 8'b11111111; // 1931 : 255 - 0xff
      11'h78C: dout  = 8'b11111111; // 1932 : 255 - 0xff
      11'h78D: dout  = 8'b11111111; // 1933 : 255 - 0xff
      11'h78E: dout  = 8'b11111111; // 1934 : 255 - 0xff
      11'h78F: dout  = 8'b11111111; // 1935 : 255 - 0xff
      11'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Background 0xf2
      11'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      11'h792: dout  = 8'b11111111; // 1938 : 255 - 0xff
      11'h793: dout  = 8'b11111111; // 1939 : 255 - 0xff
      11'h794: dout  = 8'b11111111; // 1940 : 255 - 0xff
      11'h795: dout  = 8'b11111111; // 1941 : 255 - 0xff
      11'h796: dout  = 8'b11111111; // 1942 : 255 - 0xff
      11'h797: dout  = 8'b11111111; // 1943 : 255 - 0xff
      11'h798: dout  = 8'b11111111; // 1944 : 255 - 0xff -- Background 0xf3
      11'h799: dout  = 8'b11111111; // 1945 : 255 - 0xff
      11'h79A: dout  = 8'b11111111; // 1946 : 255 - 0xff
      11'h79B: dout  = 8'b11111111; // 1947 : 255 - 0xff
      11'h79C: dout  = 8'b11111111; // 1948 : 255 - 0xff
      11'h79D: dout  = 8'b11111111; // 1949 : 255 - 0xff
      11'h79E: dout  = 8'b11111111; // 1950 : 255 - 0xff
      11'h79F: dout  = 8'b11111111; // 1951 : 255 - 0xff
      11'h7A0: dout  = 8'b11111111; // 1952 : 255 - 0xff -- Background 0xf4
      11'h7A1: dout  = 8'b11111111; // 1953 : 255 - 0xff
      11'h7A2: dout  = 8'b11111111; // 1954 : 255 - 0xff
      11'h7A3: dout  = 8'b11111111; // 1955 : 255 - 0xff
      11'h7A4: dout  = 8'b11111111; // 1956 : 255 - 0xff
      11'h7A5: dout  = 8'b11111111; // 1957 : 255 - 0xff
      11'h7A6: dout  = 8'b11111111; // 1958 : 255 - 0xff
      11'h7A7: dout  = 8'b11111111; // 1959 : 255 - 0xff
      11'h7A8: dout  = 8'b11111111; // 1960 : 255 - 0xff -- Background 0xf5
      11'h7A9: dout  = 8'b11111111; // 1961 : 255 - 0xff
      11'h7AA: dout  = 8'b11111111; // 1962 : 255 - 0xff
      11'h7AB: dout  = 8'b11111111; // 1963 : 255 - 0xff
      11'h7AC: dout  = 8'b11111111; // 1964 : 255 - 0xff
      11'h7AD: dout  = 8'b11111111; // 1965 : 255 - 0xff
      11'h7AE: dout  = 8'b11111111; // 1966 : 255 - 0xff
      11'h7AF: dout  = 8'b11111111; // 1967 : 255 - 0xff
      11'h7B0: dout  = 8'b11111111; // 1968 : 255 - 0xff -- Background 0xf6
      11'h7B1: dout  = 8'b11111111; // 1969 : 255 - 0xff
      11'h7B2: dout  = 8'b11111111; // 1970 : 255 - 0xff
      11'h7B3: dout  = 8'b11111111; // 1971 : 255 - 0xff
      11'h7B4: dout  = 8'b11111111; // 1972 : 255 - 0xff
      11'h7B5: dout  = 8'b11111111; // 1973 : 255 - 0xff
      11'h7B6: dout  = 8'b11111111; // 1974 : 255 - 0xff
      11'h7B7: dout  = 8'b11111111; // 1975 : 255 - 0xff
      11'h7B8: dout  = 8'b11111111; // 1976 : 255 - 0xff -- Background 0xf7
      11'h7B9: dout  = 8'b11111111; // 1977 : 255 - 0xff
      11'h7BA: dout  = 8'b11111111; // 1978 : 255 - 0xff
      11'h7BB: dout  = 8'b11111111; // 1979 : 255 - 0xff
      11'h7BC: dout  = 8'b11111111; // 1980 : 255 - 0xff
      11'h7BD: dout  = 8'b11111111; // 1981 : 255 - 0xff
      11'h7BE: dout  = 8'b11111111; // 1982 : 255 - 0xff
      11'h7BF: dout  = 8'b11111111; // 1983 : 255 - 0xff
      11'h7C0: dout  = 8'b11111111; // 1984 : 255 - 0xff -- Background 0xf8
      11'h7C1: dout  = 8'b11111111; // 1985 : 255 - 0xff
      11'h7C2: dout  = 8'b11111111; // 1986 : 255 - 0xff
      11'h7C3: dout  = 8'b11111111; // 1987 : 255 - 0xff
      11'h7C4: dout  = 8'b11111111; // 1988 : 255 - 0xff
      11'h7C5: dout  = 8'b11111111; // 1989 : 255 - 0xff
      11'h7C6: dout  = 8'b11111111; // 1990 : 255 - 0xff
      11'h7C7: dout  = 8'b11111111; // 1991 : 255 - 0xff
      11'h7C8: dout  = 8'b11111111; // 1992 : 255 - 0xff -- Background 0xf9
      11'h7C9: dout  = 8'b11111111; // 1993 : 255 - 0xff
      11'h7CA: dout  = 8'b11111111; // 1994 : 255 - 0xff
      11'h7CB: dout  = 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout  = 8'b11111111; // 1996 : 255 - 0xff
      11'h7CD: dout  = 8'b11111111; // 1997 : 255 - 0xff
      11'h7CE: dout  = 8'b11111111; // 1998 : 255 - 0xff
      11'h7CF: dout  = 8'b11111111; // 1999 : 255 - 0xff
      11'h7D0: dout  = 8'b11111111; // 2000 : 255 - 0xff -- Background 0xfa
      11'h7D1: dout  = 8'b11111111; // 2001 : 255 - 0xff
      11'h7D2: dout  = 8'b11111111; // 2002 : 255 - 0xff
      11'h7D3: dout  = 8'b11111111; // 2003 : 255 - 0xff
      11'h7D4: dout  = 8'b11111111; // 2004 : 255 - 0xff
      11'h7D5: dout  = 8'b11111111; // 2005 : 255 - 0xff
      11'h7D6: dout  = 8'b11111111; // 2006 : 255 - 0xff
      11'h7D7: dout  = 8'b11111111; // 2007 : 255 - 0xff
      11'h7D8: dout  = 8'b11111111; // 2008 : 255 - 0xff -- Background 0xfb
      11'h7D9: dout  = 8'b11111111; // 2009 : 255 - 0xff
      11'h7DA: dout  = 8'b11111111; // 2010 : 255 - 0xff
      11'h7DB: dout  = 8'b11111111; // 2011 : 255 - 0xff
      11'h7DC: dout  = 8'b11111111; // 2012 : 255 - 0xff
      11'h7DD: dout  = 8'b11111111; // 2013 : 255 - 0xff
      11'h7DE: dout  = 8'b11111111; // 2014 : 255 - 0xff
      11'h7DF: dout  = 8'b11111111; // 2015 : 255 - 0xff
      11'h7E0: dout  = 8'b11111111; // 2016 : 255 - 0xff -- Background 0xfc
      11'h7E1: dout  = 8'b11111111; // 2017 : 255 - 0xff
      11'h7E2: dout  = 8'b11111111; // 2018 : 255 - 0xff
      11'h7E3: dout  = 8'b11111111; // 2019 : 255 - 0xff
      11'h7E4: dout  = 8'b11111111; // 2020 : 255 - 0xff
      11'h7E5: dout  = 8'b11111111; // 2021 : 255 - 0xff
      11'h7E6: dout  = 8'b11111111; // 2022 : 255 - 0xff
      11'h7E7: dout  = 8'b11111111; // 2023 : 255 - 0xff
      11'h7E8: dout  = 8'b11111111; // 2024 : 255 - 0xff -- Background 0xfd
      11'h7E9: dout  = 8'b11111111; // 2025 : 255 - 0xff
      11'h7EA: dout  = 8'b11111111; // 2026 : 255 - 0xff
      11'h7EB: dout  = 8'b11111111; // 2027 : 255 - 0xff
      11'h7EC: dout  = 8'b11111111; // 2028 : 255 - 0xff
      11'h7ED: dout  = 8'b11111111; // 2029 : 255 - 0xff
      11'h7EE: dout  = 8'b11111111; // 2030 : 255 - 0xff
      11'h7EF: dout  = 8'b11111111; // 2031 : 255 - 0xff
      11'h7F0: dout  = 8'b11111111; // 2032 : 255 - 0xff -- Background 0xfe
      11'h7F1: dout  = 8'b11111111; // 2033 : 255 - 0xff
      11'h7F2: dout  = 8'b11111111; // 2034 : 255 - 0xff
      11'h7F3: dout  = 8'b11111111; // 2035 : 255 - 0xff
      11'h7F4: dout  = 8'b11111111; // 2036 : 255 - 0xff
      11'h7F5: dout  = 8'b11111111; // 2037 : 255 - 0xff
      11'h7F6: dout  = 8'b11111111; // 2038 : 255 - 0xff
      11'h7F7: dout  = 8'b11111111; // 2039 : 255 - 0xff
      11'h7F8: dout  = 8'b11111111; // 2040 : 255 - 0xff -- Background 0xff
      11'h7F9: dout  = 8'b11111111; // 2041 : 255 - 0xff
      11'h7FA: dout  = 8'b11111111; // 2042 : 255 - 0xff
      11'h7FB: dout  = 8'b11111111; // 2043 : 255 - 0xff
      11'h7FC: dout  = 8'b11111111; // 2044 : 255 - 0xff
      11'h7FD: dout  = 8'b11111111; // 2045 : 255 - 0xff
      11'h7FE: dout  = 8'b11111111; // 2046 : 255 - 0xff
      11'h7FF: dout  = 8'b11111111; // 2047 : 255 - 0xff
    endcase
  end

endmodule
