//- Autcmatically generated verilog ROM from a NES memory file----
//-   ATTRIBUTE TABLE SEPARATED FROM NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_attribute_tables


//-  Original memory dump file name: smario_ntable_01.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_ATABLE_SMARIO_01
  (
     //input     clk,   // clock
     input      [7-1:0] addr,  //128 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
      7'h0: dout  = 8'b10101010; //    0 : 170 - 0xaa
      7'h1: dout  = 8'b10101010; //    1 : 170 - 0xaa
      7'h2: dout  = 8'b11101010; //    2 : 234 - 0xea
      7'h3: dout  = 8'b10101010; //    3 : 170 - 0xaa
      7'h4: dout  = 8'b10101010; //    4 : 170 - 0xaa
      7'h5: dout  = 8'b10101010; //    5 : 170 - 0xaa
      7'h6: dout  = 8'b10101010; //    6 : 170 - 0xaa
      7'h7: dout  = 8'b10101010; //    7 : 170 - 0xaa
      7'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      7'h9: dout  = 8'b01010101; //    9 :  85 - 0x55
      7'hA: dout  = 8'b01010101; //   10 :  85 - 0x55
      7'hB: dout  = 8'b01010101; //   11 :  85 - 0x55
      7'hC: dout  = 8'b01010101; //   12 :  85 - 0x55
      7'hD: dout  = 8'b01010101; //   13 :  85 - 0x55
      7'hE: dout  = 8'b01010101; //   14 :  85 - 0x55
      7'hF: dout  = 8'b01010101; //   15 :  85 - 0x55
      7'h10: dout  = 8'b01010101; //   16 :  85 - 0x55
      7'h11: dout  = 8'b01010101; //   17 :  85 - 0x55
      7'h12: dout  = 8'b01010101; //   18 :  85 - 0x55
      7'h13: dout  = 8'b01010101; //   19 :  85 - 0x55
      7'h14: dout  = 8'b01010101; //   20 :  85 - 0x55
      7'h15: dout  = 8'b01010101; //   21 :  85 - 0x55
      7'h16: dout  = 8'b01010101; //   22 :  85 - 0x55
      7'h17: dout  = 8'b01010101; //   23 :  85 - 0x55
      7'h18: dout  = 8'b01010101; //   24 :  85 - 0x55
      7'h19: dout  = 8'b01010101; //   25 :  85 - 0x55
      7'h1A: dout  = 8'b01010101; //   26 :  85 - 0x55
      7'h1B: dout  = 8'b01010101; //   27 :  85 - 0x55
      7'h1C: dout  = 8'b01010101; //   28 :  85 - 0x55
      7'h1D: dout  = 8'b01010101; //   29 :  85 - 0x55
      7'h1E: dout  = 8'b01010101; //   30 :  85 - 0x55
      7'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      7'h20: dout  = 8'b00000000; //   32 :   0 - 0x0
      7'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      7'h22: dout  = 8'b10011001; //   34 : 153 - 0x99
      7'h23: dout  = 8'b10101010; //   35 : 170 - 0xaa
      7'h24: dout  = 8'b10101010; //   36 : 170 - 0xaa
      7'h25: dout  = 8'b10101010; //   37 : 170 - 0xaa
      7'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      7'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      7'h28: dout  = 8'b00000000; //   40 :   0 - 0x0
      7'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      7'h2A: dout  = 8'b10011001; //   42 : 153 - 0x99
      7'h2B: dout  = 8'b10101010; //   43 : 170 - 0xaa
      7'h2C: dout  = 8'b10101010; //   44 : 170 - 0xaa
      7'h2D: dout  = 8'b10101010; //   45 : 170 - 0xaa
      7'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      7'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      7'h30: dout  = 8'b01010000; //   48 :  80 - 0x50
      7'h31: dout  = 8'b01010000; //   49 :  80 - 0x50
      7'h32: dout  = 8'b01010000; //   50 :  80 - 0x50
      7'h33: dout  = 8'b01010000; //   51 :  80 - 0x50
      7'h34: dout  = 8'b01010000; //   52 :  80 - 0x50
      7'h35: dout  = 8'b01010000; //   53 :  80 - 0x50
      7'h36: dout  = 8'b01010000; //   54 :  80 - 0x50
      7'h37: dout  = 8'b01010000; //   55 :  80 - 0x50
      7'h38: dout  = 8'b00000101; //   56 :   5 - 0x5
      7'h39: dout  = 8'b00000101; //   57 :   5 - 0x5
      7'h3A: dout  = 8'b00000101; //   58 :   5 - 0x5
      7'h3B: dout  = 8'b00000101; //   59 :   5 - 0x5
      7'h3C: dout  = 8'b00000101; //   60 :   5 - 0x5
      7'h3D: dout  = 8'b00000101; //   61 :   5 - 0x5
      7'h3E: dout  = 8'b00000101; //   62 :   5 - 0x5
      7'h3F: dout  = 8'b00000101; //   63 :   5 - 0x5
      7'h40: dout  = 8'b00000000; //   64 :   0 - 0x0
      7'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      7'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      7'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      7'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      7'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      7'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      7'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      7'h48: dout  = 8'b00000000; //   72 :   0 - 0x0
      7'h49: dout  = 8'b10001000; //   73 : 136 - 0x88
      7'h4A: dout  = 8'b10101010; //   74 : 170 - 0xaa
      7'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      7'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      7'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      7'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      7'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      7'h50: dout  = 8'b00000000; //   80 :   0 - 0x0
      7'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      7'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      7'h53: dout  = 8'b00110000; //   83 :  48 - 0x30
      7'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      7'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      7'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      7'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      7'h58: dout  = 8'b00000000; //   88 :   0 - 0x0
      7'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      7'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      7'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      7'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      7'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      7'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      7'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      7'h60: dout  = 8'b00110000; //   96 :  48 - 0x30
      7'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      7'h62: dout  = 8'b11010000; //   98 : 208 - 0xd0
      7'h63: dout  = 8'b11010000; //   99 : 208 - 0xd0
      7'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      7'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      7'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      7'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      7'h68: dout  = 8'b00000000; //  104 :   0 - 0x0
      7'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      7'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      7'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      7'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      7'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      7'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      7'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      7'h70: dout  = 8'b01010000; //  112 :  80 - 0x50
      7'h71: dout  = 8'b01010000; //  113 :  80 - 0x50
      7'h72: dout  = 8'b01010000; //  114 :  80 - 0x50
      7'h73: dout  = 8'b01010000; //  115 :  80 - 0x50
      7'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      7'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      7'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      7'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      7'h78: dout  = 8'b00000101; //  120 :   5 - 0x5
      7'h79: dout  = 8'b00000101; //  121 :   5 - 0x5
      7'h7A: dout  = 8'b00000101; //  122 :   5 - 0x5
      7'h7B: dout  = 8'b00000101; //  123 :   5 - 0x5
      7'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      7'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      7'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      7'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
    endcase
  end

endmodule
