//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: sprilo_racet3.bin --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE_SPRILO_RACE3
  (
     //input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout  = 8'b11111010; //    0 : 250 - 0xfa -- line 0x0
      10'h1: dout  = 8'b11111010; //    1 : 250 - 0xfa
      10'h2: dout  = 8'b11111010; //    2 : 250 - 0xfa
      10'h3: dout  = 8'b11101010; //    3 : 234 - 0xea
      10'h4: dout  = 8'b11111010; //    4 : 250 - 0xfa
      10'h5: dout  = 8'b11111010; //    5 : 250 - 0xfa
      10'h6: dout  = 8'b11111010; //    6 : 250 - 0xfa
      10'h7: dout  = 8'b11111010; //    7 : 250 - 0xfa
      10'h8: dout  = 8'b11111010; //    8 : 250 - 0xfa
      10'h9: dout  = 8'b11111010; //    9 : 250 - 0xfa
      10'hA: dout  = 8'b11111010; //   10 : 250 - 0xfa
      10'hB: dout  = 8'b11111010; //   11 : 250 - 0xfa
      10'hC: dout  = 8'b11111010; //   12 : 250 - 0xfa
      10'hD: dout  = 8'b11111010; //   13 : 250 - 0xfa
      10'hE: dout  = 8'b11101010; //   14 : 234 - 0xea
      10'hF: dout  = 8'b11111010; //   15 : 250 - 0xfa
      10'h10: dout  = 8'b11111010; //   16 : 250 - 0xfa
      10'h11: dout  = 8'b11111010; //   17 : 250 - 0xfa
      10'h12: dout  = 8'b11111010; //   18 : 250 - 0xfa
      10'h13: dout  = 8'b11111010; //   19 : 250 - 0xfa
      10'h14: dout  = 8'b11111010; //   20 : 250 - 0xfa
      10'h15: dout  = 8'b11111010; //   21 : 250 - 0xfa
      10'h16: dout  = 8'b11101001; //   22 : 233 - 0xe9
      10'h17: dout  = 8'b11111010; //   23 : 250 - 0xfa
      10'h18: dout  = 8'b11111010; //   24 : 250 - 0xfa
      10'h19: dout  = 8'b11111010; //   25 : 250 - 0xfa
      10'h1A: dout  = 8'b11111010; //   26 : 250 - 0xfa
      10'h1B: dout  = 8'b11111010; //   27 : 250 - 0xfa
      10'h1C: dout  = 8'b11101010; //   28 : 234 - 0xea
      10'h1D: dout  = 8'b11111010; //   29 : 250 - 0xfa
      10'h1E: dout  = 8'b11111010; //   30 : 250 - 0xfa
      10'h1F: dout  = 8'b11111010; //   31 : 250 - 0xfa
      10'h20: dout  = 8'b11111010; //   32 : 250 - 0xfa -- line 0x1
      10'h21: dout  = 8'b11111010; //   33 : 250 - 0xfa
      10'h22: dout  = 8'b11111010; //   34 : 250 - 0xfa
      10'h23: dout  = 8'b11100111; //   35 : 231 - 0xe7
      10'h24: dout  = 8'b11111011; //   36 : 251 - 0xfb
      10'h25: dout  = 8'b11111011; //   37 : 251 - 0xfb
      10'h26: dout  = 8'b11111011; //   38 : 251 - 0xfb
      10'h27: dout  = 8'b11111011; //   39 : 251 - 0xfb
      10'h28: dout  = 8'b11111011; //   40 : 251 - 0xfb
      10'h29: dout  = 8'b11111011; //   41 : 251 - 0xfb
      10'h2A: dout  = 8'b11111011; //   42 : 251 - 0xfb
      10'h2B: dout  = 8'b11111011; //   43 : 251 - 0xfb
      10'h2C: dout  = 8'b11111011; //   44 : 251 - 0xfb
      10'h2D: dout  = 8'b11111011; //   45 : 251 - 0xfb
      10'h2E: dout  = 8'b11111011; //   46 : 251 - 0xfb
      10'h2F: dout  = 8'b11111011; //   47 : 251 - 0xfb
      10'h30: dout  = 8'b11101000; //   48 : 232 - 0xe8
      10'h31: dout  = 8'b11111010; //   49 : 250 - 0xfa
      10'h32: dout  = 8'b11101010; //   50 : 234 - 0xea
      10'h33: dout  = 8'b11111010; //   51 : 250 - 0xfa
      10'h34: dout  = 8'b11111010; //   52 : 250 - 0xfa
      10'h35: dout  = 8'b11111010; //   53 : 250 - 0xfa
      10'h36: dout  = 8'b11111010; //   54 : 250 - 0xfa
      10'h37: dout  = 8'b11111010; //   55 : 250 - 0xfa
      10'h38: dout  = 8'b11111010; //   56 : 250 - 0xfa
      10'h39: dout  = 8'b11111001; //   57 : 249 - 0xf9
      10'h3A: dout  = 8'b11111010; //   58 : 250 - 0xfa
      10'h3B: dout  = 8'b11111010; //   59 : 250 - 0xfa
      10'h3C: dout  = 8'b11111010; //   60 : 250 - 0xfa
      10'h3D: dout  = 8'b11111010; //   61 : 250 - 0xfa
      10'h3E: dout  = 8'b11111010; //   62 : 250 - 0xfa
      10'h3F: dout  = 8'b11101010; //   63 : 234 - 0xea
      10'h40: dout  = 8'b11101010; //   64 : 234 - 0xea -- line 0x2
      10'h41: dout  = 8'b11111010; //   65 : 250 - 0xfa
      10'h42: dout  = 8'b11111010; //   66 : 250 - 0xfa
      10'h43: dout  = 8'b11111100; //   67 : 252 - 0xfc
      10'h44: dout  = 8'b11111111; //   68 : 255 - 0xff
      10'h45: dout  = 8'b11111111; //   69 : 255 - 0xff
      10'h46: dout  = 8'b11111111; //   70 : 255 - 0xff
      10'h47: dout  = 8'b11111111; //   71 : 255 - 0xff
      10'h48: dout  = 8'b11111111; //   72 : 255 - 0xff
      10'h49: dout  = 8'b11111111; //   73 : 255 - 0xff
      10'h4A: dout  = 8'b11111111; //   74 : 255 - 0xff
      10'h4B: dout  = 8'b11111111; //   75 : 255 - 0xff
      10'h4C: dout  = 8'b11111111; //   76 : 255 - 0xff
      10'h4D: dout  = 8'b11111111; //   77 : 255 - 0xff
      10'h4E: dout  = 8'b11111111; //   78 : 255 - 0xff
      10'h4F: dout  = 8'b11111111; //   79 : 255 - 0xff
      10'h50: dout  = 8'b11101100; //   80 : 236 - 0xec
      10'h51: dout  = 8'b11111010; //   81 : 250 - 0xfa
      10'h52: dout  = 8'b11111010; //   82 : 250 - 0xfa
      10'h53: dout  = 8'b11111001; //   83 : 249 - 0xf9
      10'h54: dout  = 8'b11111010; //   84 : 250 - 0xfa
      10'h55: dout  = 8'b11111010; //   85 : 250 - 0xfa
      10'h56: dout  = 8'b11101001; //   86 : 233 - 0xe9
      10'h57: dout  = 8'b11111010; //   87 : 250 - 0xfa
      10'h58: dout  = 8'b11111010; //   88 : 250 - 0xfa
      10'h59: dout  = 8'b11111010; //   89 : 250 - 0xfa
      10'h5A: dout  = 8'b11111010; //   90 : 250 - 0xfa
      10'h5B: dout  = 8'b11101010; //   91 : 234 - 0xea
      10'h5C: dout  = 8'b11111010; //   92 : 250 - 0xfa
      10'h5D: dout  = 8'b11101001; //   93 : 233 - 0xe9
      10'h5E: dout  = 8'b11111010; //   94 : 250 - 0xfa
      10'h5F: dout  = 8'b11111010; //   95 : 250 - 0xfa
      10'h60: dout  = 8'b11111010; //   96 : 250 - 0xfa -- line 0x3
      10'h61: dout  = 8'b11100111; //   97 : 231 - 0xe7
      10'h62: dout  = 8'b11111011; //   98 : 251 - 0xfb
      10'h63: dout  = 8'b11110110; //   99 : 246 - 0xf6
      10'h64: dout  = 8'b11111111; //  100 : 255 - 0xff
      10'h65: dout  = 8'b11111111; //  101 : 255 - 0xff
      10'h66: dout  = 8'b11111101; //  102 : 253 - 0xfd
      10'h67: dout  = 8'b11111111; //  103 : 255 - 0xff
      10'h68: dout  = 8'b11111101; //  104 : 253 - 0xfd
      10'h69: dout  = 8'b11111111; //  105 : 255 - 0xff
      10'h6A: dout  = 8'b11111101; //  106 : 253 - 0xfd
      10'h6B: dout  = 8'b11111111; //  107 : 255 - 0xff
      10'h6C: dout  = 8'b11111101; //  108 : 253 - 0xfd
      10'h6D: dout  = 8'b11111111; //  109 : 255 - 0xff
      10'h6E: dout  = 8'b11111111; //  110 : 255 - 0xff
      10'h6F: dout  = 8'b11111111; //  111 : 255 - 0xff
      10'h70: dout  = 8'b11101100; //  112 : 236 - 0xec
      10'h71: dout  = 8'b11111010; //  113 : 250 - 0xfa
      10'h72: dout  = 8'b11111010; //  114 : 250 - 0xfa
      10'h73: dout  = 8'b11111010; //  115 : 250 - 0xfa
      10'h74: dout  = 8'b11111010; //  116 : 250 - 0xfa
      10'h75: dout  = 8'b11111010; //  117 : 250 - 0xfa
      10'h76: dout  = 8'b11111010; //  118 : 250 - 0xfa
      10'h77: dout  = 8'b11111010; //  119 : 250 - 0xfa
      10'h78: dout  = 8'b11101001; //  120 : 233 - 0xe9
      10'h79: dout  = 8'b11111010; //  121 : 250 - 0xfa
      10'h7A: dout  = 8'b11111010; //  122 : 250 - 0xfa
      10'h7B: dout  = 8'b11111010; //  123 : 250 - 0xfa
      10'h7C: dout  = 8'b11111010; //  124 : 250 - 0xfa
      10'h7D: dout  = 8'b11111010; //  125 : 250 - 0xfa
      10'h7E: dout  = 8'b11111010; //  126 : 250 - 0xfa
      10'h7F: dout  = 8'b11111010; //  127 : 250 - 0xfa
      10'h80: dout  = 8'b11101001; //  128 : 233 - 0xe9 -- line 0x4
      10'h81: dout  = 8'b11111100; //  129 : 252 - 0xfc
      10'h82: dout  = 8'b11111111; //  130 : 255 - 0xff
      10'h83: dout  = 8'b11111111; //  131 : 255 - 0xff
      10'h84: dout  = 8'b11111111; //  132 : 255 - 0xff
      10'h85: dout  = 8'b11111111; //  133 : 255 - 0xff
      10'h86: dout  = 8'b11111101; //  134 : 253 - 0xfd
      10'h87: dout  = 8'b11111111; //  135 : 255 - 0xff
      10'h88: dout  = 8'b11111101; //  136 : 253 - 0xfd
      10'h89: dout  = 8'b11111111; //  137 : 255 - 0xff
      10'h8A: dout  = 8'b11111101; //  138 : 253 - 0xfd
      10'h8B: dout  = 8'b11111111; //  139 : 255 - 0xff
      10'h8C: dout  = 8'b11111101; //  140 : 253 - 0xfd
      10'h8D: dout  = 8'b11111111; //  141 : 255 - 0xff
      10'h8E: dout  = 8'b11111111; //  142 : 255 - 0xff
      10'h8F: dout  = 8'b11111111; //  143 : 255 - 0xff
      10'h90: dout  = 8'b11101100; //  144 : 236 - 0xec
      10'h91: dout  = 8'b11111010; //  145 : 250 - 0xfa
      10'h92: dout  = 8'b11111010; //  146 : 250 - 0xfa
      10'h93: dout  = 8'b11101001; //  147 : 233 - 0xe9
      10'h94: dout  = 8'b11111010; //  148 : 250 - 0xfa
      10'h95: dout  = 8'b11111010; //  149 : 250 - 0xfa
      10'h96: dout  = 8'b11111010; //  150 : 250 - 0xfa
      10'h97: dout  = 8'b11111010; //  151 : 250 - 0xfa
      10'h98: dout  = 8'b11111010; //  152 : 250 - 0xfa
      10'h99: dout  = 8'b11111010; //  153 : 250 - 0xfa
      10'h9A: dout  = 8'b11111010; //  154 : 250 - 0xfa
      10'h9B: dout  = 8'b11111010; //  155 : 250 - 0xfa
      10'h9C: dout  = 8'b11111010; //  156 : 250 - 0xfa
      10'h9D: dout  = 8'b11111010; //  157 : 250 - 0xfa
      10'h9E: dout  = 8'b11111010; //  158 : 250 - 0xfa
      10'h9F: dout  = 8'b11111010; //  159 : 250 - 0xfa
      10'hA0: dout  = 8'b11111010; //  160 : 250 - 0xfa -- line 0x5
      10'hA1: dout  = 8'b11111100; //  161 : 252 - 0xfc
      10'hA2: dout  = 8'b11111111; //  162 : 255 - 0xff
      10'hA3: dout  = 8'b11111111; //  163 : 255 - 0xff
      10'hA4: dout  = 8'b11111111; //  164 : 255 - 0xff
      10'hA5: dout  = 8'b11111111; //  165 : 255 - 0xff
      10'hA6: dout  = 8'b11111111; //  166 : 255 - 0xff
      10'hA7: dout  = 8'b11111111; //  167 : 255 - 0xff
      10'hA8: dout  = 8'b11111111; //  168 : 255 - 0xff
      10'hA9: dout  = 8'b11111111; //  169 : 255 - 0xff
      10'hAA: dout  = 8'b11111111; //  170 : 255 - 0xff
      10'hAB: dout  = 8'b11111111; //  171 : 255 - 0xff
      10'hAC: dout  = 8'b11111111; //  172 : 255 - 0xff
      10'hAD: dout  = 8'b11111111; //  173 : 255 - 0xff
      10'hAE: dout  = 8'b11111111; //  174 : 255 - 0xff
      10'hAF: dout  = 8'b11111111; //  175 : 255 - 0xff
      10'hB0: dout  = 8'b11101100; //  176 : 236 - 0xec
      10'hB1: dout  = 8'b11111010; //  177 : 250 - 0xfa
      10'hB2: dout  = 8'b11111010; //  178 : 250 - 0xfa
      10'hB3: dout  = 8'b11111010; //  179 : 250 - 0xfa
      10'hB4: dout  = 8'b11111010; //  180 : 250 - 0xfa
      10'hB5: dout  = 8'b11111010; //  181 : 250 - 0xfa
      10'hB6: dout  = 8'b11101010; //  182 : 234 - 0xea
      10'hB7: dout  = 8'b11111010; //  183 : 250 - 0xfa
      10'hB8: dout  = 8'b11111001; //  184 : 249 - 0xf9
      10'hB9: dout  = 8'b11111010; //  185 : 250 - 0xfa
      10'hBA: dout  = 8'b11111010; //  186 : 250 - 0xfa
      10'hBB: dout  = 8'b11101001; //  187 : 233 - 0xe9
      10'hBC: dout  = 8'b11111010; //  188 : 250 - 0xfa
      10'hBD: dout  = 8'b11111010; //  189 : 250 - 0xfa
      10'hBE: dout  = 8'b11111010; //  190 : 250 - 0xfa
      10'hBF: dout  = 8'b11111010; //  191 : 250 - 0xfa
      10'hC0: dout  = 8'b11111010; //  192 : 250 - 0xfa -- line 0x6
      10'hC1: dout  = 8'b11111100; //  193 : 252 - 0xfc
      10'hC2: dout  = 8'b11111111; //  194 : 255 - 0xff
      10'hC3: dout  = 8'b11111110; //  195 : 254 - 0xfe
      10'hC4: dout  = 8'b11111110; //  196 : 254 - 0xfe
      10'hC5: dout  = 8'b11111111; //  197 : 255 - 0xff
      10'hC6: dout  = 8'b11100101; //  198 : 229 - 0xe5
      10'hC7: dout  = 8'b11101011; //  199 : 235 - 0xeb
      10'hC8: dout  = 8'b11101011; //  200 : 235 - 0xeb
      10'hC9: dout  = 8'b11101011; //  201 : 235 - 0xeb
      10'hCA: dout  = 8'b11101011; //  202 : 235 - 0xeb
      10'hCB: dout  = 8'b11100110; //  203 : 230 - 0xe6
      10'hCC: dout  = 8'b11111111; //  204 : 255 - 0xff
      10'hCD: dout  = 8'b11111110; //  205 : 254 - 0xfe
      10'hCE: dout  = 8'b11111110; //  206 : 254 - 0xfe
      10'hCF: dout  = 8'b11111111; //  207 : 255 - 0xff
      10'hD0: dout  = 8'b11101100; //  208 : 236 - 0xec
      10'hD1: dout  = 8'b11111010; //  209 : 250 - 0xfa
      10'hD2: dout  = 8'b11111001; //  210 : 249 - 0xf9
      10'hD3: dout  = 8'b11111010; //  211 : 250 - 0xfa
      10'hD4: dout  = 8'b11111010; //  212 : 250 - 0xfa
      10'hD5: dout  = 8'b11111010; //  213 : 250 - 0xfa
      10'hD6: dout  = 8'b11111010; //  214 : 250 - 0xfa
      10'hD7: dout  = 8'b11111010; //  215 : 250 - 0xfa
      10'hD8: dout  = 8'b11111010; //  216 : 250 - 0xfa
      10'hD9: dout  = 8'b11111001; //  217 : 249 - 0xf9
      10'hDA: dout  = 8'b11111010; //  218 : 250 - 0xfa
      10'hDB: dout  = 8'b11111010; //  219 : 250 - 0xfa
      10'hDC: dout  = 8'b11111010; //  220 : 250 - 0xfa
      10'hDD: dout  = 8'b11111010; //  221 : 250 - 0xfa
      10'hDE: dout  = 8'b11111010; //  222 : 250 - 0xfa
      10'hDF: dout  = 8'b11101010; //  223 : 234 - 0xea
      10'hE0: dout  = 8'b11111010; //  224 : 250 - 0xfa -- line 0x7
      10'hE1: dout  = 8'b11111100; //  225 : 252 - 0xfc
      10'hE2: dout  = 8'b11111111; //  226 : 255 - 0xff
      10'hE3: dout  = 8'b11111111; //  227 : 255 - 0xff
      10'hE4: dout  = 8'b11111111; //  228 : 255 - 0xff
      10'hE5: dout  = 8'b11111111; //  229 : 255 - 0xff
      10'hE6: dout  = 8'b11101100; //  230 : 236 - 0xec
      10'hE7: dout  = 8'b11111010; //  231 : 250 - 0xfa
      10'hE8: dout  = 8'b11111010; //  232 : 250 - 0xfa
      10'hE9: dout  = 8'b11111010; //  233 : 250 - 0xfa
      10'hEA: dout  = 8'b11111010; //  234 : 250 - 0xfa
      10'hEB: dout  = 8'b11111100; //  235 : 252 - 0xfc
      10'hEC: dout  = 8'b11111111; //  236 : 255 - 0xff
      10'hED: dout  = 8'b11111111; //  237 : 255 - 0xff
      10'hEE: dout  = 8'b11111111; //  238 : 255 - 0xff
      10'hEF: dout  = 8'b11111111; //  239 : 255 - 0xff
      10'hF0: dout  = 8'b11101100; //  240 : 236 - 0xec
      10'hF1: dout  = 8'b11111010; //  241 : 250 - 0xfa
      10'hF2: dout  = 8'b11111010; //  242 : 250 - 0xfa
      10'hF3: dout  = 8'b11111010; //  243 : 250 - 0xfa
      10'hF4: dout  = 8'b11111010; //  244 : 250 - 0xfa
      10'hF5: dout  = 8'b11111010; //  245 : 250 - 0xfa
      10'hF6: dout  = 8'b11111010; //  246 : 250 - 0xfa
      10'hF7: dout  = 8'b11111010; //  247 : 250 - 0xfa
      10'hF8: dout  = 8'b11111010; //  248 : 250 - 0xfa
      10'hF9: dout  = 8'b11111010; //  249 : 250 - 0xfa
      10'hFA: dout  = 8'b11101010; //  250 : 234 - 0xea
      10'hFB: dout  = 8'b11111010; //  251 : 250 - 0xfa
      10'hFC: dout  = 8'b11111001; //  252 : 249 - 0xf9
      10'hFD: dout  = 8'b11111010; //  253 : 250 - 0xfa
      10'hFE: dout  = 8'b11111010; //  254 : 250 - 0xfa
      10'hFF: dout  = 8'b11111010; //  255 : 250 - 0xfa
      10'h100: dout  = 8'b11111010; //  256 : 250 - 0xfa -- line 0x8
      10'h101: dout  = 8'b11111100; //  257 : 252 - 0xfc
      10'h102: dout  = 8'b11111111; //  258 : 255 - 0xff
      10'h103: dout  = 8'b11111110; //  259 : 254 - 0xfe
      10'h104: dout  = 8'b11111110; //  260 : 254 - 0xfe
      10'h105: dout  = 8'b11111111; //  261 : 255 - 0xff
      10'h106: dout  = 8'b11101100; //  262 : 236 - 0xec
      10'h107: dout  = 8'b11111010; //  263 : 250 - 0xfa
      10'h108: dout  = 8'b11111001; //  264 : 249 - 0xf9
      10'h109: dout  = 8'b11111010; //  265 : 250 - 0xfa
      10'h10A: dout  = 8'b11111010; //  266 : 250 - 0xfa
      10'h10B: dout  = 8'b11111100; //  267 : 252 - 0xfc
      10'h10C: dout  = 8'b11111111; //  268 : 255 - 0xff
      10'h10D: dout  = 8'b11111110; //  269 : 254 - 0xfe
      10'h10E: dout  = 8'b11111110; //  270 : 254 - 0xfe
      10'h10F: dout  = 8'b11111111; //  271 : 255 - 0xff
      10'h110: dout  = 8'b11101100; //  272 : 236 - 0xec
      10'h111: dout  = 8'b11111010; //  273 : 250 - 0xfa
      10'h112: dout  = 8'b11111010; //  274 : 250 - 0xfa
      10'h113: dout  = 8'b11101001; //  275 : 233 - 0xe9
      10'h114: dout  = 8'b11111010; //  276 : 250 - 0xfa
      10'h115: dout  = 8'b11101010; //  277 : 234 - 0xea
      10'h116: dout  = 8'b11111010; //  278 : 250 - 0xfa
      10'h117: dout  = 8'b11111010; //  279 : 250 - 0xfa
      10'h118: dout  = 8'b11101001; //  280 : 233 - 0xe9
      10'h119: dout  = 8'b11111010; //  281 : 250 - 0xfa
      10'h11A: dout  = 8'b11111010; //  282 : 250 - 0xfa
      10'h11B: dout  = 8'b11101010; //  283 : 234 - 0xea
      10'h11C: dout  = 8'b11111010; //  284 : 250 - 0xfa
      10'h11D: dout  = 8'b11111010; //  285 : 250 - 0xfa
      10'h11E: dout  = 8'b11101001; //  286 : 233 - 0xe9
      10'h11F: dout  = 8'b11111010; //  287 : 250 - 0xfa
      10'h120: dout  = 8'b11111010; //  288 : 250 - 0xfa -- line 0x9
      10'h121: dout  = 8'b11111100; //  289 : 252 - 0xfc
      10'h122: dout  = 8'b11111111; //  290 : 255 - 0xff
      10'h123: dout  = 8'b11111111; //  291 : 255 - 0xff
      10'h124: dout  = 8'b11111111; //  292 : 255 - 0xff
      10'h125: dout  = 8'b11111111; //  293 : 255 - 0xff
      10'h126: dout  = 8'b11101100; //  294 : 236 - 0xec
      10'h127: dout  = 8'b11111010; //  295 : 250 - 0xfa
      10'h128: dout  = 8'b11101001; //  296 : 233 - 0xe9
      10'h129: dout  = 8'b11111010; //  297 : 250 - 0xfa
      10'h12A: dout  = 8'b11101010; //  298 : 234 - 0xea
      10'h12B: dout  = 8'b11111100; //  299 : 252 - 0xfc
      10'h12C: dout  = 8'b11111111; //  300 : 255 - 0xff
      10'h12D: dout  = 8'b11111111; //  301 : 255 - 0xff
      10'h12E: dout  = 8'b11111111; //  302 : 255 - 0xff
      10'h12F: dout  = 8'b11111111; //  303 : 255 - 0xff
      10'h130: dout  = 8'b11101100; //  304 : 236 - 0xec
      10'h131: dout  = 8'b11111010; //  305 : 250 - 0xfa
      10'h132: dout  = 8'b11111010; //  306 : 250 - 0xfa
      10'h133: dout  = 8'b11111010; //  307 : 250 - 0xfa
      10'h134: dout  = 8'b11111010; //  308 : 250 - 0xfa
      10'h135: dout  = 8'b11111010; //  309 : 250 - 0xfa
      10'h136: dout  = 8'b11111010; //  310 : 250 - 0xfa
      10'h137: dout  = 8'b11111010; //  311 : 250 - 0xfa
      10'h138: dout  = 8'b11111010; //  312 : 250 - 0xfa
      10'h139: dout  = 8'b11111010; //  313 : 250 - 0xfa
      10'h13A: dout  = 8'b11111010; //  314 : 250 - 0xfa
      10'h13B: dout  = 8'b11111010; //  315 : 250 - 0xfa
      10'h13C: dout  = 8'b11111010; //  316 : 250 - 0xfa
      10'h13D: dout  = 8'b11111010; //  317 : 250 - 0xfa
      10'h13E: dout  = 8'b11111010; //  318 : 250 - 0xfa
      10'h13F: dout  = 8'b11111010; //  319 : 250 - 0xfa
      10'h140: dout  = 8'b11111010; //  320 : 250 - 0xfa -- line 0xa
      10'h141: dout  = 8'b11111100; //  321 : 252 - 0xfc
      10'h142: dout  = 8'b11111111; //  322 : 255 - 0xff
      10'h143: dout  = 8'b11111110; //  323 : 254 - 0xfe
      10'h144: dout  = 8'b11111110; //  324 : 254 - 0xfe
      10'h145: dout  = 8'b11111111; //  325 : 255 - 0xff
      10'h146: dout  = 8'b11101100; //  326 : 236 - 0xec
      10'h147: dout  = 8'b11111010; //  327 : 250 - 0xfa
      10'h148: dout  = 8'b11111010; //  328 : 250 - 0xfa
      10'h149: dout  = 8'b11111010; //  329 : 250 - 0xfa
      10'h14A: dout  = 8'b11111010; //  330 : 250 - 0xfa
      10'h14B: dout  = 8'b11111100; //  331 : 252 - 0xfc
      10'h14C: dout  = 8'b11111111; //  332 : 255 - 0xff
      10'h14D: dout  = 8'b11111110; //  333 : 254 - 0xfe
      10'h14E: dout  = 8'b11111110; //  334 : 254 - 0xfe
      10'h14F: dout  = 8'b11111111; //  335 : 255 - 0xff
      10'h150: dout  = 8'b11101100; //  336 : 236 - 0xec
      10'h151: dout  = 8'b11101001; //  337 : 233 - 0xe9
      10'h152: dout  = 8'b11111010; //  338 : 250 - 0xfa
      10'h153: dout  = 8'b11111010; //  339 : 250 - 0xfa
      10'h154: dout  = 8'b11111010; //  340 : 250 - 0xfa
      10'h155: dout  = 8'b11111010; //  341 : 250 - 0xfa
      10'h156: dout  = 8'b11111010; //  342 : 250 - 0xfa
      10'h157: dout  = 8'b11111001; //  343 : 249 - 0xf9
      10'h158: dout  = 8'b11111001; //  344 : 249 - 0xf9
      10'h159: dout  = 8'b11111001; //  345 : 249 - 0xf9
      10'h15A: dout  = 8'b11111010; //  346 : 250 - 0xfa
      10'h15B: dout  = 8'b11111010; //  347 : 250 - 0xfa
      10'h15C: dout  = 8'b11111010; //  348 : 250 - 0xfa
      10'h15D: dout  = 8'b11111010; //  349 : 250 - 0xfa
      10'h15E: dout  = 8'b11111010; //  350 : 250 - 0xfa
      10'h15F: dout  = 8'b11111010; //  351 : 250 - 0xfa
      10'h160: dout  = 8'b11111010; //  352 : 250 - 0xfa -- line 0xb
      10'h161: dout  = 8'b11111100; //  353 : 252 - 0xfc
      10'h162: dout  = 8'b11111111; //  354 : 255 - 0xff
      10'h163: dout  = 8'b11111111; //  355 : 255 - 0xff
      10'h164: dout  = 8'b11111111; //  356 : 255 - 0xff
      10'h165: dout  = 8'b11111111; //  357 : 255 - 0xff
      10'h166: dout  = 8'b11101100; //  358 : 236 - 0xec
      10'h167: dout  = 8'b11111010; //  359 : 250 - 0xfa
      10'h168: dout  = 8'b11101010; //  360 : 234 - 0xea
      10'h169: dout  = 8'b11111010; //  361 : 250 - 0xfa
      10'h16A: dout  = 8'b11111010; //  362 : 250 - 0xfa
      10'h16B: dout  = 8'b11111100; //  363 : 252 - 0xfc
      10'h16C: dout  = 8'b11111111; //  364 : 255 - 0xff
      10'h16D: dout  = 8'b11111111; //  365 : 255 - 0xff
      10'h16E: dout  = 8'b11111111; //  366 : 255 - 0xff
      10'h16F: dout  = 8'b11111111; //  367 : 255 - 0xff
      10'h170: dout  = 8'b11110101; //  368 : 245 - 0xf5
      10'h171: dout  = 8'b11111011; //  369 : 251 - 0xfb
      10'h172: dout  = 8'b11101000; //  370 : 232 - 0xe8
      10'h173: dout  = 8'b11111010; //  371 : 250 - 0xfa
      10'h174: dout  = 8'b11111001; //  372 : 249 - 0xf9
      10'h175: dout  = 8'b11101001; //  373 : 233 - 0xe9
      10'h176: dout  = 8'b11111010; //  374 : 250 - 0xfa
      10'h177: dout  = 8'b11111001; //  375 : 249 - 0xf9
      10'h178: dout  = 8'b11111010; //  376 : 250 - 0xfa
      10'h179: dout  = 8'b11111010; //  377 : 250 - 0xfa
      10'h17A: dout  = 8'b11111010; //  378 : 250 - 0xfa
      10'h17B: dout  = 8'b11101001; //  379 : 233 - 0xe9
      10'h17C: dout  = 8'b11111010; //  380 : 250 - 0xfa
      10'h17D: dout  = 8'b11101010; //  381 : 234 - 0xea
      10'h17E: dout  = 8'b11111010; //  382 : 250 - 0xfa
      10'h17F: dout  = 8'b11101001; //  383 : 233 - 0xe9
      10'h180: dout  = 8'b11101001; //  384 : 233 - 0xe9 -- line 0xc
      10'h181: dout  = 8'b11111100; //  385 : 252 - 0xfc
      10'h182: dout  = 8'b11111111; //  386 : 255 - 0xff
      10'h183: dout  = 8'b11111110; //  387 : 254 - 0xfe
      10'h184: dout  = 8'b11111110; //  388 : 254 - 0xfe
      10'h185: dout  = 8'b11111111; //  389 : 255 - 0xff
      10'h186: dout  = 8'b11101100; //  390 : 236 - 0xec
      10'h187: dout  = 8'b11101010; //  391 : 234 - 0xea
      10'h188: dout  = 8'b11111010; //  392 : 250 - 0xfa
      10'h189: dout  = 8'b11101010; //  393 : 234 - 0xea
      10'h18A: dout  = 8'b11111010; //  394 : 250 - 0xfa
      10'h18B: dout  = 8'b11111100; //  395 : 252 - 0xfc
      10'h18C: dout  = 8'b11111111; //  396 : 255 - 0xff
      10'h18D: dout  = 8'b11111110; //  397 : 254 - 0xfe
      10'h18E: dout  = 8'b11111110; //  398 : 254 - 0xfe
      10'h18F: dout  = 8'b11111111; //  399 : 255 - 0xff
      10'h190: dout  = 8'b11111111; //  400 : 255 - 0xff
      10'h191: dout  = 8'b11111111; //  401 : 255 - 0xff
      10'h192: dout  = 8'b11101100; //  402 : 236 - 0xec
      10'h193: dout  = 8'b11111010; //  403 : 250 - 0xfa
      10'h194: dout  = 8'b11111010; //  404 : 250 - 0xfa
      10'h195: dout  = 8'b11111010; //  405 : 250 - 0xfa
      10'h196: dout  = 8'b11111010; //  406 : 250 - 0xfa
      10'h197: dout  = 8'b11111010; //  407 : 250 - 0xfa
      10'h198: dout  = 8'b11111010; //  408 : 250 - 0xfa
      10'h199: dout  = 8'b11101010; //  409 : 234 - 0xea
      10'h19A: dout  = 8'b11111010; //  410 : 250 - 0xfa
      10'h19B: dout  = 8'b11111010; //  411 : 250 - 0xfa
      10'h19C: dout  = 8'b11111010; //  412 : 250 - 0xfa
      10'h19D: dout  = 8'b11111010; //  413 : 250 - 0xfa
      10'h19E: dout  = 8'b11111010; //  414 : 250 - 0xfa
      10'h19F: dout  = 8'b11111010; //  415 : 250 - 0xfa
      10'h1A0: dout  = 8'b11111010; //  416 : 250 - 0xfa -- line 0xd
      10'h1A1: dout  = 8'b11111100; //  417 : 252 - 0xfc
      10'h1A2: dout  = 8'b11111111; //  418 : 255 - 0xff
      10'h1A3: dout  = 8'b11111111; //  419 : 255 - 0xff
      10'h1A4: dout  = 8'b11111111; //  420 : 255 - 0xff
      10'h1A5: dout  = 8'b11111111; //  421 : 255 - 0xff
      10'h1A6: dout  = 8'b11101100; //  422 : 236 - 0xec
      10'h1A7: dout  = 8'b11111010; //  423 : 250 - 0xfa
      10'h1A8: dout  = 8'b11111010; //  424 : 250 - 0xfa
      10'h1A9: dout  = 8'b11111010; //  425 : 250 - 0xfa
      10'h1AA: dout  = 8'b11111010; //  426 : 250 - 0xfa
      10'h1AB: dout  = 8'b11111100; //  427 : 252 - 0xfc
      10'h1AC: dout  = 8'b11111111; //  428 : 255 - 0xff
      10'h1AD: dout  = 8'b11111111; //  429 : 255 - 0xff
      10'h1AE: dout  = 8'b11111111; //  430 : 255 - 0xff
      10'h1AF: dout  = 8'b11111111; //  431 : 255 - 0xff
      10'h1B0: dout  = 8'b11111111; //  432 : 255 - 0xff
      10'h1B1: dout  = 8'b11111111; //  433 : 255 - 0xff
      10'h1B2: dout  = 8'b11110101; //  434 : 245 - 0xf5
      10'h1B3: dout  = 8'b11111011; //  435 : 251 - 0xfb
      10'h1B4: dout  = 8'b11111011; //  436 : 251 - 0xfb
      10'h1B5: dout  = 8'b11111011; //  437 : 251 - 0xfb
      10'h1B6: dout  = 8'b11111011; //  438 : 251 - 0xfb
      10'h1B7: dout  = 8'b11111011; //  439 : 251 - 0xfb
      10'h1B8: dout  = 8'b11111011; //  440 : 251 - 0xfb
      10'h1B9: dout  = 8'b11111011; //  441 : 251 - 0xfb
      10'h1BA: dout  = 8'b11111011; //  442 : 251 - 0xfb
      10'h1BB: dout  = 8'b11111011; //  443 : 251 - 0xfb
      10'h1BC: dout  = 8'b11111011; //  444 : 251 - 0xfb
      10'h1BD: dout  = 8'b11111011; //  445 : 251 - 0xfb
      10'h1BE: dout  = 8'b11101000; //  446 : 232 - 0xe8
      10'h1BF: dout  = 8'b11101001; //  447 : 233 - 0xe9
      10'h1C0: dout  = 8'b11111010; //  448 : 250 - 0xfa -- line 0xe
      10'h1C1: dout  = 8'b11111100; //  449 : 252 - 0xfc
      10'h1C2: dout  = 8'b11111111; //  450 : 255 - 0xff
      10'h1C3: dout  = 8'b11111110; //  451 : 254 - 0xfe
      10'h1C4: dout  = 8'b11111110; //  452 : 254 - 0xfe
      10'h1C5: dout  = 8'b11111111; //  453 : 255 - 0xff
      10'h1C6: dout  = 8'b11101100; //  454 : 236 - 0xec
      10'h1C7: dout  = 8'b11111010; //  455 : 250 - 0xfa
      10'h1C8: dout  = 8'b11111010; //  456 : 250 - 0xfa
      10'h1C9: dout  = 8'b11111001; //  457 : 249 - 0xf9
      10'h1CA: dout  = 8'b11111010; //  458 : 250 - 0xfa
      10'h1CB: dout  = 8'b11111100; //  459 : 252 - 0xfc
      10'h1CC: dout  = 8'b11111111; //  460 : 255 - 0xff
      10'h1CD: dout  = 8'b11111111; //  461 : 255 - 0xff
      10'h1CE: dout  = 8'b11111111; //  462 : 255 - 0xff
      10'h1CF: dout  = 8'b11111110; //  463 : 254 - 0xfe
      10'h1D0: dout  = 8'b11111111; //  464 : 255 - 0xff
      10'h1D1: dout  = 8'b11111111; //  465 : 255 - 0xff
      10'h1D2: dout  = 8'b11111111; //  466 : 255 - 0xff
      10'h1D3: dout  = 8'b11111111; //  467 : 255 - 0xff
      10'h1D4: dout  = 8'b11111111; //  468 : 255 - 0xff
      10'h1D5: dout  = 8'b11111111; //  469 : 255 - 0xff
      10'h1D6: dout  = 8'b11111111; //  470 : 255 - 0xff
      10'h1D7: dout  = 8'b11101111; //  471 : 239 - 0xef
      10'h1D8: dout  = 8'b11111111; //  472 : 255 - 0xff
      10'h1D9: dout  = 8'b11111111; //  473 : 255 - 0xff
      10'h1DA: dout  = 8'b11111111; //  474 : 255 - 0xff
      10'h1DB: dout  = 8'b11111111; //  475 : 255 - 0xff
      10'h1DC: dout  = 8'b11111111; //  476 : 255 - 0xff
      10'h1DD: dout  = 8'b11111111; //  477 : 255 - 0xff
      10'h1DE: dout  = 8'b11101100; //  478 : 236 - 0xec
      10'h1DF: dout  = 8'b11111010; //  479 : 250 - 0xfa
      10'h1E0: dout  = 8'b11101010; //  480 : 234 - 0xea -- line 0xf
      10'h1E1: dout  = 8'b11111100; //  481 : 252 - 0xfc
      10'h1E2: dout  = 8'b11111111; //  482 : 255 - 0xff
      10'h1E3: dout  = 8'b11111111; //  483 : 255 - 0xff
      10'h1E4: dout  = 8'b11111111; //  484 : 255 - 0xff
      10'h1E5: dout  = 8'b11111111; //  485 : 255 - 0xff
      10'h1E6: dout  = 8'b11101100; //  486 : 236 - 0xec
      10'h1E7: dout  = 8'b11111010; //  487 : 250 - 0xfa
      10'h1E8: dout  = 8'b11111010; //  488 : 250 - 0xfa
      10'h1E9: dout  = 8'b11111010; //  489 : 250 - 0xfa
      10'h1EA: dout  = 8'b11111010; //  490 : 250 - 0xfa
      10'h1EB: dout  = 8'b11111100; //  491 : 252 - 0xfc
      10'h1EC: dout  = 8'b11111111; //  492 : 255 - 0xff
      10'h1ED: dout  = 8'b11111111; //  493 : 255 - 0xff
      10'h1EE: dout  = 8'b11111111; //  494 : 255 - 0xff
      10'h1EF: dout  = 8'b11111111; //  495 : 255 - 0xff
      10'h1F0: dout  = 8'b11111111; //  496 : 255 - 0xff
      10'h1F1: dout  = 8'b11111101; //  497 : 253 - 0xfd
      10'h1F2: dout  = 8'b11111111; //  498 : 255 - 0xff
      10'h1F3: dout  = 8'b11111101; //  499 : 253 - 0xfd
      10'h1F4: dout  = 8'b11111111; //  500 : 255 - 0xff
      10'h1F5: dout  = 8'b11111101; //  501 : 253 - 0xfd
      10'h1F6: dout  = 8'b11111111; //  502 : 255 - 0xff
      10'h1F7: dout  = 8'b11101111; //  503 : 239 - 0xef
      10'h1F8: dout  = 8'b11111111; //  504 : 255 - 0xff
      10'h1F9: dout  = 8'b11111101; //  505 : 253 - 0xfd
      10'h1FA: dout  = 8'b11111111; //  506 : 255 - 0xff
      10'h1FB: dout  = 8'b11111111; //  507 : 255 - 0xff
      10'h1FC: dout  = 8'b11111111; //  508 : 255 - 0xff
      10'h1FD: dout  = 8'b11111111; //  509 : 255 - 0xff
      10'h1FE: dout  = 8'b11101100; //  510 : 236 - 0xec
      10'h1FF: dout  = 8'b11111010; //  511 : 250 - 0xfa
      10'h200: dout  = 8'b11111010; //  512 : 250 - 0xfa -- line 0x10
      10'h201: dout  = 8'b11111100; //  513 : 252 - 0xfc
      10'h202: dout  = 8'b11111111; //  514 : 255 - 0xff
      10'h203: dout  = 8'b11111110; //  515 : 254 - 0xfe
      10'h204: dout  = 8'b11111110; //  516 : 254 - 0xfe
      10'h205: dout  = 8'b11111111; //  517 : 255 - 0xff
      10'h206: dout  = 8'b11101100; //  518 : 236 - 0xec
      10'h207: dout  = 8'b11101001; //  519 : 233 - 0xe9
      10'h208: dout  = 8'b11111010; //  520 : 250 - 0xfa
      10'h209: dout  = 8'b11111010; //  521 : 250 - 0xfa
      10'h20A: dout  = 8'b11111010; //  522 : 250 - 0xfa
      10'h20B: dout  = 8'b11110111; //  523 : 247 - 0xf7
      10'h20C: dout  = 8'b11101011; //  524 : 235 - 0xeb
      10'h20D: dout  = 8'b11100110; //  525 : 230 - 0xe6
      10'h20E: dout  = 8'b11111111; //  526 : 255 - 0xff
      10'h20F: dout  = 8'b11111111; //  527 : 255 - 0xff
      10'h210: dout  = 8'b11111111; //  528 : 255 - 0xff
      10'h211: dout  = 8'b11111101; //  529 : 253 - 0xfd
      10'h212: dout  = 8'b11111111; //  530 : 255 - 0xff
      10'h213: dout  = 8'b11111101; //  531 : 253 - 0xfd
      10'h214: dout  = 8'b11111111; //  532 : 255 - 0xff
      10'h215: dout  = 8'b11111101; //  533 : 253 - 0xfd
      10'h216: dout  = 8'b11111111; //  534 : 255 - 0xff
      10'h217: dout  = 8'b11101111; //  535 : 239 - 0xef
      10'h218: dout  = 8'b11111111; //  536 : 255 - 0xff
      10'h219: dout  = 8'b11111101; //  537 : 253 - 0xfd
      10'h21A: dout  = 8'b11111111; //  538 : 255 - 0xff
      10'h21B: dout  = 8'b11111111; //  539 : 255 - 0xff
      10'h21C: dout  = 8'b11111111; //  540 : 255 - 0xff
      10'h21D: dout  = 8'b11111111; //  541 : 255 - 0xff
      10'h21E: dout  = 8'b11101100; //  542 : 236 - 0xec
      10'h21F: dout  = 8'b11101010; //  543 : 234 - 0xea
      10'h220: dout  = 8'b11111010; //  544 : 250 - 0xfa -- line 0x11
      10'h221: dout  = 8'b11111100; //  545 : 252 - 0xfc
      10'h222: dout  = 8'b11111111; //  546 : 255 - 0xff
      10'h223: dout  = 8'b11111111; //  547 : 255 - 0xff
      10'h224: dout  = 8'b11111111; //  548 : 255 - 0xff
      10'h225: dout  = 8'b11111111; //  549 : 255 - 0xff
      10'h226: dout  = 8'b11101100; //  550 : 236 - 0xec
      10'h227: dout  = 8'b11111010; //  551 : 250 - 0xfa
      10'h228: dout  = 8'b11111010; //  552 : 250 - 0xfa
      10'h229: dout  = 8'b11111010; //  553 : 250 - 0xfa
      10'h22A: dout  = 8'b11101010; //  554 : 234 - 0xea
      10'h22B: dout  = 8'b11111010; //  555 : 250 - 0xfa
      10'h22C: dout  = 8'b11111010; //  556 : 250 - 0xfa
      10'h22D: dout  = 8'b11111100; //  557 : 252 - 0xfc
      10'h22E: dout  = 8'b11111111; //  558 : 255 - 0xff
      10'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      10'h230: dout  = 8'b11111111; //  560 : 255 - 0xff
      10'h231: dout  = 8'b11111111; //  561 : 255 - 0xff
      10'h232: dout  = 8'b11111111; //  562 : 255 - 0xff
      10'h233: dout  = 8'b11111111; //  563 : 255 - 0xff
      10'h234: dout  = 8'b11111111; //  564 : 255 - 0xff
      10'h235: dout  = 8'b11111111; //  565 : 255 - 0xff
      10'h236: dout  = 8'b11111111; //  566 : 255 - 0xff
      10'h237: dout  = 8'b11101111; //  567 : 239 - 0xef
      10'h238: dout  = 8'b11111111; //  568 : 255 - 0xff
      10'h239: dout  = 8'b11111111; //  569 : 255 - 0xff
      10'h23A: dout  = 8'b11111111; //  570 : 255 - 0xff
      10'h23B: dout  = 8'b11111110; //  571 : 254 - 0xfe
      10'h23C: dout  = 8'b11111110; //  572 : 254 - 0xfe
      10'h23D: dout  = 8'b11111111; //  573 : 255 - 0xff
      10'h23E: dout  = 8'b11101100; //  574 : 236 - 0xec
      10'h23F: dout  = 8'b11111010; //  575 : 250 - 0xfa
      10'h240: dout  = 8'b11111010; //  576 : 250 - 0xfa -- line 0x12
      10'h241: dout  = 8'b11111100; //  577 : 252 - 0xfc
      10'h242: dout  = 8'b11111111; //  578 : 255 - 0xff
      10'h243: dout  = 8'b11111110; //  579 : 254 - 0xfe
      10'h244: dout  = 8'b11111110; //  580 : 254 - 0xfe
      10'h245: dout  = 8'b11111111; //  581 : 255 - 0xff
      10'h246: dout  = 8'b11101100; //  582 : 236 - 0xec
      10'h247: dout  = 8'b11111001; //  583 : 249 - 0xf9
      10'h248: dout  = 8'b11111010; //  584 : 250 - 0xfa
      10'h249: dout  = 8'b11111010; //  585 : 250 - 0xfa
      10'h24A: dout  = 8'b11111010; //  586 : 250 - 0xfa
      10'h24B: dout  = 8'b11111010; //  587 : 250 - 0xfa
      10'h24C: dout  = 8'b11101010; //  588 : 234 - 0xea
      10'h24D: dout  = 8'b11110111; //  589 : 247 - 0xf7
      10'h24E: dout  = 8'b11101011; //  590 : 235 - 0xeb
      10'h24F: dout  = 8'b11101011; //  591 : 235 - 0xeb
      10'h250: dout  = 8'b11101011; //  592 : 235 - 0xeb
      10'h251: dout  = 8'b11101011; //  593 : 235 - 0xeb
      10'h252: dout  = 8'b11101011; //  594 : 235 - 0xeb
      10'h253: dout  = 8'b11101011; //  595 : 235 - 0xeb
      10'h254: dout  = 8'b11101011; //  596 : 235 - 0xeb
      10'h255: dout  = 8'b11101011; //  597 : 235 - 0xeb
      10'h256: dout  = 8'b11101011; //  598 : 235 - 0xeb
      10'h257: dout  = 8'b11101011; //  599 : 235 - 0xeb
      10'h258: dout  = 8'b11101011; //  600 : 235 - 0xeb
      10'h259: dout  = 8'b11100110; //  601 : 230 - 0xe6
      10'h25A: dout  = 8'b11111111; //  602 : 255 - 0xff
      10'h25B: dout  = 8'b11111111; //  603 : 255 - 0xff
      10'h25C: dout  = 8'b11111111; //  604 : 255 - 0xff
      10'h25D: dout  = 8'b11111111; //  605 : 255 - 0xff
      10'h25E: dout  = 8'b11101100; //  606 : 236 - 0xec
      10'h25F: dout  = 8'b11111010; //  607 : 250 - 0xfa
      10'h260: dout  = 8'b11111001; //  608 : 249 - 0xf9 -- line 0x13
      10'h261: dout  = 8'b11111100; //  609 : 252 - 0xfc
      10'h262: dout  = 8'b11111111; //  610 : 255 - 0xff
      10'h263: dout  = 8'b11111111; //  611 : 255 - 0xff
      10'h264: dout  = 8'b11111111; //  612 : 255 - 0xff
      10'h265: dout  = 8'b11111111; //  613 : 255 - 0xff
      10'h266: dout  = 8'b11110101; //  614 : 245 - 0xf5
      10'h267: dout  = 8'b11111011; //  615 : 251 - 0xfb
      10'h268: dout  = 8'b11111011; //  616 : 251 - 0xfb
      10'h269: dout  = 8'b11111011; //  617 : 251 - 0xfb
      10'h26A: dout  = 8'b11111011; //  618 : 251 - 0xfb
      10'h26B: dout  = 8'b11111011; //  619 : 251 - 0xfb
      10'h26C: dout  = 8'b11111011; //  620 : 251 - 0xfb
      10'h26D: dout  = 8'b11111011; //  621 : 251 - 0xfb
      10'h26E: dout  = 8'b11111011; //  622 : 251 - 0xfb
      10'h26F: dout  = 8'b11111011; //  623 : 251 - 0xfb
      10'h270: dout  = 8'b11111011; //  624 : 251 - 0xfb
      10'h271: dout  = 8'b11111011; //  625 : 251 - 0xfb
      10'h272: dout  = 8'b11101000; //  626 : 232 - 0xe8
      10'h273: dout  = 8'b11111010; //  627 : 250 - 0xfa
      10'h274: dout  = 8'b11111010; //  628 : 250 - 0xfa
      10'h275: dout  = 8'b11101010; //  629 : 234 - 0xea
      10'h276: dout  = 8'b11111010; //  630 : 250 - 0xfa
      10'h277: dout  = 8'b11111010; //  631 : 250 - 0xfa
      10'h278: dout  = 8'b11101001; //  632 : 233 - 0xe9
      10'h279: dout  = 8'b11111100; //  633 : 252 - 0xfc
      10'h27A: dout  = 8'b11111111; //  634 : 255 - 0xff
      10'h27B: dout  = 8'b11111110; //  635 : 254 - 0xfe
      10'h27C: dout  = 8'b11111110; //  636 : 254 - 0xfe
      10'h27D: dout  = 8'b11111111; //  637 : 255 - 0xff
      10'h27E: dout  = 8'b11101100; //  638 : 236 - 0xec
      10'h27F: dout  = 8'b11111010; //  639 : 250 - 0xfa
      10'h280: dout  = 8'b11111010; //  640 : 250 - 0xfa -- line 0x14
      10'h281: dout  = 8'b11111100; //  641 : 252 - 0xfc
      10'h282: dout  = 8'b11111111; //  642 : 255 - 0xff
      10'h283: dout  = 8'b11111110; //  643 : 254 - 0xfe
      10'h284: dout  = 8'b11111110; //  644 : 254 - 0xfe
      10'h285: dout  = 8'b11111111; //  645 : 255 - 0xff
      10'h286: dout  = 8'b11111111; //  646 : 255 - 0xff
      10'h287: dout  = 8'b11111101; //  647 : 253 - 0xfd
      10'h288: dout  = 8'b11111111; //  648 : 255 - 0xff
      10'h289: dout  = 8'b11111101; //  649 : 253 - 0xfd
      10'h28A: dout  = 8'b11111111; //  650 : 255 - 0xff
      10'h28B: dout  = 8'b11111101; //  651 : 253 - 0xfd
      10'h28C: dout  = 8'b11111111; //  652 : 255 - 0xff
      10'h28D: dout  = 8'b11111101; //  653 : 253 - 0xfd
      10'h28E: dout  = 8'b11111111; //  654 : 255 - 0xff
      10'h28F: dout  = 8'b11111101; //  655 : 253 - 0xfd
      10'h290: dout  = 8'b11111111; //  656 : 255 - 0xff
      10'h291: dout  = 8'b11111111; //  657 : 255 - 0xff
      10'h292: dout  = 8'b11101100; //  658 : 236 - 0xec
      10'h293: dout  = 8'b11101001; //  659 : 233 - 0xe9
      10'h294: dout  = 8'b11111010; //  660 : 250 - 0xfa
      10'h295: dout  = 8'b11111010; //  661 : 250 - 0xfa
      10'h296: dout  = 8'b11101010; //  662 : 234 - 0xea
      10'h297: dout  = 8'b11111010; //  663 : 250 - 0xfa
      10'h298: dout  = 8'b11111010; //  664 : 250 - 0xfa
      10'h299: dout  = 8'b11111100; //  665 : 252 - 0xfc
      10'h29A: dout  = 8'b11111111; //  666 : 255 - 0xff
      10'h29B: dout  = 8'b11111111; //  667 : 255 - 0xff
      10'h29C: dout  = 8'b11111111; //  668 : 255 - 0xff
      10'h29D: dout  = 8'b11111111; //  669 : 255 - 0xff
      10'h29E: dout  = 8'b11101100; //  670 : 236 - 0xec
      10'h29F: dout  = 8'b11101010; //  671 : 234 - 0xea
      10'h2A0: dout  = 8'b11111010; //  672 : 250 - 0xfa -- line 0x15
      10'h2A1: dout  = 8'b11111100; //  673 : 252 - 0xfc
      10'h2A2: dout  = 8'b11111111; //  674 : 255 - 0xff
      10'h2A3: dout  = 8'b11111111; //  675 : 255 - 0xff
      10'h2A4: dout  = 8'b11111111; //  676 : 255 - 0xff
      10'h2A5: dout  = 8'b11111111; //  677 : 255 - 0xff
      10'h2A6: dout  = 8'b11111111; //  678 : 255 - 0xff
      10'h2A7: dout  = 8'b11111101; //  679 : 253 - 0xfd
      10'h2A8: dout  = 8'b11111111; //  680 : 255 - 0xff
      10'h2A9: dout  = 8'b11111101; //  681 : 253 - 0xfd
      10'h2AA: dout  = 8'b11111111; //  682 : 255 - 0xff
      10'h2AB: dout  = 8'b11111101; //  683 : 253 - 0xfd
      10'h2AC: dout  = 8'b11111111; //  684 : 255 - 0xff
      10'h2AD: dout  = 8'b11111101; //  685 : 253 - 0xfd
      10'h2AE: dout  = 8'b11111111; //  686 : 255 - 0xff
      10'h2AF: dout  = 8'b11111101; //  687 : 253 - 0xfd
      10'h2B0: dout  = 8'b11111111; //  688 : 255 - 0xff
      10'h2B1: dout  = 8'b11111111; //  689 : 255 - 0xff
      10'h2B2: dout  = 8'b11101100; //  690 : 236 - 0xec
      10'h2B3: dout  = 8'b11100111; //  691 : 231 - 0xe7
      10'h2B4: dout  = 8'b11111011; //  692 : 251 - 0xfb
      10'h2B5: dout  = 8'b11111011; //  693 : 251 - 0xfb
      10'h2B6: dout  = 8'b11111011; //  694 : 251 - 0xfb
      10'h2B7: dout  = 8'b11111011; //  695 : 251 - 0xfb
      10'h2B8: dout  = 8'b11111011; //  696 : 251 - 0xfb
      10'h2B9: dout  = 8'b11110110; //  697 : 246 - 0xf6
      10'h2BA: dout  = 8'b11111111; //  698 : 255 - 0xff
      10'h2BB: dout  = 8'b11111110; //  699 : 254 - 0xfe
      10'h2BC: dout  = 8'b11111110; //  700 : 254 - 0xfe
      10'h2BD: dout  = 8'b11111111; //  701 : 255 - 0xff
      10'h2BE: dout  = 8'b11101100; //  702 : 236 - 0xec
      10'h2BF: dout  = 8'b11111010; //  703 : 250 - 0xfa
      10'h2C0: dout  = 8'b11111010; //  704 : 250 - 0xfa -- line 0x16
      10'h2C1: dout  = 8'b11111100; //  705 : 252 - 0xfc
      10'h2C2: dout  = 8'b11111111; //  706 : 255 - 0xff
      10'h2C3: dout  = 8'b11111110; //  707 : 254 - 0xfe
      10'h2C4: dout  = 8'b11111110; //  708 : 254 - 0xfe
      10'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      10'h2C6: dout  = 8'b11100101; //  710 : 229 - 0xe5
      10'h2C7: dout  = 8'b11101011; //  711 : 235 - 0xeb
      10'h2C8: dout  = 8'b11101011; //  712 : 235 - 0xeb
      10'h2C9: dout  = 8'b11101011; //  713 : 235 - 0xeb
      10'h2CA: dout  = 8'b11101011; //  714 : 235 - 0xeb
      10'h2CB: dout  = 8'b11101011; //  715 : 235 - 0xeb
      10'h2CC: dout  = 8'b11101011; //  716 : 235 - 0xeb
      10'h2CD: dout  = 8'b11101011; //  717 : 235 - 0xeb
      10'h2CE: dout  = 8'b11101011; //  718 : 235 - 0xeb
      10'h2CF: dout  = 8'b11100110; //  719 : 230 - 0xe6
      10'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff
      10'h2D1: dout  = 8'b11111111; //  721 : 255 - 0xff
      10'h2D2: dout  = 8'b11101100; //  722 : 236 - 0xec
      10'h2D3: dout  = 8'b11111100; //  723 : 252 - 0xfc
      10'h2D4: dout  = 8'b11111111; //  724 : 255 - 0xff
      10'h2D5: dout  = 8'b11111111; //  725 : 255 - 0xff
      10'h2D6: dout  = 8'b11111111; //  726 : 255 - 0xff
      10'h2D7: dout  = 8'b11111111; //  727 : 255 - 0xff
      10'h2D8: dout  = 8'b11111111; //  728 : 255 - 0xff
      10'h2D9: dout  = 8'b11111111; //  729 : 255 - 0xff
      10'h2DA: dout  = 8'b11111111; //  730 : 255 - 0xff
      10'h2DB: dout  = 8'b11111111; //  731 : 255 - 0xff
      10'h2DC: dout  = 8'b11111111; //  732 : 255 - 0xff
      10'h2DD: dout  = 8'b11111111; //  733 : 255 - 0xff
      10'h2DE: dout  = 8'b11101100; //  734 : 236 - 0xec
      10'h2DF: dout  = 8'b11111010; //  735 : 250 - 0xfa
      10'h2E0: dout  = 8'b11111010; //  736 : 250 - 0xfa -- line 0x17
      10'h2E1: dout  = 8'b11111100; //  737 : 252 - 0xfc
      10'h2E2: dout  = 8'b11111111; //  738 : 255 - 0xff
      10'h2E3: dout  = 8'b11111111; //  739 : 255 - 0xff
      10'h2E4: dout  = 8'b11111111; //  740 : 255 - 0xff
      10'h2E5: dout  = 8'b11111111; //  741 : 255 - 0xff
      10'h2E6: dout  = 8'b11110101; //  742 : 245 - 0xf5
      10'h2E7: dout  = 8'b11111011; //  743 : 251 - 0xfb
      10'h2E8: dout  = 8'b11111011; //  744 : 251 - 0xfb
      10'h2E9: dout  = 8'b11111011; //  745 : 251 - 0xfb
      10'h2EA: dout  = 8'b11111011; //  746 : 251 - 0xfb
      10'h2EB: dout  = 8'b11111011; //  747 : 251 - 0xfb
      10'h2EC: dout  = 8'b11111011; //  748 : 251 - 0xfb
      10'h2ED: dout  = 8'b11111011; //  749 : 251 - 0xfb
      10'h2EE: dout  = 8'b11111011; //  750 : 251 - 0xfb
      10'h2EF: dout  = 8'b11110110; //  751 : 246 - 0xf6
      10'h2F0: dout  = 8'b11111111; //  752 : 255 - 0xff
      10'h2F1: dout  = 8'b11111111; //  753 : 255 - 0xff
      10'h2F2: dout  = 8'b11110101; //  754 : 245 - 0xf5
      10'h2F3: dout  = 8'b11110110; //  755 : 246 - 0xf6
      10'h2F4: dout  = 8'b11111111; //  756 : 255 - 0xff
      10'h2F5: dout  = 8'b11111111; //  757 : 255 - 0xff
      10'h2F6: dout  = 8'b11111111; //  758 : 255 - 0xff
      10'h2F7: dout  = 8'b11111111; //  759 : 255 - 0xff
      10'h2F8: dout  = 8'b11111111; //  760 : 255 - 0xff
      10'h2F9: dout  = 8'b11111111; //  761 : 255 - 0xff
      10'h2FA: dout  = 8'b11111111; //  762 : 255 - 0xff
      10'h2FB: dout  = 8'b11111110; //  763 : 254 - 0xfe
      10'h2FC: dout  = 8'b11111110; //  764 : 254 - 0xfe
      10'h2FD: dout  = 8'b11111111; //  765 : 255 - 0xff
      10'h2FE: dout  = 8'b11101100; //  766 : 236 - 0xec
      10'h2FF: dout  = 8'b11111010; //  767 : 250 - 0xfa
      10'h300: dout  = 8'b11111010; //  768 : 250 - 0xfa -- line 0x18
      10'h301: dout  = 8'b11111100; //  769 : 252 - 0xfc
      10'h302: dout  = 8'b11111111; //  770 : 255 - 0xff
      10'h303: dout  = 8'b11111110; //  771 : 254 - 0xfe
      10'h304: dout  = 8'b11111110; //  772 : 254 - 0xfe
      10'h305: dout  = 8'b11111111; //  773 : 255 - 0xff
      10'h306: dout  = 8'b11111111; //  774 : 255 - 0xff
      10'h307: dout  = 8'b11111111; //  775 : 255 - 0xff
      10'h308: dout  = 8'b11111111; //  776 : 255 - 0xff
      10'h309: dout  = 8'b11111111; //  777 : 255 - 0xff
      10'h30A: dout  = 8'b11111111; //  778 : 255 - 0xff
      10'h30B: dout  = 8'b11111111; //  779 : 255 - 0xff
      10'h30C: dout  = 8'b11111111; //  780 : 255 - 0xff
      10'h30D: dout  = 8'b11111111; //  781 : 255 - 0xff
      10'h30E: dout  = 8'b11111111; //  782 : 255 - 0xff
      10'h30F: dout  = 8'b11111111; //  783 : 255 - 0xff
      10'h310: dout  = 8'b11111111; //  784 : 255 - 0xff
      10'h311: dout  = 8'b11111111; //  785 : 255 - 0xff
      10'h312: dout  = 8'b11111111; //  786 : 255 - 0xff
      10'h313: dout  = 8'b11111111; //  787 : 255 - 0xff
      10'h314: dout  = 8'b11111111; //  788 : 255 - 0xff
      10'h315: dout  = 8'b11111101; //  789 : 253 - 0xfd
      10'h316: dout  = 8'b11111111; //  790 : 255 - 0xff
      10'h317: dout  = 8'b11111101; //  791 : 253 - 0xfd
      10'h318: dout  = 8'b11111111; //  792 : 255 - 0xff
      10'h319: dout  = 8'b11111101; //  793 : 253 - 0xfd
      10'h31A: dout  = 8'b11111111; //  794 : 255 - 0xff
      10'h31B: dout  = 8'b11111111; //  795 : 255 - 0xff
      10'h31C: dout  = 8'b11111111; //  796 : 255 - 0xff
      10'h31D: dout  = 8'b11111111; //  797 : 255 - 0xff
      10'h31E: dout  = 8'b11101100; //  798 : 236 - 0xec
      10'h31F: dout  = 8'b11101001; //  799 : 233 - 0xe9
      10'h320: dout  = 8'b11101010; //  800 : 234 - 0xea -- line 0x19
      10'h321: dout  = 8'b11111100; //  801 : 252 - 0xfc
      10'h322: dout  = 8'b11111111; //  802 : 255 - 0xff
      10'h323: dout  = 8'b11111111; //  803 : 255 - 0xff
      10'h324: dout  = 8'b11111111; //  804 : 255 - 0xff
      10'h325: dout  = 8'b11111111; //  805 : 255 - 0xff
      10'h326: dout  = 8'b11111111; //  806 : 255 - 0xff
      10'h327: dout  = 8'b11111101; //  807 : 253 - 0xfd
      10'h328: dout  = 8'b11111111; //  808 : 255 - 0xff
      10'h329: dout  = 8'b11111101; //  809 : 253 - 0xfd
      10'h32A: dout  = 8'b11111111; //  810 : 255 - 0xff
      10'h32B: dout  = 8'b11111101; //  811 : 253 - 0xfd
      10'h32C: dout  = 8'b11111111; //  812 : 255 - 0xff
      10'h32D: dout  = 8'b11111101; //  813 : 253 - 0xfd
      10'h32E: dout  = 8'b11111111; //  814 : 255 - 0xff
      10'h32F: dout  = 8'b11111101; //  815 : 253 - 0xfd
      10'h330: dout  = 8'b11111111; //  816 : 255 - 0xff
      10'h331: dout  = 8'b11111101; //  817 : 253 - 0xfd
      10'h332: dout  = 8'b11111111; //  818 : 255 - 0xff
      10'h333: dout  = 8'b11111101; //  819 : 253 - 0xfd
      10'h334: dout  = 8'b11111111; //  820 : 255 - 0xff
      10'h335: dout  = 8'b11111101; //  821 : 253 - 0xfd
      10'h336: dout  = 8'b11111111; //  822 : 255 - 0xff
      10'h337: dout  = 8'b11111101; //  823 : 253 - 0xfd
      10'h338: dout  = 8'b11111111; //  824 : 255 - 0xff
      10'h339: dout  = 8'b11111101; //  825 : 253 - 0xfd
      10'h33A: dout  = 8'b11111111; //  826 : 255 - 0xff
      10'h33B: dout  = 8'b11111111; //  827 : 255 - 0xff
      10'h33C: dout  = 8'b11111111; //  828 : 255 - 0xff
      10'h33D: dout  = 8'b11111111; //  829 : 255 - 0xff
      10'h33E: dout  = 8'b11101100; //  830 : 236 - 0xec
      10'h33F: dout  = 8'b11111010; //  831 : 250 - 0xfa
      10'h340: dout  = 8'b11111010; //  832 : 250 - 0xfa -- line 0x1a
      10'h341: dout  = 8'b11110111; //  833 : 247 - 0xf7
      10'h342: dout  = 8'b11101011; //  834 : 235 - 0xeb
      10'h343: dout  = 8'b11100110; //  835 : 230 - 0xe6
      10'h344: dout  = 8'b11111111; //  836 : 255 - 0xff
      10'h345: dout  = 8'b11111111; //  837 : 255 - 0xff
      10'h346: dout  = 8'b11111111; //  838 : 255 - 0xff
      10'h347: dout  = 8'b11111101; //  839 : 253 - 0xfd
      10'h348: dout  = 8'b11111111; //  840 : 255 - 0xff
      10'h349: dout  = 8'b11111101; //  841 : 253 - 0xfd
      10'h34A: dout  = 8'b11111111; //  842 : 255 - 0xff
      10'h34B: dout  = 8'b11111101; //  843 : 253 - 0xfd
      10'h34C: dout  = 8'b11111111; //  844 : 255 - 0xff
      10'h34D: dout  = 8'b11111101; //  845 : 253 - 0xfd
      10'h34E: dout  = 8'b11111111; //  846 : 255 - 0xff
      10'h34F: dout  = 8'b11111101; //  847 : 253 - 0xfd
      10'h350: dout  = 8'b11111111; //  848 : 255 - 0xff
      10'h351: dout  = 8'b11111101; //  849 : 253 - 0xfd
      10'h352: dout  = 8'b11111111; //  850 : 255 - 0xff
      10'h353: dout  = 8'b11111101; //  851 : 253 - 0xfd
      10'h354: dout  = 8'b11111111; //  852 : 255 - 0xff
      10'h355: dout  = 8'b11111111; //  853 : 255 - 0xff
      10'h356: dout  = 8'b11111111; //  854 : 255 - 0xff
      10'h357: dout  = 8'b11111111; //  855 : 255 - 0xff
      10'h358: dout  = 8'b11111111; //  856 : 255 - 0xff
      10'h359: dout  = 8'b11111111; //  857 : 255 - 0xff
      10'h35A: dout  = 8'b11111111; //  858 : 255 - 0xff
      10'h35B: dout  = 8'b11111111; //  859 : 255 - 0xff
      10'h35C: dout  = 8'b11100101; //  860 : 229 - 0xe5
      10'h35D: dout  = 8'b11101011; //  861 : 235 - 0xeb
      10'h35E: dout  = 8'b11111000; //  862 : 248 - 0xf8
      10'h35F: dout  = 8'b11111010; //  863 : 250 - 0xfa
      10'h360: dout  = 8'b11111010; //  864 : 250 - 0xfa -- line 0x1b
      10'h361: dout  = 8'b11111010; //  865 : 250 - 0xfa
      10'h362: dout  = 8'b11111010; //  866 : 250 - 0xfa
      10'h363: dout  = 8'b11111100; //  867 : 252 - 0xfc
      10'h364: dout  = 8'b11111111; //  868 : 255 - 0xff
      10'h365: dout  = 8'b11111111; //  869 : 255 - 0xff
      10'h366: dout  = 8'b11111111; //  870 : 255 - 0xff
      10'h367: dout  = 8'b11111111; //  871 : 255 - 0xff
      10'h368: dout  = 8'b11111111; //  872 : 255 - 0xff
      10'h369: dout  = 8'b11111111; //  873 : 255 - 0xff
      10'h36A: dout  = 8'b11111111; //  874 : 255 - 0xff
      10'h36B: dout  = 8'b11111111; //  875 : 255 - 0xff
      10'h36C: dout  = 8'b11111111; //  876 : 255 - 0xff
      10'h36D: dout  = 8'b11111111; //  877 : 255 - 0xff
      10'h36E: dout  = 8'b11111111; //  878 : 255 - 0xff
      10'h36F: dout  = 8'b11111111; //  879 : 255 - 0xff
      10'h370: dout  = 8'b11111111; //  880 : 255 - 0xff
      10'h371: dout  = 8'b11111111; //  881 : 255 - 0xff
      10'h372: dout  = 8'b11111111; //  882 : 255 - 0xff
      10'h373: dout  = 8'b11111111; //  883 : 255 - 0xff
      10'h374: dout  = 8'b11111111; //  884 : 255 - 0xff
      10'h375: dout  = 8'b11111111; //  885 : 255 - 0xff
      10'h376: dout  = 8'b11111111; //  886 : 255 - 0xff
      10'h377: dout  = 8'b11111111; //  887 : 255 - 0xff
      10'h378: dout  = 8'b11111111; //  888 : 255 - 0xff
      10'h379: dout  = 8'b11111111; //  889 : 255 - 0xff
      10'h37A: dout  = 8'b11111111; //  890 : 255 - 0xff
      10'h37B: dout  = 8'b11111111; //  891 : 255 - 0xff
      10'h37C: dout  = 8'b11101100; //  892 : 236 - 0xec
      10'h37D: dout  = 8'b11111010; //  893 : 250 - 0xfa
      10'h37E: dout  = 8'b11111010; //  894 : 250 - 0xfa
      10'h37F: dout  = 8'b11111001; //  895 : 249 - 0xf9
      10'h380: dout  = 8'b11111010; //  896 : 250 - 0xfa -- line 0x1c
      10'h381: dout  = 8'b11111010; //  897 : 250 - 0xfa
      10'h382: dout  = 8'b11111010; //  898 : 250 - 0xfa
      10'h383: dout  = 8'b11110111; //  899 : 247 - 0xf7
      10'h384: dout  = 8'b11101011; //  900 : 235 - 0xeb
      10'h385: dout  = 8'b11101011; //  901 : 235 - 0xeb
      10'h386: dout  = 8'b11101011; //  902 : 235 - 0xeb
      10'h387: dout  = 8'b11101011; //  903 : 235 - 0xeb
      10'h388: dout  = 8'b11101011; //  904 : 235 - 0xeb
      10'h389: dout  = 8'b11101011; //  905 : 235 - 0xeb
      10'h38A: dout  = 8'b11101011; //  906 : 235 - 0xeb
      10'h38B: dout  = 8'b11101011; //  907 : 235 - 0xeb
      10'h38C: dout  = 8'b11101011; //  908 : 235 - 0xeb
      10'h38D: dout  = 8'b11101011; //  909 : 235 - 0xeb
      10'h38E: dout  = 8'b11101011; //  910 : 235 - 0xeb
      10'h38F: dout  = 8'b11101011; //  911 : 235 - 0xeb
      10'h390: dout  = 8'b11101011; //  912 : 235 - 0xeb
      10'h391: dout  = 8'b11101011; //  913 : 235 - 0xeb
      10'h392: dout  = 8'b11101011; //  914 : 235 - 0xeb
      10'h393: dout  = 8'b11101011; //  915 : 235 - 0xeb
      10'h394: dout  = 8'b11101011; //  916 : 235 - 0xeb
      10'h395: dout  = 8'b11101011; //  917 : 235 - 0xeb
      10'h396: dout  = 8'b11101011; //  918 : 235 - 0xeb
      10'h397: dout  = 8'b11101011; //  919 : 235 - 0xeb
      10'h398: dout  = 8'b11101011; //  920 : 235 - 0xeb
      10'h399: dout  = 8'b11101011; //  921 : 235 - 0xeb
      10'h39A: dout  = 8'b11101011; //  922 : 235 - 0xeb
      10'h39B: dout  = 8'b11101011; //  923 : 235 - 0xeb
      10'h39C: dout  = 8'b11111000; //  924 : 248 - 0xf8
      10'h39D: dout  = 8'b11111010; //  925 : 250 - 0xfa
      10'h39E: dout  = 8'b11111010; //  926 : 250 - 0xfa
      10'h39F: dout  = 8'b11111010; //  927 : 250 - 0xfa
      10'h3A0: dout  = 8'b11111010; //  928 : 250 - 0xfa -- line 0x1d
      10'h3A1: dout  = 8'b11111001; //  929 : 249 - 0xf9
      10'h3A2: dout  = 8'b11111010; //  930 : 250 - 0xfa
      10'h3A3: dout  = 8'b11111010; //  931 : 250 - 0xfa
      10'h3A4: dout  = 8'b11111010; //  932 : 250 - 0xfa
      10'h3A5: dout  = 8'b11111010; //  933 : 250 - 0xfa
      10'h3A6: dout  = 8'b11111010; //  934 : 250 - 0xfa
      10'h3A7: dout  = 8'b11111010; //  935 : 250 - 0xfa
      10'h3A8: dout  = 8'b11111010; //  936 : 250 - 0xfa
      10'h3A9: dout  = 8'b11111010; //  937 : 250 - 0xfa
      10'h3AA: dout  = 8'b11111010; //  938 : 250 - 0xfa
      10'h3AB: dout  = 8'b11111010; //  939 : 250 - 0xfa
      10'h3AC: dout  = 8'b11111010; //  940 : 250 - 0xfa
      10'h3AD: dout  = 8'b11111010; //  941 : 250 - 0xfa
      10'h3AE: dout  = 8'b11111010; //  942 : 250 - 0xfa
      10'h3AF: dout  = 8'b11111010; //  943 : 250 - 0xfa
      10'h3B0: dout  = 8'b11111010; //  944 : 250 - 0xfa
      10'h3B1: dout  = 8'b11111010; //  945 : 250 - 0xfa
      10'h3B2: dout  = 8'b11111010; //  946 : 250 - 0xfa
      10'h3B3: dout  = 8'b11111010; //  947 : 250 - 0xfa
      10'h3B4: dout  = 8'b11111010; //  948 : 250 - 0xfa
      10'h3B5: dout  = 8'b11101001; //  949 : 233 - 0xe9
      10'h3B6: dout  = 8'b11111010; //  950 : 250 - 0xfa
      10'h3B7: dout  = 8'b11111010; //  951 : 250 - 0xfa
      10'h3B8: dout  = 8'b11111010; //  952 : 250 - 0xfa
      10'h3B9: dout  = 8'b11111010; //  953 : 250 - 0xfa
      10'h3BA: dout  = 8'b11111010; //  954 : 250 - 0xfa
      10'h3BB: dout  = 8'b11111010; //  955 : 250 - 0xfa
      10'h3BC: dout  = 8'b11101010; //  956 : 234 - 0xea
      10'h3BD: dout  = 8'b11111010; //  957 : 250 - 0xfa
      10'h3BE: dout  = 8'b11111010; //  958 : 250 - 0xfa
      10'h3BF: dout  = 8'b11111010; //  959 : 250 - 0xfa
        //-- Attribute Table 0----
      10'h3C0: dout  = 8'b01010101; //  960 :  85 - 0x55
      10'h3C1: dout  = 8'b00000101; //  961 :   5 - 0x5
      10'h3C2: dout  = 8'b00000101; //  962 :   5 - 0x5
      10'h3C3: dout  = 8'b00000101; //  963 :   5 - 0x5
      10'h3C4: dout  = 8'b01010101; //  964 :  85 - 0x55
      10'h3C5: dout  = 8'b01010101; //  965 :  85 - 0x55
      10'h3C6: dout  = 8'b01010101; //  966 :  85 - 0x55
      10'h3C7: dout  = 8'b01010101; //  967 :  85 - 0x55
      10'h3C8: dout  = 8'b00010001; //  968 :  17 - 0x11
      10'h3C9: dout  = 8'b01000000; //  969 :  64 - 0x40
      10'h3CA: dout  = 8'b01010000; //  970 :  80 - 0x50
      10'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      10'h3CC: dout  = 8'b01010101; //  972 :  85 - 0x55
      10'h3CD: dout  = 8'b01010101; //  973 :  85 - 0x55
      10'h3CE: dout  = 8'b01010101; //  974 :  85 - 0x55
      10'h3CF: dout  = 8'b01010101; //  975 :  85 - 0x55
      10'h3D0: dout  = 8'b00010001; //  976 :  17 - 0x11
      10'h3D1: dout  = 8'b01000100; //  977 :  68 - 0x44
      10'h3D2: dout  = 8'b01010101; //  978 :  85 - 0x55
      10'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      10'h3D4: dout  = 8'b01010101; //  980 :  85 - 0x55
      10'h3D5: dout  = 8'b01010101; //  981 :  85 - 0x55
      10'h3D6: dout  = 8'b01010101; //  982 :  85 - 0x55
      10'h3D7: dout  = 8'b01010101; //  983 :  85 - 0x55
      10'h3D8: dout  = 8'b00010001; //  984 :  17 - 0x11
      10'h3D9: dout  = 8'b01000100; //  985 :  68 - 0x44
      10'h3DA: dout  = 8'b01010101; //  986 :  85 - 0x55
      10'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      10'h3DC: dout  = 8'b00000100; //  988 :   4 - 0x4
      10'h3DD: dout  = 8'b00000101; //  989 :   5 - 0x5
      10'h3DE: dout  = 8'b00000101; //  990 :   5 - 0x5
      10'h3DF: dout  = 8'b01000101; //  991 :  69 - 0x45
      10'h3E0: dout  = 8'b00010001; //  992 :  17 - 0x11
      10'h3E1: dout  = 8'b01000100; //  993 :  68 - 0x44
      10'h3E2: dout  = 8'b01010101; //  994 :  85 - 0x55
      10'h3E3: dout  = 8'b01010001; //  995 :  81 - 0x51
      10'h3E4: dout  = 8'b01010000; //  996 :  80 - 0x50
      10'h3E5: dout  = 8'b01010000; //  997 :  80 - 0x50
      10'h3E6: dout  = 8'b00010000; //  998 :  16 - 0x10
      10'h3E7: dout  = 8'b01000100; //  999 :  68 - 0x44
      10'h3E8: dout  = 8'b00010001; // 1000 :  17 - 0x11
      10'h3E9: dout  = 8'b01000000; // 1001 :  64 - 0x40
      10'h3EA: dout  = 8'b01010000; // 1002 :  80 - 0x50
      10'h3EB: dout  = 8'b01010000; // 1003 :  80 - 0x50
      10'h3EC: dout  = 8'b01000100; // 1004 :  68 - 0x44
      10'h3ED: dout  = 8'b00000101; // 1005 :   5 - 0x5
      10'h3EE: dout  = 8'b00000001; // 1006 :   1 - 0x1
      10'h3EF: dout  = 8'b01000100; // 1007 :  68 - 0x44
      10'h3F0: dout  = 8'b01010001; // 1008 :  81 - 0x51
      10'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      10'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      10'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      10'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      10'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      10'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      10'h3F7: dout  = 8'b01010100; // 1015 :  84 - 0x54
      10'h3F8: dout  = 8'b00000101; // 1016 :   5 - 0x5
      10'h3F9: dout  = 8'b00000101; // 1017 :   5 - 0x5
      10'h3FA: dout  = 8'b00000101; // 1018 :   5 - 0x5
      10'h3FB: dout  = 8'b00000101; // 1019 :   5 - 0x5
      10'h3FC: dout  = 8'b00000101; // 1020 :   5 - 0x5
      10'h3FD: dout  = 8'b00000101; // 1021 :   5 - 0x5
      10'h3FE: dout  = 8'b00000101; // 1022 :   5 - 0x5
      10'h3FF: dout  = 8'b00000101; // 1023 :   5 - 0x5
    endcase
  end

endmodule
