--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_color1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_color1;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_color1 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "01111111", --    1 -  0x1  :  127 - 0x7f
    "01111111", --    2 -  0x2  :  127 - 0x7f
    "01111111", --    3 -  0x3  :  127 - 0x7f
    "01111111", --    4 -  0x4  :  127 - 0x7f
    "01111111", --    5 -  0x5  :  127 - 0x7f
    "01101010", --    6 -  0x6  :  106 - 0x6a
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "01111011", --    9 -  0x9  :  123 - 0x7b
    "01110011", --   10 -  0xa  :  115 - 0x73
    "01111011", --   11 -  0xb  :  123 - 0x7b
    "01110011", --   12 -  0xc  :  115 - 0x73
    "01111011", --   13 -  0xd  :  123 - 0x7b
    "01010011", --   14 -  0xe  :   83 - 0x53
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x2
    "11011110", --   17 - 0x11  :  222 - 0xde
    "10011110", --   18 - 0x12  :  158 - 0x9e
    "11011100", --   19 - 0x13  :  220 - 0xdc
    "10011110", --   20 - 0x14  :  158 - 0x9e
    "11011100", --   21 - 0x15  :  220 - 0xdc
    "10011010", --   22 - 0x16  :  154 - 0x9a
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Sprite 0x3
    "11111110", --   25 - 0x19  :  254 - 0xfe
    "11111100", --   26 - 0x1a  :  252 - 0xfc
    "11111110", --   27 - 0x1b  :  254 - 0xfe
    "11111100", --   28 - 0x1c  :  252 - 0xfc
    "11111110", --   29 - 0x1d  :  254 - 0xfe
    "01010100", --   30 - 0x1e  :   84 - 0x54
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x4
    "01111111", --   33 - 0x21  :  127 - 0x7f
    "01011111", --   34 - 0x22  :   95 - 0x5f
    "01111001", --   35 - 0x23  :  121 - 0x79
    "01111001", --   36 - 0x24  :  121 - 0x79
    "01001001", --   37 - 0x25  :   73 - 0x49
    "01001111", --   38 - 0x26  :   79 - 0x4f
    "01001110", --   39 - 0x27  :   78 - 0x4e
    "01111000", --   40 - 0x28  :  120 - 0x78 -- Sprite 0x5
    "01110000", --   41 - 0x29  :  112 - 0x70
    "01100000", --   42 - 0x2a  :   96 - 0x60
    "01100000", --   43 - 0x2b  :   96 - 0x60
    "01110001", --   44 - 0x2c  :  113 - 0x71
    "01011111", --   45 - 0x2d  :   95 - 0x5f
    "01111111", --   46 - 0x2e  :  127 - 0x7f
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x6
    "11111110", --   49 - 0x31  :  254 - 0xfe
    "11111010", --   50 - 0x32  :  250 - 0xfa
    "10011110", --   51 - 0x33  :  158 - 0x9e
    "10011110", --   52 - 0x34  :  158 - 0x9e
    "10010010", --   53 - 0x35  :  146 - 0x92
    "11110010", --   54 - 0x36  :  242 - 0xf2
    "01110010", --   55 - 0x37  :  114 - 0x72
    "00011110", --   56 - 0x38  :   30 - 0x1e -- Sprite 0x7
    "00001110", --   57 - 0x39  :   14 - 0xe
    "00000110", --   58 - 0x3a  :    6 - 0x6
    "00000110", --   59 - 0x3b  :    6 - 0x6
    "10001110", --   60 - 0x3c  :  142 - 0x8e
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111110", --   62 - 0x3e  :  254 - 0xfe
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "01111111", --   65 - 0x41  :  127 - 0x7f
    "01011111", --   66 - 0x42  :   95 - 0x5f
    "01111111", --   67 - 0x43  :  127 - 0x7f
    "01111111", --   68 - 0x44  :  127 - 0x7f
    "01111111", --   69 - 0x45  :  127 - 0x7f
    "01111111", --   70 - 0x46  :  127 - 0x7f
    "01111111", --   71 - 0x47  :  127 - 0x7f
    "01111111", --   72 - 0x48  :  127 - 0x7f -- Sprite 0x9
    "01111111", --   73 - 0x49  :  127 - 0x7f
    "01111111", --   74 - 0x4a  :  127 - 0x7f
    "01111111", --   75 - 0x4b  :  127 - 0x7f
    "01111111", --   76 - 0x4c  :  127 - 0x7f
    "01011111", --   77 - 0x4d  :   95 - 0x5f
    "01111111", --   78 - 0x4e  :  127 - 0x7f
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0xa
    "11111110", --   81 - 0x51  :  254 - 0xfe
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111110", --   83 - 0x53  :  254 - 0xfe
    "11111110", --   84 - 0x54  :  254 - 0xfe
    "11111110", --   85 - 0x55  :  254 - 0xfe
    "11111110", --   86 - 0x56  :  254 - 0xfe
    "11111110", --   87 - 0x57  :  254 - 0xfe
    "11111110", --   88 - 0x58  :  254 - 0xfe -- Sprite 0xb
    "11111110", --   89 - 0x59  :  254 - 0xfe
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111110", --   91 - 0x5b  :  254 - 0xfe
    "11111110", --   92 - 0x5c  :  254 - 0xfe
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111110", --   94 - 0x5e  :  254 - 0xfe
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0xc
    "00111111", --   97 - 0x61  :   63 - 0x3f
    "01011111", --   98 - 0x62  :   95 - 0x5f
    "01101111", --   99 - 0x63  :  111 - 0x6f
    "01110000", --  100 - 0x64  :  112 - 0x70
    "01110111", --  101 - 0x65  :  119 - 0x77
    "01110111", --  102 - 0x66  :  119 - 0x77
    "01110111", --  103 - 0x67  :  119 - 0x77
    "01110111", --  104 - 0x68  :  119 - 0x77 -- Sprite 0xd
    "01110111", --  105 - 0x69  :  119 - 0x77
    "01110111", --  106 - 0x6a  :  119 - 0x77
    "01110000", --  107 - 0x6b  :  112 - 0x70
    "01101111", --  108 - 0x6c  :  111 - 0x6f
    "01011111", --  109 - 0x6d  :   95 - 0x5f
    "00010101", --  110 - 0x6e  :   21 - 0x15
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0xe
    "11111100", --  113 - 0x71  :  252 - 0xfc
    "11111000", --  114 - 0x72  :  248 - 0xf8
    "11110110", --  115 - 0x73  :  246 - 0xf6
    "00001100", --  116 - 0x74  :   12 - 0xc
    "11101110", --  117 - 0x75  :  238 - 0xee
    "11101100", --  118 - 0x76  :  236 - 0xec
    "11101110", --  119 - 0x77  :  238 - 0xee
    "11101100", --  120 - 0x78  :  236 - 0xec -- Sprite 0xf
    "11101110", --  121 - 0x79  :  238 - 0xee
    "11101100", --  122 - 0x7a  :  236 - 0xec
    "00001110", --  123 - 0x7b  :   14 - 0xe
    "11110100", --  124 - 0x7c  :  244 - 0xf4
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "01010100", --  126 - 0x7e  :   84 - 0x54
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "01100000", --  128 - 0x80  :   96 - 0x60 -- Sprite 0x10
    "01100000", --  129 - 0x81  :   96 - 0x60
    "01100000", --  130 - 0x82  :   96 - 0x60
    "01101111", --  131 - 0x83  :  111 - 0x6f
    "01101010", --  132 - 0x84  :  106 - 0x6a
    "01100000", --  133 - 0x85  :   96 - 0x60
    "01100000", --  134 - 0x86  :   96 - 0x60
    "01100000", --  135 - 0x87  :   96 - 0x60
    "00000110", --  136 - 0x88  :    6 - 0x6 -- Sprite 0x11
    "00000100", --  137 - 0x89  :    4 - 0x4
    "00000110", --  138 - 0x8a  :    6 - 0x6
    "11110100", --  139 - 0x8b  :  244 - 0xf4
    "10100110", --  140 - 0x8c  :  166 - 0xa6
    "00000100", --  141 - 0x8d  :    4 - 0x4
    "00000110", --  142 - 0x8e  :    6 - 0x6
    "00000100", --  143 - 0x8f  :    4 - 0x4
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x12
    "00001000", --  145 - 0x91  :    8 - 0x8
    "00001000", --  146 - 0x92  :    8 - 0x8
    "00011100", --  147 - 0x93  :   28 - 0x1c
    "00011100", --  148 - 0x94  :   28 - 0x1c
    "00111100", --  149 - 0x95  :   60 - 0x3c
    "00111100", --  150 - 0x96  :   60 - 0x3c
    "00111100", --  151 - 0x97  :   60 - 0x3c
    "00111100", --  152 - 0x98  :   60 - 0x3c -- Sprite 0x13
    "01111110", --  153 - 0x99  :  126 - 0x7e
    "01111110", --  154 - 0x9a  :  126 - 0x7e
    "01111110", --  155 - 0x9b  :  126 - 0x7e
    "01111110", --  156 - 0x9c  :  126 - 0x7e
    "01111110", --  157 - 0x9d  :  126 - 0x7e
    "01111110", --  158 - 0x9e  :  126 - 0x7e
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000101", --  162 - 0xa2  :    5 - 0x5
    "00000011", --  163 - 0xa3  :    3 - 0x3
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000010", --  166 - 0xa6  :    2 - 0x2
    "00001111", --  167 - 0xa7  :   15 - 0xf
    "00011100", --  168 - 0xa8  :   28 - 0x1c -- Sprite 0x15
    "00111010", --  169 - 0xa9  :   58 - 0x3a
    "00111100", --  170 - 0xaa  :   60 - 0x3c
    "00111111", --  171 - 0xab  :   63 - 0x3f
    "00111000", --  172 - 0xac  :   56 - 0x38
    "00011110", --  173 - 0xad  :   30 - 0x1e
    "00001111", --  174 - 0xae  :   15 - 0xf
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "01000000", --  178 - 0xb2  :   64 - 0x40
    "11000000", --  179 - 0xb3  :  192 - 0xc0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "10000000", --  181 - 0xb5  :  128 - 0x80
    "11000000", --  182 - 0xb6  :  192 - 0xc0
    "01110000", --  183 - 0xb7  :  112 - 0x70
    "00011000", --  184 - 0xb8  :   24 - 0x18 -- Sprite 0x17
    "11111100", --  185 - 0xb9  :  252 - 0xfc
    "00111100", --  186 - 0xba  :   60 - 0x3c
    "01011100", --  187 - 0xbb  :   92 - 0x5c
    "00111100", --  188 - 0xbc  :   60 - 0x3c
    "11111000", --  189 - 0xbd  :  248 - 0xf8
    "11110000", --  190 - 0xbe  :  240 - 0xf0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0x18
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "00111111", --  194 - 0xc2  :   63 - 0x3f
    "01111111", --  195 - 0xc3  :  127 - 0x7f
    "01111111", --  196 - 0xc4  :  127 - 0x7f
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Sprite 0x19
    "11111100", --  201 - 0xc9  :  252 - 0xfc
    "11111100", --  202 - 0xca  :  252 - 0xfc
    "11111110", --  203 - 0xcb  :  254 - 0xfe
    "11111110", --  204 - 0xcc  :  254 - 0xfe
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00111111", --  211 - 0xd3  :   63 - 0x3f
    "00111111", --  212 - 0xd4  :   63 - 0x3f
    "01111111", --  213 - 0xd5  :  127 - 0x7f
    "01111111", --  214 - 0xd6  :  127 - 0x7f
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "11111100", --  219 - 0xdb  :  252 - 0xfc
    "11111100", --  220 - 0xdc  :  252 - 0xfc
    "11111110", --  221 - 0xdd  :  254 - 0xfe
    "11111110", --  222 - 0xde  :  254 - 0xfe
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0x1c
    "01111111", --  225 - 0xe1  :  127 - 0x7f
    "01111111", --  226 - 0xe2  :  127 - 0x7f
    "01111111", --  227 - 0xe3  :  127 - 0x7f
    "01100100", --  228 - 0xe4  :  100 - 0x64
    "01011011", --  229 - 0xe5  :   91 - 0x5b
    "01011001", --  230 - 0xe6  :   89 - 0x59
    "01111111", --  231 - 0xe7  :  127 - 0x7f
    "01111111", --  232 - 0xe8  :  127 - 0x7f -- Sprite 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000001", --  234 - 0xea  :    1 - 0x1
    "00000001", --  235 - 0xeb  :    1 - 0x1
    "00000001", --  236 - 0xec  :    1 - 0x1
    "00000001", --  237 - 0xed  :    1 - 0x1
    "00000001", --  238 - 0xee  :    1 - 0x1
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0x1e
    "11111110", --  241 - 0xf1  :  254 - 0xfe
    "11111110", --  242 - 0xf2  :  254 - 0xfe
    "11111110", --  243 - 0xf3  :  254 - 0xfe
    "10111110", --  244 - 0xf4  :  190 - 0xbe
    "00001010", --  245 - 0xf5  :   10 - 0xa
    "11100010", --  246 - 0xf6  :  226 - 0xe2
    "11111110", --  247 - 0xf7  :  254 - 0xfe
    "11111110", --  248 - 0xf8  :  254 - 0xfe -- Sprite 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "10000000", --  250 - 0xfa  :  128 - 0x80
    "10000000", --  251 - 0xfb  :  128 - 0x80
    "10000000", --  252 - 0xfc  :  128 - 0x80
    "10000000", --  253 - 0xfd  :  128 - 0x80
    "10000000", --  254 - 0xfe  :  128 - 0x80
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00011000", --  274 - 0x112  :   24 - 0x18
    "00010000", --  275 - 0x113  :   16 - 0x10
    "00011010", --  276 - 0x114  :   26 - 0x1a
    "00010001", --  277 - 0x115  :   17 - 0x11
    "00011010", --  278 - 0x116  :   26 - 0x1a
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- Sprite 0x23
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00101000", --  283 - 0x11b  :   40 - 0x28
    "10001100", --  284 - 0x11c  :  140 - 0x8c
    "00101000", --  285 - 0x11d  :   40 - 0x28
    "10101100", --  286 - 0x11e  :  172 - 0xac
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00011100", --  296 - 0x128  :   28 - 0x1c -- Sprite 0x25
    "00111001", --  297 - 0x129  :   57 - 0x39
    "00111111", --  298 - 0x12a  :   63 - 0x3f
    "00111110", --  299 - 0x12b  :   62 - 0x3e
    "00111111", --  300 - 0x12c  :   63 - 0x3f
    "00011110", --  301 - 0x12d  :   30 - 0x1e
    "00001111", --  302 - 0x12e  :   15 - 0xf
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "01000000", --  306 - 0x132  :   64 - 0x40
    "11000000", --  307 - 0x133  :  192 - 0xc0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "10000000", --  309 - 0x135  :  128 - 0x80
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "11110000", --  311 - 0x137  :  240 - 0xf0
    "00111000", --  312 - 0x138  :   56 - 0x38 -- Sprite 0x27
    "10011100", --  313 - 0x139  :  156 - 0x9c
    "10011100", --  314 - 0x13a  :  156 - 0x9c
    "00111100", --  315 - 0x13b  :   60 - 0x3c
    "11111100", --  316 - 0x13c  :  252 - 0xfc
    "01111000", --  317 - 0x13d  :  120 - 0x78
    "11110000", --  318 - 0x13e  :  240 - 0xf0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00111110", --  321 - 0x141  :   62 - 0x3e
    "01011101", --  322 - 0x142  :   93 - 0x5d
    "01101011", --  323 - 0x143  :  107 - 0x6b
    "01110101", --  324 - 0x144  :  117 - 0x75
    "01110001", --  325 - 0x145  :  113 - 0x71
    "01110101", --  326 - 0x146  :  117 - 0x75
    "01110100", --  327 - 0x147  :  116 - 0x74
    "01110000", --  328 - 0x148  :  112 - 0x70 -- Sprite 0x29
    "01110111", --  329 - 0x149  :  119 - 0x77
    "01110111", --  330 - 0x14a  :  119 - 0x77
    "01110000", --  331 - 0x14b  :  112 - 0x70
    "01101111", --  332 - 0x14c  :  111 - 0x6f
    "01011111", --  333 - 0x14d  :   95 - 0x5f
    "00010101", --  334 - 0x14e  :   21 - 0x15
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Sprite 0x2a
    "01111100", --  337 - 0x151  :  124 - 0x7c
    "10111000", --  338 - 0x152  :  184 - 0xb8
    "11010110", --  339 - 0x153  :  214 - 0xd6
    "10101100", --  340 - 0x154  :  172 - 0xac
    "10001110", --  341 - 0x155  :  142 - 0x8e
    "10101100", --  342 - 0x156  :  172 - 0xac
    "00101110", --  343 - 0x157  :   46 - 0x2e
    "00001100", --  344 - 0x158  :   12 - 0xc -- Sprite 0x2b
    "11101110", --  345 - 0x159  :  238 - 0xee
    "11101100", --  346 - 0x15a  :  236 - 0xec
    "00001110", --  347 - 0x15b  :   14 - 0xe
    "11110100", --  348 - 0x15c  :  244 - 0xf4
    "11111010", --  349 - 0x15d  :  250 - 0xfa
    "01010100", --  350 - 0x15e  :   84 - 0x54
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00011110", --  360 - 0x168  :   30 - 0x1e -- Sprite 0x2d
    "00111110", --  361 - 0x169  :   62 - 0x3e
    "00111110", --  362 - 0x16a  :   62 - 0x3e
    "00111110", --  363 - 0x16b  :   62 - 0x3e
    "00111111", --  364 - 0x16c  :   63 - 0x3f
    "00011110", --  365 - 0x16d  :   30 - 0x1e
    "00001111", --  366 - 0x16e  :   15 - 0xf
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "01111000", --  376 - 0x178  :  120 - 0x78 -- Sprite 0x2f
    "01111100", --  377 - 0x179  :  124 - 0x7c
    "01111100", --  378 - 0x17a  :  124 - 0x7c
    "01111100", --  379 - 0x17b  :  124 - 0x7c
    "11111100", --  380 - 0x17c  :  252 - 0xfc
    "01111000", --  381 - 0x17d  :  120 - 0x78
    "11110000", --  382 - 0x17e  :  240 - 0xf0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x30
    "00011000", --  385 - 0x181  :   24 - 0x18
    "00111100", --  386 - 0x182  :   60 - 0x3c
    "01011010", --  387 - 0x183  :   90 - 0x5a
    "00011000", --  388 - 0x184  :   24 - 0x18
    "00011000", --  389 - 0x185  :   24 - 0x18
    "00011000", --  390 - 0x186  :   24 - 0x18
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Sprite 0x31
    "00011000", --  393 - 0x189  :   24 - 0x18
    "00011000", --  394 - 0x18a  :   24 - 0x18
    "00011000", --  395 - 0x18b  :   24 - 0x18
    "01011010", --  396 - 0x18c  :   90 - 0x5a
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00011000", --  398 - 0x18e  :   24 - 0x18
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000001", --  400 - 0x190  :    1 - 0x1 -- Sprite 0x32
    "00000001", --  401 - 0x191  :    1 - 0x1
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000001", --  403 - 0x193  :    1 - 0x1
    "00000001", --  404 - 0x194  :    1 - 0x1
    "00000001", --  405 - 0x195  :    1 - 0x1
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000001", --  407 - 0x197  :    1 - 0x1
    "10000000", --  408 - 0x198  :  128 - 0x80 -- Sprite 0x33
    "00000000", --  409 - 0x199  :    0 - 0x0
    "10000000", --  410 - 0x19a  :  128 - 0x80
    "10000000", --  411 - 0x19b  :  128 - 0x80
    "10000000", --  412 - 0x19c  :  128 - 0x80
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "10000000", --  414 - 0x19e  :  128 - 0x80
    "10000000", --  415 - 0x19f  :  128 - 0x80
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00011000", --  418 - 0x1a2  :   24 - 0x18
    "00111100", --  419 - 0x1a3  :   60 - 0x3c
    "00111110", --  420 - 0x1a4  :   62 - 0x3e
    "01111111", --  421 - 0x1a5  :  127 - 0x7f
    "01111111", --  422 - 0x1a6  :  127 - 0x7f
    "01111111", --  423 - 0x1a7  :  127 - 0x7f
    "00111111", --  424 - 0x1a8  :   63 - 0x3f -- Sprite 0x35
    "00111111", --  425 - 0x1a9  :   63 - 0x3f
    "00011111", --  426 - 0x1aa  :   31 - 0x1f
    "00001111", --  427 - 0x1ab  :   15 - 0xf
    "00000111", --  428 - 0x1ac  :    7 - 0x7
    "00000011", --  429 - 0x1ad  :    3 - 0x3
    "00000001", --  430 - 0x1ae  :    1 - 0x1
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00011000", --  434 - 0x1b2  :   24 - 0x18
    "00111100", --  435 - 0x1b3  :   60 - 0x3c
    "01111100", --  436 - 0x1b4  :  124 - 0x7c
    "11111110", --  437 - 0x1b5  :  254 - 0xfe
    "11111110", --  438 - 0x1b6  :  254 - 0xfe
    "11111110", --  439 - 0x1b7  :  254 - 0xfe
    "11111100", --  440 - 0x1b8  :  252 - 0xfc -- Sprite 0x37
    "11111100", --  441 - 0x1b9  :  252 - 0xfc
    "11111000", --  442 - 0x1ba  :  248 - 0xf8
    "11110000", --  443 - 0x1bb  :  240 - 0xf0
    "11100000", --  444 - 0x1bc  :  224 - 0xe0
    "11000000", --  445 - 0x1bd  :  192 - 0xc0
    "10000000", --  446 - 0x1be  :  128 - 0x80
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000110", --  450 - 0x1c2  :    6 - 0x6
    "00000111", --  451 - 0x1c3  :    7 - 0x7
    "00000111", --  452 - 0x1c4  :    7 - 0x7
    "00000011", --  453 - 0x1c5  :    3 - 0x3
    "00000001", --  454 - 0x1c6  :    1 - 0x1
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "01100000", --  466 - 0x1d2  :   96 - 0x60
    "11100000", --  467 - 0x1d3  :  224 - 0xe0
    "11100000", --  468 - 0x1d4  :  224 - 0xe0
    "11000000", --  469 - 0x1d5  :  192 - 0xc0
    "10000000", --  470 - 0x1d6  :  128 - 0x80
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "00101010", --  473 - 0x1d9  :   42 - 0x2a
    "01000000", --  474 - 0x1da  :   64 - 0x40
    "00000010", --  475 - 0x1db  :    2 - 0x2
    "01000000", --  476 - 0x1dc  :   64 - 0x40
    "00000010", --  477 - 0x1dd  :    2 - 0x2
    "01010100", --  478 - 0x1de  :   84 - 0x54
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "11111111", --  488 - 0x1e8  :  255 - 0xff -- Sprite 0x3d
    "11111111", --  489 - 0x1e9  :  255 - 0xff
    "11111111", --  490 - 0x1ea  :  255 - 0xff
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "11111111", --  492 - 0x1ec  :  255 - 0xff
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "11111111", --  494 - 0x1ee  :  255 - 0xff
    "11111111", --  495 - 0x1ef  :  255 - 0xff
    "11111111", --  496 - 0x1f0  :  255 - 0xff -- Sprite 0x3e
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111111", --  499 - 0x1f3  :  255 - 0xff
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Sprite 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Sprite 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Sprite 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Sprite 0x46
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Sprite 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Sprite 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Sprite 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Sprite 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Sprite 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Sprite 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00111111", --  641 - 0x281  :   63 - 0x3f
    "01111111", --  642 - 0x282  :  127 - 0x7f
    "01111111", --  643 - 0x283  :  127 - 0x7f
    "01111111", --  644 - 0x284  :  127 - 0x7f
    "00111100", --  645 - 0x285  :   60 - 0x3c
    "00000000", --  646 - 0x286  :    0 - 0x0
    "01000000", --  647 - 0x287  :   64 - 0x40
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "11111100", --  649 - 0x289  :  252 - 0xfc
    "11111110", --  650 - 0x28a  :  254 - 0xfe
    "11111110", --  651 - 0x28b  :  254 - 0xfe
    "11111110", --  652 - 0x28c  :  254 - 0xfe
    "00111100", --  653 - 0x28d  :   60 - 0x3c
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000010", --  655 - 0x28f  :    2 - 0x2
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000011", --  658 - 0x292  :    3 - 0x3
    "00000111", --  659 - 0x293  :    7 - 0x7
    "00001111", --  660 - 0x294  :   15 - 0xf
    "00011111", --  661 - 0x295  :   31 - 0x1f
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00110000", --  663 - 0x297  :   48 - 0x30
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "10100000", --  666 - 0x29a  :  160 - 0xa0
    "10110000", --  667 - 0x29b  :  176 - 0xb0
    "10110000", --  668 - 0x29c  :  176 - 0xb0
    "10111000", --  669 - 0x29d  :  184 - 0xb8
    "01111100", --  670 - 0x29e  :  124 - 0x7c
    "01111100", --  671 - 0x29f  :  124 - 0x7c
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x54
    "00100001", --  673 - 0x2a1  :   33 - 0x21
    "01110001", --  674 - 0x2a2  :  113 - 0x71
    "00111010", --  675 - 0x2a3  :   58 - 0x3a
    "01101101", --  676 - 0x2a4  :  109 - 0x6d
    "00111000", --  677 - 0x2a5  :   56 - 0x38
    "00011101", --  678 - 0x2a6  :   29 - 0x1d
    "00101111", --  679 - 0x2a7  :   47 - 0x2f
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00100001", --  681 - 0x2a9  :   33 - 0x21
    "01110001", --  682 - 0x2aa  :  113 - 0x71
    "00111010", --  683 - 0x2ab  :   58 - 0x3a
    "01101101", --  684 - 0x2ac  :  109 - 0x6d
    "10111000", --  685 - 0x2ad  :  184 - 0xb8
    "00011101", --  686 - 0x2ae  :   29 - 0x1d
    "10101111", --  687 - 0x2af  :  175 - 0xaf
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Sprite 0x56
    "00100000", --  689 - 0x2b1  :   32 - 0x20
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "00111010", --  691 - 0x2b3  :   58 - 0x3a
    "01101100", --  692 - 0x2b4  :  108 - 0x6c
    "10111000", --  693 - 0x2b5  :  184 - 0xb8
    "00011100", --  694 - 0x2b6  :   28 - 0x1c
    "10101110", --  695 - 0x2b7  :  174 - 0xae
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Sprite 0x57
    "01111111", --  697 - 0x2b9  :  127 - 0x7f
    "01001100", --  698 - 0x2ba  :   76 - 0x4c
    "00110011", --  699 - 0x2bb  :   51 - 0x33
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x58
    "11111111", --  705 - 0x2c1  :  255 - 0xff
    "11001100", --  706 - 0x2c2  :  204 - 0xcc
    "00110011", --  707 - 0x2c3  :   51 - 0x33
    "11001100", --  708 - 0x2c4  :  204 - 0xcc
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Sprite 0x59
    "11111110", --  713 - 0x2c9  :  254 - 0xfe
    "11001100", --  714 - 0x2ca  :  204 - 0xcc
    "00110000", --  715 - 0x2cb  :   48 - 0x30
    "11000000", --  716 - 0x2cc  :  192 - 0xc0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000001", --  732 - 0x2dc  :    1 - 0x1
    "00000001", --  733 - 0x2dd  :    1 - 0x1
    "00000011", --  734 - 0x2de  :    3 - 0x3
    "00000011", --  735 - 0x2df  :    3 - 0x3
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000001", --  738 - 0x2e2  :    1 - 0x1
    "01111110", --  739 - 0x2e3  :  126 - 0x7e
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11111111", --  743 - 0x2e7  :  255 - 0xff
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Sprite 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "01111111", --  748 - 0x2ec  :  127 - 0x7f
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111111", --  751 - 0x2ef  :  255 - 0xff
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "10000000", --  754 - 0x2f2  :  128 - 0x80
    "01111110", --  755 - 0x2f3  :  126 - 0x7e
    "10111111", --  756 - 0x2f4  :  191 - 0xbf
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Sprite 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "10000000", --  764 - 0x2fc  :  128 - 0x80
    "10000000", --  765 - 0x2fd  :  128 - 0x80
    "11000000", --  766 - 0x2fe  :  192 - 0xc0
    "11000000", --  767 - 0x2ff  :  192 - 0xc0
    "01111111", --  768 - 0x300  :  127 - 0x7f -- Sprite 0x60
    "01111111", --  769 - 0x301  :  127 - 0x7f
    "01111101", --  770 - 0x302  :  125 - 0x7d
    "01111111", --  771 - 0x303  :  127 - 0x7f
    "00111111", --  772 - 0x304  :   63 - 0x3f
    "01111111", --  773 - 0x305  :  127 - 0x7f
    "01111111", --  774 - 0x306  :  127 - 0x7f
    "01110111", --  775 - 0x307  :  119 - 0x77
    "11111110", --  776 - 0x308  :  254 - 0xfe -- Sprite 0x61
    "11111110", --  777 - 0x309  :  254 - 0xfe
    "11111100", --  778 - 0x30a  :  252 - 0xfc
    "11111110", --  779 - 0x30b  :  254 - 0xfe
    "10111110", --  780 - 0x30c  :  190 - 0xbe
    "11111110", --  781 - 0x30d  :  254 - 0xfe
    "11111110", --  782 - 0x30e  :  254 - 0xfe
    "11110110", --  783 - 0x30f  :  246 - 0xf6
    "00000111", --  784 - 0x310  :    7 - 0x7 -- Sprite 0x62
    "00011111", --  785 - 0x311  :   31 - 0x1f
    "00111111", --  786 - 0x312  :   63 - 0x3f
    "00111111", --  787 - 0x313  :   63 - 0x3f
    "00111111", --  788 - 0x314  :   63 - 0x3f
    "00011111", --  789 - 0x315  :   31 - 0x1f
    "00001111", --  790 - 0x316  :   15 - 0xf
    "00000000", --  791 - 0x317  :    0 - 0x0
    "01111110", --  792 - 0x318  :  126 - 0x7e -- Sprite 0x63
    "01111100", --  793 - 0x319  :  124 - 0x7c
    "00111110", --  794 - 0x31a  :   62 - 0x3e
    "10111100", --  795 - 0x31b  :  188 - 0xbc
    "10111110", --  796 - 0x31c  :  190 - 0xbe
    "10011100", --  797 - 0x31d  :  156 - 0x9c
    "11011000", --  798 - 0x31e  :  216 - 0xd8
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "01000110", --  800 - 0x320  :   70 - 0x46 -- Sprite 0x64
    "01101011", --  801 - 0x321  :  107 - 0x6b
    "01110001", --  802 - 0x322  :  113 - 0x71
    "00111010", --  803 - 0x323  :   58 - 0x3a
    "01101101", --  804 - 0x324  :  109 - 0x6d
    "00111000", --  805 - 0x325  :   56 - 0x38
    "00011101", --  806 - 0x326  :   29 - 0x1d
    "00101111", --  807 - 0x327  :   47 - 0x2f
    "01000110", --  808 - 0x328  :   70 - 0x46 -- Sprite 0x65
    "11101011", --  809 - 0x329  :  235 - 0xeb
    "01110001", --  810 - 0x32a  :  113 - 0x71
    "00111010", --  811 - 0x32b  :   58 - 0x3a
    "01101101", --  812 - 0x32c  :  109 - 0x6d
    "10111000", --  813 - 0x32d  :  184 - 0xb8
    "00011101", --  814 - 0x32e  :   29 - 0x1d
    "10101111", --  815 - 0x32f  :  175 - 0xaf
    "01000110", --  816 - 0x330  :   70 - 0x46 -- Sprite 0x66
    "11101010", --  817 - 0x331  :  234 - 0xea
    "01110000", --  818 - 0x332  :  112 - 0x70
    "00111010", --  819 - 0x333  :   58 - 0x3a
    "01101100", --  820 - 0x334  :  108 - 0x6c
    "10111000", --  821 - 0x335  :  184 - 0xb8
    "00011100", --  822 - 0x336  :   28 - 0x1c
    "10101110", --  823 - 0x337  :  174 - 0xae
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Sprite 0x67
    "01111111", --  825 - 0x339  :  127 - 0x7f
    "01111111", --  826 - 0x33a  :  127 - 0x7f
    "00110011", --  827 - 0x33b  :   51 - 0x33
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "11111111", --  833 - 0x341  :  255 - 0xff
    "11111111", --  834 - 0x342  :  255 - 0xff
    "11111111", --  835 - 0x343  :  255 - 0xff
    "11001100", --  836 - 0x344  :  204 - 0xcc
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "11111110", --  841 - 0x349  :  254 - 0xfe
    "11111110", --  842 - 0x34a  :  254 - 0xfe
    "11110000", --  843 - 0x34b  :  240 - 0xf0
    "11000000", --  844 - 0x34c  :  192 - 0xc0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00111101", --  856 - 0x358  :   61 - 0x3d -- Sprite 0x6b
    "01111111", --  857 - 0x359  :  127 - 0x7f
    "01111111", --  858 - 0x35a  :  127 - 0x7f
    "01111111", --  859 - 0x35b  :  127 - 0x7f
    "00111111", --  860 - 0x35c  :   63 - 0x3f
    "00001111", --  861 - 0x35d  :   15 - 0xf
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111111", --  864 - 0x360  :  255 - 0xff -- Sprite 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111110", --  870 - 0x366  :  254 - 0xfe
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "10111000", --  888 - 0x378  :  184 - 0xb8 -- Sprite 0x6f
    "11111100", --  889 - 0x379  :  252 - 0xfc
    "11111110", --  890 - 0x37a  :  254 - 0xfe
    "11111110", --  891 - 0x37b  :  254 - 0xfe
    "11111100", --  892 - 0x37c  :  252 - 0xfc
    "11110000", --  893 - 0x37d  :  240 - 0xf0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x70
    "00111111", --  897 - 0x381  :   63 - 0x3f
    "01111111", --  898 - 0x382  :  127 - 0x7f
    "01111111", --  899 - 0x383  :  127 - 0x7f
    "00011100", --  900 - 0x384  :   28 - 0x1c
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Sprite 0x71
    "11111111", --  905 - 0x389  :  255 - 0xff
    "11111111", --  906 - 0x38a  :  255 - 0xff
    "11111111", --  907 - 0x38b  :  255 - 0xff
    "11111111", --  908 - 0x38c  :  255 - 0xff
    "00111100", --  909 - 0x38d  :   60 - 0x3c
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x72
    "11111100", --  913 - 0x391  :  252 - 0xfc
    "11111110", --  914 - 0x392  :  254 - 0xfe
    "11111110", --  915 - 0x393  :  254 - 0xfe
    "00111000", --  916 - 0x394  :   56 - 0x38
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111101", --  922 - 0x39a  :  253 - 0xfd
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "10111111", --  924 - 0x39c  :  191 - 0xbf
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11110111", --  927 - 0x39f  :  247 - 0xf7
    "01000110", --  928 - 0x3a0  :   70 - 0x46 -- Sprite 0x74
    "01101011", --  929 - 0x3a1  :  107 - 0x6b
    "01110001", --  930 - 0x3a2  :  113 - 0x71
    "00111010", --  931 - 0x3a3  :   58 - 0x3a
    "01101101", --  932 - 0x3a4  :  109 - 0x6d
    "00111000", --  933 - 0x3a5  :   56 - 0x38
    "00011101", --  934 - 0x3a6  :   29 - 0x1d
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "01000110", --  936 - 0x3a8  :   70 - 0x46 -- Sprite 0x75
    "11101011", --  937 - 0x3a9  :  235 - 0xeb
    "01110001", --  938 - 0x3aa  :  113 - 0x71
    "00111010", --  939 - 0x3ab  :   58 - 0x3a
    "01101101", --  940 - 0x3ac  :  109 - 0x6d
    "10111000", --  941 - 0x3ad  :  184 - 0xb8
    "00011101", --  942 - 0x3ae  :   29 - 0x1d
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "01000110", --  944 - 0x3b0  :   70 - 0x46 -- Sprite 0x76
    "11101010", --  945 - 0x3b1  :  234 - 0xea
    "01110000", --  946 - 0x3b2  :  112 - 0x70
    "00111010", --  947 - 0x3b3  :   58 - 0x3a
    "01101100", --  948 - 0x3b4  :  108 - 0x6c
    "10111000", --  949 - 0x3b5  :  184 - 0xb8
    "00011100", --  950 - 0x3b6  :   28 - 0x1c
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "10000001", --  952 - 0x3b8  :  129 - 0x81 -- Sprite 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111101", --  954 - 0x3ba  :  253 - 0xfd
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "10111111", --  956 - 0x3bc  :  191 - 0xbf
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11110111", --  959 - 0x3bf  :  247 - 0xf7
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00100010", --  993 - 0x3e1  :   34 - 0x22
    "01110111", --  994 - 0x3e2  :  119 - 0x77
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111011", --  996 - 0x3e4  :  251 - 0xfb
    "11110101", --  997 - 0x3e5  :  245 - 0xf5
    "11101111", --  998 - 0x3e6  :  239 - 0xef
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "01110011", -- 1001 - 0x3e9  :  115 - 0x73
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111011", -- 1004 - 0x3ec  :  251 - 0xfb
    "11111101", -- 1005 - 0x3ed  :  253 - 0xfd
    "11101111", -- 1006 - 0x3ee  :  239 - 0xef
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "11011111", -- 1008 - 0x3f0  :  223 - 0xdf -- Sprite 0x7e
    "10101111", -- 1009 - 0x3f1  :  175 - 0xaf
    "01111111", -- 1010 - 0x3f2  :  127 - 0x7f
    "11111111", -- 1011 - 0x3f3  :  255 - 0xff
    "11111011", -- 1012 - 0x3f4  :  251 - 0xfb
    "11110101", -- 1013 - 0x3f5  :  245 - 0xf5
    "11101111", -- 1014 - 0x3f6  :  239 - 0xef
    "11111111", -- 1015 - 0x3f7  :  255 - 0xff
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "10101111", -- 1017 - 0x3f9  :  175 - 0xaf
    "01111111", -- 1018 - 0x3fa  :  127 - 0x7f
    "11111111", -- 1019 - 0x3fb  :  255 - 0xff
    "11111011", -- 1020 - 0x3fc  :  251 - 0xfb
    "11110101", -- 1021 - 0x3fd  :  245 - 0xf5
    "11101111", -- 1022 - 0x3fe  :  239 - 0xef
    "11111111", -- 1023 - 0x3ff  :  255 - 0xff
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x80
    "01111111", -- 1025 - 0x401  :  127 - 0x7f
    "00110000", -- 1026 - 0x402  :   48 - 0x30
    "00110000", -- 1027 - 0x403  :   48 - 0x30
    "00110000", -- 1028 - 0x404  :   48 - 0x30
    "01111111", -- 1029 - 0x405  :  127 - 0x7f
    "00110000", -- 1030 - 0x406  :   48 - 0x30
    "00110000", -- 1031 - 0x407  :   48 - 0x30
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Sprite 0x81
    "01111111", -- 1033 - 0x409  :  127 - 0x7f
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "01111111", -- 1035 - 0x40b  :  127 - 0x7f
    "01111111", -- 1036 - 0x40c  :  127 - 0x7f
    "00100000", -- 1037 - 0x40d  :   32 - 0x20
    "01000000", -- 1038 - 0x40e  :   64 - 0x40
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x82
    "11111110", -- 1041 - 0x411  :  254 - 0xfe
    "00001100", -- 1042 - 0x412  :   12 - 0xc
    "00001100", -- 1043 - 0x413  :   12 - 0xc
    "00001100", -- 1044 - 0x414  :   12 - 0xc
    "11111110", -- 1045 - 0x415  :  254 - 0xfe
    "00001100", -- 1046 - 0x416  :   12 - 0xc
    "00001100", -- 1047 - 0x417  :   12 - 0xc
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Sprite 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "11111111", -- 1051 - 0x41b  :  255 - 0xff
    "11111111", -- 1052 - 0x41c  :  255 - 0xff
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Sprite 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11101111", -- 1061 - 0x425  :  239 - 0xef
    "10111011", -- 1062 - 0x426  :  187 - 0xbb
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Sprite 0x85
    "11111110", -- 1065 - 0x429  :  254 - 0xfe
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "11111110", -- 1067 - 0x42b  :  254 - 0xfe
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "00001100", -- 1069 - 0x42d  :   12 - 0xc
    "00000010", -- 1070 - 0x42e  :    2 - 0x2
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Sprite 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x88
    "00000111", -- 1089 - 0x441  :    7 - 0x7
    "00011111", -- 1090 - 0x442  :   31 - 0x1f
    "00111100", -- 1091 - 0x443  :   60 - 0x3c
    "00110001", -- 1092 - 0x444  :   49 - 0x31
    "01110100", -- 1093 - 0x445  :  116 - 0x74
    "01100101", -- 1094 - 0x446  :  101 - 0x65
    "01101010", -- 1095 - 0x447  :  106 - 0x6a
    "01100100", -- 1096 - 0x448  :  100 - 0x64 -- Sprite 0x89
    "01101101", -- 1097 - 0x449  :  109 - 0x6d
    "01110010", -- 1098 - 0x44a  :  114 - 0x72
    "00110000", -- 1099 - 0x44b  :   48 - 0x30
    "00111100", -- 1100 - 0x44c  :   60 - 0x3c
    "00011111", -- 1101 - 0x44d  :   31 - 0x1f
    "00000111", -- 1102 - 0x44e  :    7 - 0x7
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x8a
    "11100000", -- 1105 - 0x451  :  224 - 0xe0
    "11111000", -- 1106 - 0x452  :  248 - 0xf8
    "00111100", -- 1107 - 0x453  :   60 - 0x3c
    "01001100", -- 1108 - 0x454  :   76 - 0x4c
    "01101110", -- 1109 - 0x455  :  110 - 0x6e
    "00100110", -- 1110 - 0x456  :   38 - 0x26
    "01000110", -- 1111 - 0x457  :   70 - 0x46
    "10010110", -- 1112 - 0x458  :  150 - 0x96 -- Sprite 0x8b
    "01100110", -- 1113 - 0x459  :  102 - 0x66
    "10101110", -- 1114 - 0x45a  :  174 - 0xae
    "01001100", -- 1115 - 0x45b  :   76 - 0x4c
    "00111100", -- 1116 - 0x45c  :   60 - 0x3c
    "11111000", -- 1117 - 0x45d  :  248 - 0xf8
    "11100000", -- 1118 - 0x45e  :  224 - 0xe0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x8c
    "00000111", -- 1121 - 0x461  :    7 - 0x7
    "00011111", -- 1122 - 0x462  :   31 - 0x1f
    "00111111", -- 1123 - 0x463  :   63 - 0x3f
    "00111111", -- 1124 - 0x464  :   63 - 0x3f
    "01111111", -- 1125 - 0x465  :  127 - 0x7f
    "01111111", -- 1126 - 0x466  :  127 - 0x7f
    "01111111", -- 1127 - 0x467  :  127 - 0x7f
    "01111111", -- 1128 - 0x468  :  127 - 0x7f -- Sprite 0x8d
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "01111111", -- 1130 - 0x46a  :  127 - 0x7f
    "00111111", -- 1131 - 0x46b  :   63 - 0x3f
    "00111111", -- 1132 - 0x46c  :   63 - 0x3f
    "00011111", -- 1133 - 0x46d  :   31 - 0x1f
    "00000111", -- 1134 - 0x46e  :    7 - 0x7
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Sprite 0x8e
    "11100000", -- 1137 - 0x471  :  224 - 0xe0
    "11111000", -- 1138 - 0x472  :  248 - 0xf8
    "11111100", -- 1139 - 0x473  :  252 - 0xfc
    "11111100", -- 1140 - 0x474  :  252 - 0xfc
    "11111110", -- 1141 - 0x475  :  254 - 0xfe
    "11111110", -- 1142 - 0x476  :  254 - 0xfe
    "11111110", -- 1143 - 0x477  :  254 - 0xfe
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- Sprite 0x8f
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111110", -- 1146 - 0x47a  :  254 - 0xfe
    "11111100", -- 1147 - 0x47b  :  252 - 0xfc
    "11111100", -- 1148 - 0x47c  :  252 - 0xfc
    "11111000", -- 1149 - 0x47d  :  248 - 0xf8
    "11100000", -- 1150 - 0x47e  :  224 - 0xe0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00010000", -- 1156 - 0x484  :   16 - 0x10
    "00011100", -- 1157 - 0x485  :   28 - 0x1c
    "00001110", -- 1158 - 0x486  :   14 - 0xe
    "00000111", -- 1159 - 0x487  :    7 - 0x7
    "00000011", -- 1160 - 0x488  :    3 - 0x3 -- Sprite 0x91
    "00000001", -- 1161 - 0x489  :    1 - 0x1
    "00110000", -- 1162 - 0x48a  :   48 - 0x30
    "00001111", -- 1163 - 0x48b  :   15 - 0xf
    "00000011", -- 1164 - 0x48c  :    3 - 0x3
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "01111111", -- 1166 - 0x48e  :  127 - 0x7f
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x92
    "01000010", -- 1169 - 0x491  :   66 - 0x42
    "01000010", -- 1170 - 0x492  :   66 - 0x42
    "01100110", -- 1171 - 0x493  :  102 - 0x66
    "01100110", -- 1172 - 0x494  :  102 - 0x66
    "01100110", -- 1173 - 0x495  :  102 - 0x66
    "11111110", -- 1174 - 0x496  :  254 - 0xfe
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "01111110", -- 1176 - 0x498  :  126 - 0x7e -- Sprite 0x93
    "01111110", -- 1177 - 0x499  :  126 - 0x7e
    "01111110", -- 1178 - 0x49a  :  126 - 0x7e
    "01111110", -- 1179 - 0x49b  :  126 - 0x7e
    "01111110", -- 1180 - 0x49c  :  126 - 0x7e
    "01111110", -- 1181 - 0x49d  :  126 - 0x7e
    "01111110", -- 1182 - 0x49e  :  126 - 0x7e
    "01111110", -- 1183 - 0x49f  :  126 - 0x7e
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00001000", -- 1188 - 0x4a4  :    8 - 0x8
    "00111000", -- 1189 - 0x4a5  :   56 - 0x38
    "01110000", -- 1190 - 0x4a6  :  112 - 0x70
    "11100000", -- 1191 - 0x4a7  :  224 - 0xe0
    "11000000", -- 1192 - 0x4a8  :  192 - 0xc0 -- Sprite 0x95
    "10000000", -- 1193 - 0x4a9  :  128 - 0x80
    "00001100", -- 1194 - 0x4aa  :   12 - 0xc
    "11110000", -- 1195 - 0x4ab  :  240 - 0xf0
    "11000000", -- 1196 - 0x4ac  :  192 - 0xc0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "11111110", -- 1198 - 0x4ae  :  254 - 0xfe
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "00111111", -- 1201 - 0x4b1  :   63 - 0x3f
    "01111111", -- 1202 - 0x4b2  :  127 - 0x7f
    "01111111", -- 1203 - 0x4b3  :  127 - 0x7f
    "01111111", -- 1204 - 0x4b4  :  127 - 0x7f
    "01111111", -- 1205 - 0x4b5  :  127 - 0x7f
    "01111111", -- 1206 - 0x4b6  :  127 - 0x7f
    "01111111", -- 1207 - 0x4b7  :  127 - 0x7f
    "01111111", -- 1208 - 0x4b8  :  127 - 0x7f -- Sprite 0x97
    "01111111", -- 1209 - 0x4b9  :  127 - 0x7f
    "00111111", -- 1210 - 0x4ba  :   63 - 0x3f
    "01111111", -- 1211 - 0x4bb  :  127 - 0x7f
    "01111111", -- 1212 - 0x4bc  :  127 - 0x7f
    "01111111", -- 1213 - 0x4bd  :  127 - 0x7f
    "01111111", -- 1214 - 0x4be  :  127 - 0x7f
    "01111111", -- 1215 - 0x4bf  :  127 - 0x7f
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x98
    "11011111", -- 1217 - 0x4c1  :  223 - 0xdf
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "10111111", -- 1226 - 0x4ca  :  191 - 0xbf
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "11111111", -- 1228 - 0x4cc  :  255 - 0xff
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "10111100", -- 1233 - 0x4d1  :  188 - 0xbc
    "11111110", -- 1234 - 0x4d2  :  254 - 0xfe
    "11111110", -- 1235 - 0x4d3  :  254 - 0xfe
    "11111110", -- 1236 - 0x4d4  :  254 - 0xfe
    "11111110", -- 1237 - 0x4d5  :  254 - 0xfe
    "11111110", -- 1238 - 0x4d6  :  254 - 0xfe
    "11111110", -- 1239 - 0x4d7  :  254 - 0xfe
    "11111110", -- 1240 - 0x4d8  :  254 - 0xfe -- Sprite 0x9b
    "11111110", -- 1241 - 0x4d9  :  254 - 0xfe
    "10111110", -- 1242 - 0x4da  :  190 - 0xbe
    "11111110", -- 1243 - 0x4db  :  254 - 0xfe
    "11111110", -- 1244 - 0x4dc  :  254 - 0xfe
    "11111110", -- 1245 - 0x4dd  :  254 - 0xfe
    "11111110", -- 1246 - 0x4de  :  254 - 0xfe
    "11111110", -- 1247 - 0x4df  :  254 - 0xfe
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Sprite 0x9c
    "00111111", -- 1249 - 0x4e1  :   63 - 0x3f
    "01011111", -- 1250 - 0x4e2  :   95 - 0x5f
    "01101111", -- 1251 - 0x4e3  :  111 - 0x6f
    "01110111", -- 1252 - 0x4e4  :  119 - 0x77
    "01111011", -- 1253 - 0x4e5  :  123 - 0x7b
    "00010101", -- 1254 - 0x4e6  :   21 - 0x15
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- Sprite 0x9d
    "10111110", -- 1257 - 0x4e9  :  190 - 0xbe
    "11011110", -- 1258 - 0x4ea  :  222 - 0xde
    "11101110", -- 1259 - 0x4eb  :  238 - 0xee
    "11110110", -- 1260 - 0x4ec  :  246 - 0xf6
    "11111010", -- 1261 - 0x4ed  :  250 - 0xfa
    "01010100", -- 1262 - 0x4ee  :   84 - 0x54
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x9e
    "10111111", -- 1265 - 0x4f1  :  191 - 0xbf
    "11011111", -- 1266 - 0x4f2  :  223 - 0xdf
    "11101111", -- 1267 - 0x4f3  :  239 - 0xef
    "11110111", -- 1268 - 0x4f4  :  247 - 0xf7
    "11111011", -- 1269 - 0x4f5  :  251 - 0xfb
    "01010101", -- 1270 - 0x4f6  :   85 - 0x55
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0xa0
    "01111111", -- 1281 - 0x501  :  127 - 0x7f
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000001", -- 1283 - 0x503  :    1 - 0x1
    "00000001", -- 1284 - 0x504  :    1 - 0x1
    "00000001", -- 1285 - 0x505  :    1 - 0x1
    "00000001", -- 1286 - 0x506  :    1 - 0x1
    "00000001", -- 1287 - 0x507  :    1 - 0x1
    "00000001", -- 1288 - 0x508  :    1 - 0x1 -- Sprite 0xa1
    "00000001", -- 1289 - 0x509  :    1 - 0x1
    "00000001", -- 1290 - 0x50a  :    1 - 0x1
    "00000001", -- 1291 - 0x50b  :    1 - 0x1
    "00000001", -- 1292 - 0x50c  :    1 - 0x1
    "00000001", -- 1293 - 0x50d  :    1 - 0x1
    "00000001", -- 1294 - 0x50e  :    1 - 0x1
    "00000001", -- 1295 - 0x50f  :    1 - 0x1
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Sprite 0xa2
    "11111110", -- 1297 - 0x511  :  254 - 0xfe
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "10000000", -- 1299 - 0x513  :  128 - 0x80
    "10000000", -- 1300 - 0x514  :  128 - 0x80
    "10000000", -- 1301 - 0x515  :  128 - 0x80
    "10000000", -- 1302 - 0x516  :  128 - 0x80
    "10000000", -- 1303 - 0x517  :  128 - 0x80
    "10000000", -- 1304 - 0x518  :  128 - 0x80 -- Sprite 0xa3
    "10000000", -- 1305 - 0x519  :  128 - 0x80
    "10000000", -- 1306 - 0x51a  :  128 - 0x80
    "10000000", -- 1307 - 0x51b  :  128 - 0x80
    "10000000", -- 1308 - 0x51c  :  128 - 0x80
    "10000000", -- 1309 - 0x51d  :  128 - 0x80
    "10000000", -- 1310 - 0x51e  :  128 - 0x80
    "10000000", -- 1311 - 0x51f  :  128 - 0x80
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0xa4
    "00110000", -- 1313 - 0x521  :   48 - 0x30
    "00111000", -- 1314 - 0x522  :   56 - 0x38
    "01111000", -- 1315 - 0x523  :  120 - 0x78
    "01111100", -- 1316 - 0x524  :  124 - 0x7c
    "01111101", -- 1317 - 0x525  :  125 - 0x7d
    "00011101", -- 1318 - 0x526  :   29 - 0x1d
    "00001101", -- 1319 - 0x527  :   13 - 0xd
    "00001101", -- 1320 - 0x528  :   13 - 0xd -- Sprite 0xa5
    "00011101", -- 1321 - 0x529  :   29 - 0x1d
    "00111101", -- 1322 - 0x52a  :   61 - 0x3d
    "00111111", -- 1323 - 0x52b  :   63 - 0x3f
    "00111111", -- 1324 - 0x52c  :   63 - 0x3f
    "00011111", -- 1325 - 0x52d  :   31 - 0x1f
    "00000001", -- 1326 - 0x52e  :    1 - 0x1
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "11100000", -- 1330 - 0x532  :  224 - 0xe0
    "11111000", -- 1331 - 0x533  :  248 - 0xf8
    "11111000", -- 1332 - 0x534  :  248 - 0xf8
    "11110000", -- 1333 - 0x535  :  240 - 0xf0
    "11000000", -- 1334 - 0x536  :  192 - 0xc0
    "11000000", -- 1335 - 0x537  :  192 - 0xc0
    "11000000", -- 1336 - 0x538  :  192 - 0xc0 -- Sprite 0xa7
    "11110000", -- 1337 - 0x539  :  240 - 0xf0
    "11110000", -- 1338 - 0x53a  :  240 - 0xf0
    "11000000", -- 1339 - 0x53b  :  192 - 0xc0
    "11000000", -- 1340 - 0x53c  :  192 - 0xc0
    "11000000", -- 1341 - 0x53d  :  192 - 0xc0
    "11000000", -- 1342 - 0x53e  :  192 - 0xc0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0xa8
    "01100000", -- 1345 - 0x541  :   96 - 0x60
    "01100000", -- 1346 - 0x542  :   96 - 0x60
    "01100000", -- 1347 - 0x543  :   96 - 0x60
    "01100000", -- 1348 - 0x544  :   96 - 0x60
    "01100000", -- 1349 - 0x545  :   96 - 0x60
    "01100000", -- 1350 - 0x546  :   96 - 0x60
    "01100000", -- 1351 - 0x547  :   96 - 0x60
    "01100000", -- 1352 - 0x548  :   96 - 0x60 -- Sprite 0xa9
    "01100000", -- 1353 - 0x549  :   96 - 0x60
    "01100000", -- 1354 - 0x54a  :   96 - 0x60
    "01100000", -- 1355 - 0x54b  :   96 - 0x60
    "01100000", -- 1356 - 0x54c  :   96 - 0x60
    "01100000", -- 1357 - 0x54d  :   96 - 0x60
    "01100000", -- 1358 - 0x54e  :   96 - 0x60
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Sprite 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000110", -- 1377 - 0x561  :    6 - 0x6
    "00000110", -- 1378 - 0x562  :    6 - 0x6
    "00000110", -- 1379 - 0x563  :    6 - 0x6
    "00000110", -- 1380 - 0x564  :    6 - 0x6
    "00000110", -- 1381 - 0x565  :    6 - 0x6
    "00000110", -- 1382 - 0x566  :    6 - 0x6
    "00000110", -- 1383 - 0x567  :    6 - 0x6
    "00000110", -- 1384 - 0x568  :    6 - 0x6 -- Sprite 0xad
    "00000110", -- 1385 - 0x569  :    6 - 0x6
    "00000110", -- 1386 - 0x56a  :    6 - 0x6
    "00000110", -- 1387 - 0x56b  :    6 - 0x6
    "00000110", -- 1388 - 0x56c  :    6 - 0x6
    "00000110", -- 1389 - 0x56d  :    6 - 0x6
    "00000110", -- 1390 - 0x56e  :    6 - 0x6
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000001", -- 1393 - 0x571  :    1 - 0x1
    "00000011", -- 1394 - 0x572  :    3 - 0x3
    "00000010", -- 1395 - 0x573  :    2 - 0x2
    "00000010", -- 1396 - 0x574  :    2 - 0x2
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000011", -- 1398 - 0x576  :    3 - 0x3
    "00000010", -- 1399 - 0x577  :    2 - 0x2
    "00000001", -- 1400 - 0x578  :    1 - 0x1 -- Sprite 0xaf
    "00000011", -- 1401 - 0x579  :    3 - 0x3
    "00000101", -- 1402 - 0x57a  :    5 - 0x5
    "00000100", -- 1403 - 0x57b  :    4 - 0x4
    "00000101", -- 1404 - 0x57c  :    5 - 0x5
    "00001101", -- 1405 - 0x57d  :   13 - 0xd
    "00001100", -- 1406 - 0x57e  :   12 - 0xc
    "00000001", -- 1407 - 0x57f  :    1 - 0x1
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "01000000", -- 1410 - 0x582  :   64 - 0x40
    "11110000", -- 1411 - 0x583  :  240 - 0xf0
    "11101000", -- 1412 - 0x584  :  232 - 0xe8
    "10010000", -- 1413 - 0x585  :  144 - 0x90
    "01010000", -- 1414 - 0x586  :   80 - 0x50
    "11010000", -- 1415 - 0x587  :  208 - 0xd0
    "11111000", -- 1416 - 0x588  :  248 - 0xf8 -- Sprite 0xb1
    "11000000", -- 1417 - 0x589  :  192 - 0xc0
    "11100000", -- 1418 - 0x58a  :  224 - 0xe0
    "01000000", -- 1419 - 0x58b  :   64 - 0x40
    "10000000", -- 1420 - 0x58c  :  128 - 0x80
    "11000000", -- 1421 - 0x58d  :  192 - 0xc0
    "11100000", -- 1422 - 0x58e  :  224 - 0xe0
    "01110000", -- 1423 - 0x58f  :  112 - 0x70
    "00000001", -- 1424 - 0x590  :    1 - 0x1 -- Sprite 0xb2
    "00001101", -- 1425 - 0x591  :   13 - 0xd
    "00001101", -- 1426 - 0x592  :   13 - 0xd
    "00000011", -- 1427 - 0x593  :    3 - 0x3
    "00000011", -- 1428 - 0x594  :    3 - 0x3
    "00000111", -- 1429 - 0x595  :    7 - 0x7
    "00000111", -- 1430 - 0x596  :    7 - 0x7
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00111111", -- 1432 - 0x598  :   63 - 0x3f -- Sprite 0xb3
    "00111111", -- 1433 - 0x599  :   63 - 0x3f
    "00111111", -- 1434 - 0x59a  :   63 - 0x3f
    "00111111", -- 1435 - 0x59b  :   63 - 0x3f
    "00111111", -- 1436 - 0x59c  :   63 - 0x3f
    "00111111", -- 1437 - 0x59d  :   63 - 0x3f
    "00110101", -- 1438 - 0x59e  :   53 - 0x35
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "10110000", -- 1440 - 0x5a0  :  176 - 0xb0 -- Sprite 0xb4
    "11000000", -- 1441 - 0x5a1  :  192 - 0xc0
    "11100000", -- 1442 - 0x5a2  :  224 - 0xe0
    "11100000", -- 1443 - 0x5a3  :  224 - 0xe0
    "11110000", -- 1444 - 0x5a4  :  240 - 0xf0
    "11110000", -- 1445 - 0x5a5  :  240 - 0xf0
    "11110000", -- 1446 - 0x5a6  :  240 - 0xf0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "11111100", -- 1448 - 0x5a8  :  252 - 0xfc -- Sprite 0xb5
    "11111000", -- 1449 - 0x5a9  :  248 - 0xf8
    "11111100", -- 1450 - 0x5aa  :  252 - 0xfc
    "11111000", -- 1451 - 0x5ab  :  248 - 0xf8
    "11111100", -- 1452 - 0x5ac  :  252 - 0xfc
    "11111000", -- 1453 - 0x5ad  :  248 - 0xf8
    "01010100", -- 1454 - 0x5ae  :   84 - 0x54
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "01111111", -- 1457 - 0x5b1  :  127 - 0x7f
    "01111111", -- 1458 - 0x5b2  :  127 - 0x7f
    "01111111", -- 1459 - 0x5b3  :  127 - 0x7f
    "01111111", -- 1460 - 0x5b4  :  127 - 0x7f
    "01111111", -- 1461 - 0x5b5  :  127 - 0x7f
    "01101010", -- 1462 - 0x5b6  :  106 - 0x6a
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- Sprite 0xb7
    "01111011", -- 1465 - 0x5b9  :  123 - 0x7b
    "01110011", -- 1466 - 0x5ba  :  115 - 0x73
    "01111011", -- 1467 - 0x5bb  :  123 - 0x7b
    "01110011", -- 1468 - 0x5bc  :  115 - 0x73
    "01111011", -- 1469 - 0x5bd  :  123 - 0x7b
    "01010011", -- 1470 - 0x5be  :   83 - 0x53
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0xb8
    "11011110", -- 1473 - 0x5c1  :  222 - 0xde
    "10011110", -- 1474 - 0x5c2  :  158 - 0x9e
    "11011100", -- 1475 - 0x5c3  :  220 - 0xdc
    "10011110", -- 1476 - 0x5c4  :  158 - 0x9e
    "11011100", -- 1477 - 0x5c5  :  220 - 0xdc
    "10011010", -- 1478 - 0x5c6  :  154 - 0x9a
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- Sprite 0xb9
    "11111110", -- 1481 - 0x5c9  :  254 - 0xfe
    "11111100", -- 1482 - 0x5ca  :  252 - 0xfc
    "11111110", -- 1483 - 0x5cb  :  254 - 0xfe
    "11111100", -- 1484 - 0x5cc  :  252 - 0xfc
    "11111110", -- 1485 - 0x5cd  :  254 - 0xfe
    "01010100", -- 1486 - 0x5ce  :   84 - 0x54
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0xba
    "01111111", -- 1489 - 0x5d1  :  127 - 0x7f
    "01111111", -- 1490 - 0x5d2  :  127 - 0x7f
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "01111111", -- 1492 - 0x5d4  :  127 - 0x7f
    "01111111", -- 1493 - 0x5d5  :  127 - 0x7f
    "01101010", -- 1494 - 0x5d6  :  106 - 0x6a
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0xbc
    "11111110", -- 1505 - 0x5e1  :  254 - 0xfe
    "11111110", -- 1506 - 0x5e2  :  254 - 0xfe
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "10011110", -- 1508 - 0x5e4  :  158 - 0x9e
    "11011100", -- 1509 - 0x5e5  :  220 - 0xdc
    "10011010", -- 1510 - 0x5e6  :  154 - 0x9a
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- Sprite 0xc5
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000001", -- 1579 - 0x62b  :    1 - 0x1
    "00000111", -- 1580 - 0x62c  :    7 - 0x7
    "00001111", -- 1581 - 0x62d  :   15 - 0xf
    "00001111", -- 1582 - 0x62e  :   15 - 0xf
    "00011111", -- 1583 - 0x62f  :   31 - 0x1f
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0xc6
    "00011111", -- 1585 - 0x631  :   31 - 0x1f
    "01111111", -- 1586 - 0x632  :  127 - 0x7f
    "11111111", -- 1587 - 0x633  :  255 - 0xff
    "11111111", -- 1588 - 0x634  :  255 - 0xff
    "11111111", -- 1589 - 0x635  :  255 - 0xff
    "11111111", -- 1590 - 0x636  :  255 - 0xff
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "00011111", -- 1592 - 0x638  :   31 - 0x1f -- Sprite 0xc7
    "00111111", -- 1593 - 0x639  :   63 - 0x3f
    "00111111", -- 1594 - 0x63a  :   63 - 0x3f
    "01111111", -- 1595 - 0x63b  :  127 - 0x7f
    "01111111", -- 1596 - 0x63c  :  127 - 0x7f
    "01111111", -- 1597 - 0x63d  :  127 - 0x7f
    "01111111", -- 1598 - 0x63e  :  127 - 0x7f
    "01111111", -- 1599 - 0x63f  :  127 - 0x7f
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "11111111", -- 1601 - 0x641  :  255 - 0xff
    "11111111", -- 1602 - 0x642  :  255 - 0xff
    "11111111", -- 1603 - 0x643  :  255 - 0xff
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "11111111", -- 1605 - 0x645  :  255 - 0xff
    "11111111", -- 1606 - 0x646  :  255 - 0xff
    "11111111", -- 1607 - 0x647  :  255 - 0xff
    "11101000", -- 1608 - 0x648  :  232 - 0xe8 -- Sprite 0xc9
    "11010100", -- 1609 - 0x649  :  212 - 0xd4
    "11101000", -- 1610 - 0x64a  :  232 - 0xe8
    "11010100", -- 1611 - 0x64b  :  212 - 0xd4
    "11101010", -- 1612 - 0x64c  :  234 - 0xea
    "11010100", -- 1613 - 0x64d  :  212 - 0xd4
    "11101010", -- 1614 - 0x64e  :  234 - 0xea
    "11010100", -- 1615 - 0x64f  :  212 - 0xd4
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000101", -- 1636 - 0x664  :    5 - 0x5
    "00000010", -- 1637 - 0x665  :    2 - 0x2
    "00000001", -- 1638 - 0x666  :    1 - 0x1
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "10000000", -- 1643 - 0x66b  :  128 - 0x80
    "01010000", -- 1644 - 0x66c  :   80 - 0x50
    "10100000", -- 1645 - 0x66d  :  160 - 0xa0
    "01000000", -- 1646 - 0x66e  :   64 - 0x40
    "10000000", -- 1647 - 0x66f  :  128 - 0x80
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00110000", -- 1652 - 0x674  :   48 - 0x30
    "01111111", -- 1653 - 0x675  :  127 - 0x7f
    "00110000", -- 1654 - 0x676  :   48 - 0x30
    "00110000", -- 1655 - 0x677  :   48 - 0x30
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00001100", -- 1660 - 0x67c  :   12 - 0xc
    "11111110", -- 1661 - 0x67d  :  254 - 0xfe
    "00001100", -- 1662 - 0x67e  :   12 - 0xc
    "00001100", -- 1663 - 0x67f  :   12 - 0xc
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Sprite 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000111", -- 1680 - 0x690  :    7 - 0x7 -- Sprite 0xd2
    "00000111", -- 1681 - 0x691  :    7 - 0x7
    "00000111", -- 1682 - 0x692  :    7 - 0x7
    "00000111", -- 1683 - 0x693  :    7 - 0x7
    "00000111", -- 1684 - 0x694  :    7 - 0x7
    "00000111", -- 1685 - 0x695  :    7 - 0x7
    "00000111", -- 1686 - 0x696  :    7 - 0x7
    "00000111", -- 1687 - 0x697  :    7 - 0x7
    "11100000", -- 1688 - 0x698  :  224 - 0xe0 -- Sprite 0xd3
    "11100000", -- 1689 - 0x699  :  224 - 0xe0
    "11000000", -- 1690 - 0x69a  :  192 - 0xc0
    "11100000", -- 1691 - 0x69b  :  224 - 0xe0
    "10100000", -- 1692 - 0x69c  :  160 - 0xa0
    "11100000", -- 1693 - 0x69d  :  224 - 0xe0
    "11000000", -- 1694 - 0x69e  :  192 - 0xc0
    "11100000", -- 1695 - 0x69f  :  224 - 0xe0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "11111000", -- 1705 - 0x6a9  :  248 - 0xf8
    "11111110", -- 1706 - 0x6aa  :  254 - 0xfe
    "11111111", -- 1707 - 0x6ab  :  255 - 0xff
    "11111111", -- 1708 - 0x6ac  :  255 - 0xff
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "10000000", -- 1715 - 0x6b3  :  128 - 0x80
    "10100000", -- 1716 - 0x6b4  :  160 - 0xa0
    "01010000", -- 1717 - 0x6b5  :   80 - 0x50
    "10100000", -- 1718 - 0x6b6  :  160 - 0xa0
    "11010000", -- 1719 - 0x6b7  :  208 - 0xd0
    "01111111", -- 1720 - 0x6b8  :  127 - 0x7f -- Sprite 0xd7
    "01111111", -- 1721 - 0x6b9  :  127 - 0x7f
    "01111111", -- 1722 - 0x6ba  :  127 - 0x7f
    "00111111", -- 1723 - 0x6bb  :   63 - 0x3f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00001111", -- 1725 - 0x6bd  :   15 - 0xf
    "00000111", -- 1726 - 0x6be  :    7 - 0x7
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11111111", -- 1732 - 0x6c4  :  255 - 0xff
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111111", -- 1734 - 0x6c6  :  255 - 0xff
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "11101010", -- 1736 - 0x6c8  :  234 - 0xea -- Sprite 0xd9
    "11010100", -- 1737 - 0x6c9  :  212 - 0xd4
    "11101010", -- 1738 - 0x6ca  :  234 - 0xea
    "11010100", -- 1739 - 0x6cb  :  212 - 0xd4
    "10101000", -- 1740 - 0x6cc  :  168 - 0xa8
    "01010000", -- 1741 - 0x6cd  :   80 - 0x50
    "10100000", -- 1742 - 0x6ce  :  160 - 0xa0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00001100", -- 1746 - 0x6d2  :   12 - 0xc
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Sprite 0xdb
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "10000000", -- 1754 - 0x6da  :  128 - 0x80
    "10000000", -- 1755 - 0x6db  :  128 - 0x80
    "10011000", -- 1756 - 0x6dc  :  152 - 0x98
    "10000000", -- 1757 - 0x6dd  :  128 - 0x80
    "10000000", -- 1758 - 0x6de  :  128 - 0x80
    "10000000", -- 1759 - 0x6df  :  128 - 0x80
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000010", -- 1764 - 0x6e4  :    2 - 0x2
    "00000011", -- 1765 - 0x6e5  :    3 - 0x3
    "00000011", -- 1766 - 0x6e6  :    3 - 0x3
    "00000001", -- 1767 - 0x6e7  :    1 - 0x1
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "10100000", -- 1772 - 0x6ec  :  160 - 0xa0
    "11100000", -- 1773 - 0x6ed  :  224 - 0xe0
    "11100000", -- 1774 - 0x6ee  :  224 - 0xe0
    "11000000", -- 1775 - 0x6ef  :  192 - 0xc0
    "00110000", -- 1776 - 0x6f0  :   48 - 0x30 -- Sprite 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00110000", -- 1778 - 0x6f2  :   48 - 0x30
    "00110000", -- 1779 - 0x6f3  :   48 - 0x30
    "00110000", -- 1780 - 0x6f4  :   48 - 0x30
    "00110000", -- 1781 - 0x6f5  :   48 - 0x30
    "00110000", -- 1782 - 0x6f6  :   48 - 0x30
    "00110000", -- 1783 - 0x6f7  :   48 - 0x30
    "00001100", -- 1784 - 0x6f8  :   12 - 0xc -- Sprite 0xdf
    "11111110", -- 1785 - 0x6f9  :  254 - 0xfe
    "00001100", -- 1786 - 0x6fa  :   12 - 0xc
    "00001100", -- 1787 - 0x6fb  :   12 - 0xc
    "00001100", -- 1788 - 0x6fc  :   12 - 0xc
    "00001100", -- 1789 - 0x6fd  :   12 - 0xc
    "00001100", -- 1790 - 0x6fe  :   12 - 0xc
    "00001100", -- 1791 - 0x6ff  :   12 - 0xc
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- Sprite 0xe1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0xe2
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- Sprite 0xe3
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Sprite 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Sprite 0xf1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Sprite 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Sprite 0xf5
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
          -- Background pattern Table
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Background 0x0
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000011", -- 2050 - 0x802  :    3 - 0x3
    "00000001", -- 2051 - 0x803  :    1 - 0x1
    "00000001", -- 2052 - 0x804  :    1 - 0x1
    "00000000", -- 2053 - 0x805  :    0 - 0x0
    "00000011", -- 2054 - 0x806  :    3 - 0x3
    "00000001", -- 2055 - 0x807  :    1 - 0x1
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- Background 0x1
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00111000", -- 2058 - 0x80a  :   56 - 0x38
    "10110100", -- 2059 - 0x80b  :  180 - 0xb4
    "10101000", -- 2060 - 0x80c  :  168 - 0xa8
    "11010100", -- 2061 - 0x80d  :  212 - 0xd4
    "01110100", -- 2062 - 0x80e  :  116 - 0x74
    "01111110", -- 2063 - 0x80f  :  126 - 0x7e
    "00111000", -- 2064 - 0x810  :   56 - 0x38 -- Background 0x2
    "01111000", -- 2065 - 0x811  :  120 - 0x78
    "01111100", -- 2066 - 0x812  :  124 - 0x7c
    "01111110", -- 2067 - 0x813  :  126 - 0x7e
    "01111110", -- 2068 - 0x814  :  126 - 0x7e
    "01111110", -- 2069 - 0x815  :  126 - 0x7e
    "00111110", -- 2070 - 0x816  :   62 - 0x3e
    "00011110", -- 2071 - 0x817  :   30 - 0x1e
    "11110110", -- 2072 - 0x818  :  246 - 0xf6 -- Background 0x3
    "11110000", -- 2073 - 0x819  :  240 - 0xf0
    "00111000", -- 2074 - 0x81a  :   56 - 0x38
    "11010000", -- 2075 - 0x81b  :  208 - 0xd0
    "11100000", -- 2076 - 0x81c  :  224 - 0xe0
    "01110000", -- 2077 - 0x81d  :  112 - 0x70
    "10111000", -- 2078 - 0x81e  :  184 - 0xb8
    "01000000", -- 2079 - 0x81f  :   64 - 0x40
    "00011100", -- 2080 - 0x820  :   28 - 0x1c -- Background 0x4
    "00011100", -- 2081 - 0x821  :   28 - 0x1c
    "00011110", -- 2082 - 0x822  :   30 - 0x1e
    "00011111", -- 2083 - 0x823  :   31 - 0x1f
    "00001100", -- 2084 - 0x824  :   12 - 0xc
    "00000000", -- 2085 - 0x825  :    0 - 0x0
    "00000000", -- 2086 - 0x826  :    0 - 0x0
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "10101000", -- 2088 - 0x828  :  168 - 0xa8 -- Background 0x5
    "01010000", -- 2089 - 0x829  :   80 - 0x50
    "10101000", -- 2090 - 0x82a  :  168 - 0xa8
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "01100000", -- 2092 - 0x82c  :   96 - 0x60
    "01100000", -- 2093 - 0x82d  :   96 - 0x60
    "01110000", -- 2094 - 0x82e  :  112 - 0x70
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00011100", -- 2096 - 0x830  :   28 - 0x1c -- Background 0x6
    "00011100", -- 2097 - 0x831  :   28 - 0x1c
    "00011110", -- 2098 - 0x832  :   30 - 0x1e
    "00011111", -- 2099 - 0x833  :   31 - 0x1f
    "00001100", -- 2100 - 0x834  :   12 - 0xc
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000001", -- 2102 - 0x836  :    1 - 0x1
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "10101000", -- 2104 - 0x838  :  168 - 0xa8 -- Background 0x7
    "01010000", -- 2105 - 0x839  :   80 - 0x50
    "10101000", -- 2106 - 0x83a  :  168 - 0xa8
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "01011000", -- 2108 - 0x83c  :   88 - 0x58
    "11011000", -- 2109 - 0x83d  :  216 - 0xd8
    "10001100", -- 2110 - 0x83e  :  140 - 0x8c
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00011100", -- 2112 - 0x840  :   28 - 0x1c -- Background 0x8
    "00011100", -- 2113 - 0x841  :   28 - 0x1c
    "00011110", -- 2114 - 0x842  :   30 - 0x1e
    "00011111", -- 2115 - 0x843  :   31 - 0x1f
    "00001100", -- 2116 - 0x844  :   12 - 0xc
    "00000000", -- 2117 - 0x845  :    0 - 0x0
    "00000000", -- 2118 - 0x846  :    0 - 0x0
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "10101000", -- 2120 - 0x848  :  168 - 0xa8 -- Background 0x9
    "01010100", -- 2121 - 0x849  :   84 - 0x54
    "10101000", -- 2122 - 0x84a  :  168 - 0xa8
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "01101110", -- 2124 - 0x84c  :  110 - 0x6e
    "11000000", -- 2125 - 0x84d  :  192 - 0xc0
    "10000000", -- 2126 - 0x84e  :  128 - 0x80
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00011100", -- 2128 - 0x850  :   28 - 0x1c -- Background 0xa
    "00011100", -- 2129 - 0x851  :   28 - 0x1c
    "00011110", -- 2130 - 0x852  :   30 - 0x1e
    "00011111", -- 2131 - 0x853  :   31 - 0x1f
    "00001100", -- 2132 - 0x854  :   12 - 0xc
    "00000001", -- 2133 - 0x855  :    1 - 0x1
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "10101000", -- 2136 - 0x858  :  168 - 0xa8 -- Background 0xb
    "01010100", -- 2137 - 0x859  :   84 - 0x54
    "10101000", -- 2138 - 0x85a  :  168 - 0xa8
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "11011000", -- 2140 - 0x85c  :  216 - 0xd8
    "11011100", -- 2141 - 0x85d  :  220 - 0xdc
    "00001100", -- 2142 - 0x85e  :   12 - 0xc
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "11110110", -- 2144 - 0x860  :  246 - 0xf6 -- Background 0xc
    "11110000", -- 2145 - 0x861  :  240 - 0xf0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "11111100", -- 2147 - 0x863  :  252 - 0xfc
    "11111000", -- 2148 - 0x864  :  248 - 0xf8
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "10101000", -- 2150 - 0x866  :  168 - 0xa8
    "01010100", -- 2151 - 0x867  :   84 - 0x54
    "00111000", -- 2152 - 0x868  :   56 - 0x38 -- Background 0xd
    "01111000", -- 2153 - 0x869  :  120 - 0x78
    "01111100", -- 2154 - 0x86a  :  124 - 0x7c
    "01111101", -- 2155 - 0x86b  :  125 - 0x7d
    "01111101", -- 2156 - 0x86c  :  125 - 0x7d
    "01111011", -- 2157 - 0x86d  :  123 - 0x7b
    "00111011", -- 2158 - 0x86e  :   59 - 0x3b
    "00011011", -- 2159 - 0x86f  :   27 - 0x1b
    "11110110", -- 2160 - 0x870  :  246 - 0xf6 -- Background 0xe
    "11110000", -- 2161 - 0x871  :  240 - 0xf0
    "01111000", -- 2162 - 0x872  :  120 - 0x78
    "01110000", -- 2163 - 0x873  :  112 - 0x70
    "10100000", -- 2164 - 0x874  :  160 - 0xa0
    "10010000", -- 2165 - 0x875  :  144 - 0x90
    "00101000", -- 2166 - 0x876  :   40 - 0x28
    "01010100", -- 2167 - 0x877  :   84 - 0x54
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- Background 0xf
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000011", -- 2170 - 0x87a  :    3 - 0x3
    "00000001", -- 2171 - 0x87b  :    1 - 0x1
    "00000001", -- 2172 - 0x87c  :    1 - 0x1
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000011", -- 2174 - 0x87e  :    3 - 0x3
    "00000001", -- 2175 - 0x87f  :    1 - 0x1
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Background 0x10
    "00000011", -- 2177 - 0x881  :    3 - 0x3
    "00001111", -- 2178 - 0x882  :   15 - 0xf
    "00001111", -- 2179 - 0x883  :   15 - 0xf
    "00001111", -- 2180 - 0x884  :   15 - 0xf
    "00011111", -- 2181 - 0x885  :   31 - 0x1f
    "00011111", -- 2182 - 0x886  :   31 - 0x1f
    "00011110", -- 2183 - 0x887  :   30 - 0x1e
    "00110110", -- 2184 - 0x888  :   54 - 0x36 -- Background 0x11
    "10110000", -- 2185 - 0x889  :  176 - 0xb0
    "10111000", -- 2186 - 0x88a  :  184 - 0xb8
    "10010000", -- 2187 - 0x88b  :  144 - 0x90
    "10100000", -- 2188 - 0x88c  :  160 - 0xa0
    "01110000", -- 2189 - 0x88d  :  112 - 0x70
    "00111000", -- 2190 - 0x88e  :   56 - 0x38
    "01000000", -- 2191 - 0x88f  :   64 - 0x40
    "00011100", -- 2192 - 0x890  :   28 - 0x1c -- Background 0x12
    "00011100", -- 2193 - 0x891  :   28 - 0x1c
    "00011110", -- 2194 - 0x892  :   30 - 0x1e
    "00011111", -- 2195 - 0x893  :   31 - 0x1f
    "00001100", -- 2196 - 0x894  :   12 - 0xc
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000000", -- 2200 - 0x898  :    0 - 0x0 -- Background 0x13
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000011", -- 2203 - 0x89b  :    3 - 0x3
    "00000111", -- 2204 - 0x89c  :    7 - 0x7
    "00001111", -- 2205 - 0x89d  :   15 - 0xf
    "00001111", -- 2206 - 0x89e  :   15 - 0xf
    "00011111", -- 2207 - 0x89f  :   31 - 0x1f
    "11110110", -- 2208 - 0x8a0  :  246 - 0xf6 -- Background 0x14
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "11111000", -- 2210 - 0x8a2  :  248 - 0xf8
    "11111110", -- 2211 - 0x8a3  :  254 - 0xfe
    "11111110", -- 2212 - 0x8a4  :  254 - 0xfe
    "11111110", -- 2213 - 0x8a5  :  254 - 0xfe
    "11111000", -- 2214 - 0x8a6  :  248 - 0xf8
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "00000011", -- 2216 - 0x8a8  :    3 - 0x3 -- Background 0x15
    "00000011", -- 2217 - 0x8a9  :    3 - 0x3
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000011", -- 2219 - 0x8ab  :    3 - 0x3
    "00000011", -- 2220 - 0x8ac  :    3 - 0x3
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00001111", -- 2222 - 0x8ae  :   15 - 0xf
    "00111111", -- 2223 - 0x8af  :   63 - 0x3f
    "11011000", -- 2224 - 0x8b0  :  216 - 0xd8 -- Background 0x16
    "11000000", -- 2225 - 0x8b1  :  192 - 0xc0
    "11100000", -- 2226 - 0x8b2  :  224 - 0xe0
    "01000000", -- 2227 - 0x8b3  :   64 - 0x40
    "10000000", -- 2228 - 0x8b4  :  128 - 0x80
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "11100000", -- 2230 - 0x8b6  :  224 - 0xe0
    "11111100", -- 2231 - 0x8b7  :  252 - 0xfc
    "01111111", -- 2232 - 0x8b8  :  127 - 0x7f -- Background 0x17
    "01111111", -- 2233 - 0x8b9  :  127 - 0x7f
    "01111111", -- 2234 - 0x8ba  :  127 - 0x7f
    "01111100", -- 2235 - 0x8bb  :  124 - 0x7c
    "00110000", -- 2236 - 0x8bc  :   48 - 0x30
    "00000001", -- 2237 - 0x8bd  :    1 - 0x1
    "00000001", -- 2238 - 0x8be  :    1 - 0x1
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "11111100", -- 2240 - 0x8c0  :  252 - 0xfc -- Background 0x18
    "11111110", -- 2241 - 0x8c1  :  254 - 0xfe
    "11111100", -- 2242 - 0x8c2  :  252 - 0xfc
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000000", -- 2244 - 0x8c4  :    0 - 0x0
    "10000000", -- 2245 - 0x8c5  :  128 - 0x80
    "11000000", -- 2246 - 0x8c6  :  192 - 0xc0
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "00000111", -- 2248 - 0x8c8  :    7 - 0x7 -- Background 0x19
    "00000111", -- 2249 - 0x8c9  :    7 - 0x7
    "00000001", -- 2250 - 0x8ca  :    1 - 0x1
    "00000110", -- 2251 - 0x8cb  :    6 - 0x6
    "00000111", -- 2252 - 0x8cc  :    7 - 0x7
    "00000110", -- 2253 - 0x8cd  :    6 - 0x6
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00001111", -- 2255 - 0x8cf  :   15 - 0xf
    "10110000", -- 2256 - 0x8d0  :  176 - 0xb0 -- Background 0x1a
    "10000000", -- 2257 - 0x8d1  :  128 - 0x80
    "11000000", -- 2258 - 0x8d2  :  192 - 0xc0
    "10000000", -- 2259 - 0x8d3  :  128 - 0x80
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "11100000", -- 2263 - 0x8d7  :  224 - 0xe0
    "00111111", -- 2264 - 0x8d8  :   63 - 0x3f -- Background 0x1b
    "00111111", -- 2265 - 0x8d9  :   63 - 0x3f
    "01111111", -- 2266 - 0x8da  :  127 - 0x7f
    "01111111", -- 2267 - 0x8db  :  127 - 0x7f
    "00111111", -- 2268 - 0x8dc  :   63 - 0x3f
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000011", -- 2270 - 0x8de  :    3 - 0x3
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "11111111", -- 2272 - 0x8e0  :  255 - 0xff -- Background 0x1c
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11111111", -- 2274 - 0x8e2  :  255 - 0xff
    "11111111", -- 2275 - 0x8e3  :  255 - 0xff
    "11111111", -- 2276 - 0x8e4  :  255 - 0xff
    "00000000", -- 2277 - 0x8e5  :    0 - 0x0
    "10000000", -- 2278 - 0x8e6  :  128 - 0x80
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- Background 0x1d
    "11000000", -- 2281 - 0x8e9  :  192 - 0xc0
    "11000000", -- 2282 - 0x8ea  :  192 - 0xc0
    "11000000", -- 2283 - 0x8eb  :  192 - 0xc0
    "10000000", -- 2284 - 0x8ec  :  128 - 0x80
    "00000000", -- 2285 - 0x8ed  :    0 - 0x0
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "11100000", -- 2288 - 0x8f0  :  224 - 0xe0 -- Background 0x1e
    "10011100", -- 2289 - 0x8f1  :  156 - 0x9c
    "00111000", -- 2290 - 0x8f2  :   56 - 0x38
    "11100000", -- 2291 - 0x8f3  :  224 - 0xe0
    "11001000", -- 2292 - 0x8f4  :  200 - 0xc8
    "00010100", -- 2293 - 0x8f5  :   20 - 0x14
    "10101000", -- 2294 - 0x8f6  :  168 - 0xa8
    "01010100", -- 2295 - 0x8f7  :   84 - 0x54
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0 -- Background 0x1f
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00111000", -- 2298 - 0x8fa  :   56 - 0x38
    "10110100", -- 2299 - 0x8fb  :  180 - 0xb4
    "10101000", -- 2300 - 0x8fc  :  168 - 0xa8
    "11010100", -- 2301 - 0x8fd  :  212 - 0xd4
    "01110100", -- 2302 - 0x8fe  :  116 - 0x74
    "00011110", -- 2303 - 0x8ff  :   30 - 0x1e
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x20
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00001100", -- 2306 - 0x902  :   12 - 0xc
    "00000111", -- 2307 - 0x903  :    7 - 0x7
    "00001111", -- 2308 - 0x904  :   15 - 0xf
    "00000111", -- 2309 - 0x905  :    7 - 0x7
    "00001111", -- 2310 - 0x906  :   15 - 0xf
    "00001111", -- 2311 - 0x907  :   15 - 0xf
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- Background 0x21
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00110000", -- 2314 - 0x90a  :   48 - 0x30
    "11100000", -- 2315 - 0x90b  :  224 - 0xe0
    "11110000", -- 2316 - 0x90c  :  240 - 0xf0
    "11100000", -- 2317 - 0x90d  :  224 - 0xe0
    "11110000", -- 2318 - 0x90e  :  240 - 0xf0
    "11110000", -- 2319 - 0x90f  :  240 - 0xf0
    "00000111", -- 2320 - 0x910  :    7 - 0x7 -- Background 0x22
    "00000011", -- 2321 - 0x911  :    3 - 0x3
    "00011000", -- 2322 - 0x912  :   24 - 0x18
    "00010101", -- 2323 - 0x913  :   21 - 0x15
    "00000010", -- 2324 - 0x914  :    2 - 0x2
    "00000101", -- 2325 - 0x915  :    5 - 0x5
    "00000010", -- 2326 - 0x916  :    2 - 0x2
    "00000100", -- 2327 - 0x917  :    4 - 0x4
    "11100000", -- 2328 - 0x918  :  224 - 0xe0 -- Background 0x23
    "11000000", -- 2329 - 0x919  :  192 - 0xc0
    "00111100", -- 2330 - 0x91a  :   60 - 0x3c
    "01111100", -- 2331 - 0x91b  :  124 - 0x7c
    "01111100", -- 2332 - 0x91c  :  124 - 0x7c
    "01111100", -- 2333 - 0x91d  :  124 - 0x7c
    "11101100", -- 2334 - 0x91e  :  236 - 0xec
    "11100000", -- 2335 - 0x91f  :  224 - 0xe0
    "00000010", -- 2336 - 0x920  :    2 - 0x2 -- Background 0x24
    "00000101", -- 2337 - 0x921  :    5 - 0x5
    "00001011", -- 2338 - 0x922  :   11 - 0xb
    "00001011", -- 2339 - 0x923  :   11 - 0xb
    "00001101", -- 2340 - 0x924  :   13 - 0xd
    "00011000", -- 2341 - 0x925  :   24 - 0x18
    "00111000", -- 2342 - 0x926  :   56 - 0x38
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "11100000", -- 2344 - 0x928  :  224 - 0xe0 -- Background 0x25
    "11100000", -- 2345 - 0x929  :  224 - 0xe0
    "11100000", -- 2346 - 0x92a  :  224 - 0xe0
    "11010000", -- 2347 - 0x92b  :  208 - 0xd0
    "10111000", -- 2348 - 0x92c  :  184 - 0xb8
    "00111000", -- 2349 - 0x92d  :   56 - 0x38
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "00000000", -- 2353 - 0x931  :    0 - 0x0
    "00000000", -- 2354 - 0x932  :    0 - 0x0
    "00000000", -- 2355 - 0x933  :    0 - 0x0
    "00000000", -- 2356 - 0x934  :    0 - 0x0
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0 -- Background 0x27
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "00000000", -- 2362 - 0x93a  :    0 - 0x0
    "00000000", -- 2363 - 0x93b  :    0 - 0x0
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00000000", -- 2372 - 0x944  :    0 - 0x0
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00011111", -- 2376 - 0x948  :   31 - 0x1f -- Background 0x29
    "00011111", -- 2377 - 0x949  :   31 - 0x1f
    "00011111", -- 2378 - 0x94a  :   31 - 0x1f
    "00011111", -- 2379 - 0x94b  :   31 - 0x1f
    "00001100", -- 2380 - 0x94c  :   12 - 0xc
    "00000000", -- 2381 - 0x94d  :    0 - 0x0
    "00000001", -- 2382 - 0x94e  :    1 - 0x1
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00011111", -- 2384 - 0x950  :   31 - 0x1f -- Background 0x2a
    "00011111", -- 2385 - 0x951  :   31 - 0x1f
    "00011111", -- 2386 - 0x952  :   31 - 0x1f
    "00011111", -- 2387 - 0x953  :   31 - 0x1f
    "00001100", -- 2388 - 0x954  :   12 - 0xc
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "00000000", -- 2391 - 0x957  :    0 - 0x0
    "00000000", -- 2392 - 0x958  :    0 - 0x0 -- Background 0x2b
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- Background 0x2d
    "01111110", -- 2409 - 0x969  :  126 - 0x7e
    "01000010", -- 2410 - 0x96a  :   66 - 0x42
    "01000010", -- 2411 - 0x96b  :   66 - 0x42
    "01000010", -- 2412 - 0x96c  :   66 - 0x42
    "01000010", -- 2413 - 0x96d  :   66 - 0x42
    "01111110", -- 2414 - 0x96e  :  126 - 0x7e
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "01100110", -- 2424 - 0x978  :  102 - 0x66 -- Background 0x2f
    "01100000", -- 2425 - 0x979  :   96 - 0x60
    "01101000", -- 2426 - 0x97a  :  104 - 0x68
    "11100000", -- 2427 - 0x97b  :  224 - 0xe0
    "11000000", -- 2428 - 0x97c  :  192 - 0xc0
    "00010000", -- 2429 - 0x97d  :   16 - 0x10
    "00101000", -- 2430 - 0x97e  :   40 - 0x28
    "01010000", -- 2431 - 0x97f  :   80 - 0x50
    "11110110", -- 2432 - 0x980  :  246 - 0xf6 -- Background 0x30
    "11110000", -- 2433 - 0x981  :  240 - 0xf0
    "00111000", -- 2434 - 0x982  :   56 - 0x38
    "11010000", -- 2435 - 0x983  :  208 - 0xd0
    "11000000", -- 2436 - 0x984  :  192 - 0xc0
    "11111000", -- 2437 - 0x985  :  248 - 0xf8
    "01111000", -- 2438 - 0x986  :  120 - 0x78
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "11110110", -- 2440 - 0x988  :  246 - 0xf6 -- Background 0x31
    "11110000", -- 2441 - 0x989  :  240 - 0xf0
    "00111000", -- 2442 - 0x98a  :   56 - 0x38
    "11010000", -- 2443 - 0x98b  :  208 - 0xd0
    "11000000", -- 2444 - 0x98c  :  192 - 0xc0
    "11100000", -- 2445 - 0x98d  :  224 - 0xe0
    "01111000", -- 2446 - 0x98e  :  120 - 0x78
    "00111000", -- 2447 - 0x98f  :   56 - 0x38
    "11110110", -- 2448 - 0x990  :  246 - 0xf6 -- Background 0x32
    "11110000", -- 2449 - 0x991  :  240 - 0xf0
    "00111000", -- 2450 - 0x992  :   56 - 0x38
    "11000000", -- 2451 - 0x993  :  192 - 0xc0
    "11011000", -- 2452 - 0x994  :  216 - 0xd8
    "11111000", -- 2453 - 0x995  :  248 - 0xf8
    "01100000", -- 2454 - 0x996  :   96 - 0x60
    "00010000", -- 2455 - 0x997  :   16 - 0x10
    "00011100", -- 2456 - 0x998  :   28 - 0x1c -- Background 0x33
    "00011100", -- 2457 - 0x999  :   28 - 0x1c
    "00011110", -- 2458 - 0x99a  :   30 - 0x1e
    "00011111", -- 2459 - 0x99b  :   31 - 0x1f
    "00001100", -- 2460 - 0x99c  :   12 - 0xc
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "10000000", -- 2464 - 0x9a0  :  128 - 0x80 -- Background 0x34
    "01010000", -- 2465 - 0x9a1  :   80 - 0x50
    "10101000", -- 2466 - 0x9a2  :  168 - 0xa8
    "00000000", -- 2467 - 0x9a3  :    0 - 0x0
    "01011000", -- 2468 - 0x9a4  :   88 - 0x58
    "11011000", -- 2469 - 0x9a5  :  216 - 0xd8
    "11101100", -- 2470 - 0x9a6  :  236 - 0xec
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00011100", -- 2472 - 0x9a8  :   28 - 0x1c -- Background 0x35
    "00011100", -- 2473 - 0x9a9  :   28 - 0x1c
    "00011110", -- 2474 - 0x9aa  :   30 - 0x1e
    "00011111", -- 2475 - 0x9ab  :   31 - 0x1f
    "00001100", -- 2476 - 0x9ac  :   12 - 0xc
    "00000001", -- 2477 - 0x9ad  :    1 - 0x1
    "00000001", -- 2478 - 0x9ae  :    1 - 0x1
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "10101000", -- 2480 - 0x9b0  :  168 - 0xa8 -- Background 0x36
    "01010000", -- 2481 - 0x9b1  :   80 - 0x50
    "10101000", -- 2482 - 0x9b2  :  168 - 0xa8
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "01011000", -- 2484 - 0x9b4  :   88 - 0x58
    "11001110", -- 2485 - 0x9b5  :  206 - 0xce
    "10000110", -- 2486 - 0x9b6  :  134 - 0x86
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "10101000", -- 2488 - 0x9b8  :  168 - 0xa8 -- Background 0x37
    "01010000", -- 2489 - 0x9b9  :   80 - 0x50
    "10101000", -- 2490 - 0x9ba  :  168 - 0xa8
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "01011000", -- 2492 - 0x9bc  :   88 - 0x58
    "11011000", -- 2493 - 0x9bd  :  216 - 0xd8
    "11101100", -- 2494 - 0x9be  :  236 - 0xec
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00111100", -- 2560 - 0xa00  :   60 - 0x3c -- Background 0x40
    "01111100", -- 2561 - 0xa01  :  124 - 0x7c
    "11100110", -- 2562 - 0xa02  :  230 - 0xe6
    "11101110", -- 2563 - 0xa03  :  238 - 0xee
    "11110110", -- 2564 - 0xa04  :  246 - 0xf6
    "11100110", -- 2565 - 0xa05  :  230 - 0xe6
    "00111100", -- 2566 - 0xa06  :   60 - 0x3c
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00111000", -- 2568 - 0xa08  :   56 - 0x38 -- Background 0x41
    "01111000", -- 2569 - 0xa09  :  120 - 0x78
    "00111000", -- 2570 - 0xa0a  :   56 - 0x38
    "00111000", -- 2571 - 0xa0b  :   56 - 0x38
    "00111000", -- 2572 - 0xa0c  :   56 - 0x38
    "00111000", -- 2573 - 0xa0d  :   56 - 0x38
    "00111000", -- 2574 - 0xa0e  :   56 - 0x38
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "01111100", -- 2576 - 0xa10  :  124 - 0x7c -- Background 0x42
    "11111110", -- 2577 - 0xa11  :  254 - 0xfe
    "11100110", -- 2578 - 0xa12  :  230 - 0xe6
    "00011110", -- 2579 - 0xa13  :   30 - 0x1e
    "01111100", -- 2580 - 0xa14  :  124 - 0x7c
    "11100000", -- 2581 - 0xa15  :  224 - 0xe0
    "11111110", -- 2582 - 0xa16  :  254 - 0xfe
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "01111100", -- 2584 - 0xa18  :  124 - 0x7c -- Background 0x43
    "11111100", -- 2585 - 0xa19  :  252 - 0xfc
    "11100110", -- 2586 - 0xa1a  :  230 - 0xe6
    "00011100", -- 2587 - 0xa1b  :   28 - 0x1c
    "01100110", -- 2588 - 0xa1c  :  102 - 0x66
    "11101110", -- 2589 - 0xa1d  :  238 - 0xee
    "11111100", -- 2590 - 0xa1e  :  252 - 0xfc
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00001100", -- 2592 - 0xa20  :   12 - 0xc -- Background 0x44
    "00011100", -- 2593 - 0xa21  :   28 - 0x1c
    "00111100", -- 2594 - 0xa22  :   60 - 0x3c
    "01111100", -- 2595 - 0xa23  :  124 - 0x7c
    "11101100", -- 2596 - 0xa24  :  236 - 0xec
    "11111110", -- 2597 - 0xa25  :  254 - 0xfe
    "00001100", -- 2598 - 0xa26  :   12 - 0xc
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "11111110", -- 2600 - 0xa28  :  254 - 0xfe -- Background 0x45
    "11111110", -- 2601 - 0xa29  :  254 - 0xfe
    "11100000", -- 2602 - 0xa2a  :  224 - 0xe0
    "11111110", -- 2603 - 0xa2b  :  254 - 0xfe
    "00000110", -- 2604 - 0xa2c  :    6 - 0x6
    "11101110", -- 2605 - 0xa2d  :  238 - 0xee
    "11111100", -- 2606 - 0xa2e  :  252 - 0xfc
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00111100", -- 2608 - 0xa30  :   60 - 0x3c -- Background 0x46
    "01111100", -- 2609 - 0xa31  :  124 - 0x7c
    "11100000", -- 2610 - 0xa32  :  224 - 0xe0
    "11111110", -- 2611 - 0xa33  :  254 - 0xfe
    "11100110", -- 2612 - 0xa34  :  230 - 0xe6
    "11101110", -- 2613 - 0xa35  :  238 - 0xee
    "00111100", -- 2614 - 0xa36  :   60 - 0x3c
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "11111110", -- 2616 - 0xa38  :  254 - 0xfe -- Background 0x47
    "11111100", -- 2617 - 0xa39  :  252 - 0xfc
    "00001100", -- 2618 - 0xa3a  :   12 - 0xc
    "00111000", -- 2619 - 0xa3b  :   56 - 0x38
    "00111000", -- 2620 - 0xa3c  :   56 - 0x38
    "01110000", -- 2621 - 0xa3d  :  112 - 0x70
    "01110000", -- 2622 - 0xa3e  :  112 - 0x70
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00111110", -- 2624 - 0xa40  :   62 - 0x3e -- Background 0x48
    "01111100", -- 2625 - 0xa41  :  124 - 0x7c
    "11100110", -- 2626 - 0xa42  :  230 - 0xe6
    "10111100", -- 2627 - 0xa43  :  188 - 0xbc
    "11100110", -- 2628 - 0xa44  :  230 - 0xe6
    "11101110", -- 2629 - 0xa45  :  238 - 0xee
    "00111100", -- 2630 - 0xa46  :   60 - 0x3c
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00111100", -- 2632 - 0xa48  :   60 - 0x3c -- Background 0x49
    "01111100", -- 2633 - 0xa49  :  124 - 0x7c
    "11100110", -- 2634 - 0xa4a  :  230 - 0xe6
    "11101110", -- 2635 - 0xa4b  :  238 - 0xee
    "11111110", -- 2636 - 0xa4c  :  254 - 0xfe
    "10000110", -- 2637 - 0xa4d  :  134 - 0x86
    "01111100", -- 2638 - 0xa4e  :  124 - 0x7c
    "01000000", -- 2639 - 0xa4f  :   64 - 0x40
    "11101110", -- 2640 - 0xa50  :  238 - 0xee -- Background 0x4a
    "11101110", -- 2641 - 0xa51  :  238 - 0xee
    "11101110", -- 2642 - 0xa52  :  238 - 0xee
    "11101110", -- 2643 - 0xa53  :  238 - 0xee
    "11101110", -- 2644 - 0xa54  :  238 - 0xee
    "11101110", -- 2645 - 0xa55  :  238 - 0xee
    "11101110", -- 2646 - 0xa56  :  238 - 0xee
    "10001000", -- 2647 - 0xa57  :  136 - 0x88
    "11100000", -- 2648 - 0xa58  :  224 - 0xe0 -- Background 0x4b
    "11100000", -- 2649 - 0xa59  :  224 - 0xe0
    "11100000", -- 2650 - 0xa5a  :  224 - 0xe0
    "11100000", -- 2651 - 0xa5b  :  224 - 0xe0
    "11100000", -- 2652 - 0xa5c  :  224 - 0xe0
    "11100000", -- 2653 - 0xa5d  :  224 - 0xe0
    "11100000", -- 2654 - 0xa5e  :  224 - 0xe0
    "10000000", -- 2655 - 0xa5f  :  128 - 0x80
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0x4c
    "01111111", -- 2657 - 0xa61  :  127 - 0x7f
    "01111111", -- 2658 - 0xa62  :  127 - 0x7f
    "01111111", -- 2659 - 0xa63  :  127 - 0x7f
    "01111111", -- 2660 - 0xa64  :  127 - 0x7f
    "01111111", -- 2661 - 0xa65  :  127 - 0x7f
    "01111111", -- 2662 - 0xa66  :  127 - 0x7f
    "01111111", -- 2663 - 0xa67  :  127 - 0x7f
    "01111111", -- 2664 - 0xa68  :  127 - 0x7f -- Background 0x4d
    "01111111", -- 2665 - 0xa69  :  127 - 0x7f
    "01111111", -- 2666 - 0xa6a  :  127 - 0x7f
    "01111111", -- 2667 - 0xa6b  :  127 - 0x7f
    "01111111", -- 2668 - 0xa6c  :  127 - 0x7f
    "01111111", -- 2669 - 0xa6d  :  127 - 0x7f
    "01111111", -- 2670 - 0xa6e  :  127 - 0x7f
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0 -- Background 0x4e
    "11111110", -- 2673 - 0xa71  :  254 - 0xfe
    "11111110", -- 2674 - 0xa72  :  254 - 0xfe
    "11111110", -- 2675 - 0xa73  :  254 - 0xfe
    "11111110", -- 2676 - 0xa74  :  254 - 0xfe
    "11111110", -- 2677 - 0xa75  :  254 - 0xfe
    "11111110", -- 2678 - 0xa76  :  254 - 0xfe
    "11111110", -- 2679 - 0xa77  :  254 - 0xfe
    "11111110", -- 2680 - 0xa78  :  254 - 0xfe -- Background 0x4f
    "11111110", -- 2681 - 0xa79  :  254 - 0xfe
    "11111110", -- 2682 - 0xa7a  :  254 - 0xfe
    "11111110", -- 2683 - 0xa7b  :  254 - 0xfe
    "11111110", -- 2684 - 0xa7c  :  254 - 0xfe
    "11111110", -- 2685 - 0xa7d  :  254 - 0xfe
    "11111110", -- 2686 - 0xa7e  :  254 - 0xfe
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Background 0x50
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00000000", -- 2693 - 0xa85  :    0 - 0x0
    "00000000", -- 2694 - 0xa86  :    0 - 0x0
    "00000000", -- 2695 - 0xa87  :    0 - 0x0
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- Background 0x51
    "00010000", -- 2697 - 0xa89  :   16 - 0x10
    "00010000", -- 2698 - 0xa8a  :   16 - 0x10
    "01111100", -- 2699 - 0xa8b  :  124 - 0x7c
    "00111000", -- 2700 - 0xa8c  :   56 - 0x38
    "00111000", -- 2701 - 0xa8d  :   56 - 0x38
    "01101100", -- 2702 - 0xa8e  :  108 - 0x6c
    "00000000", -- 2703 - 0xa8f  :    0 - 0x0
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00010000", -- 2705 - 0xa91  :   16 - 0x10
    "00010000", -- 2706 - 0xa92  :   16 - 0x10
    "01111100", -- 2707 - 0xa93  :  124 - 0x7c
    "00111000", -- 2708 - 0xa94  :   56 - 0x38
    "00111000", -- 2709 - 0xa95  :   56 - 0x38
    "01101100", -- 2710 - 0xa96  :  108 - 0x6c
    "00000000", -- 2711 - 0xa97  :    0 - 0x0
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- Background 0x53
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "11111111", -- 2720 - 0xaa0  :  255 - 0xff -- Background 0x54
    "11111111", -- 2721 - 0xaa1  :  255 - 0xff
    "11111111", -- 2722 - 0xaa2  :  255 - 0xff
    "11111111", -- 2723 - 0xaa3  :  255 - 0xff
    "11111111", -- 2724 - 0xaa4  :  255 - 0xff
    "11111111", -- 2725 - 0xaa5  :  255 - 0xff
    "11111111", -- 2726 - 0xaa6  :  255 - 0xff
    "11111111", -- 2727 - 0xaa7  :  255 - 0xff
    "11111111", -- 2728 - 0xaa8  :  255 - 0xff -- Background 0x55
    "11111111", -- 2729 - 0xaa9  :  255 - 0xff
    "11111111", -- 2730 - 0xaaa  :  255 - 0xff
    "11111111", -- 2731 - 0xaab  :  255 - 0xff
    "11111111", -- 2732 - 0xaac  :  255 - 0xff
    "11111111", -- 2733 - 0xaad  :  255 - 0xff
    "11111111", -- 2734 - 0xaae  :  255 - 0xff
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "00000010", -- 2736 - 0xab0  :    2 - 0x2 -- Background 0x56
    "00000101", -- 2737 - 0xab1  :    5 - 0x5
    "10101010", -- 2738 - 0xab2  :  170 - 0xaa
    "01010001", -- 2739 - 0xab3  :   81 - 0x51
    "10101010", -- 2740 - 0xab4  :  170 - 0xaa
    "01010001", -- 2741 - 0xab5  :   81 - 0x51
    "10100010", -- 2742 - 0xab6  :  162 - 0xa2
    "00000100", -- 2743 - 0xab7  :    4 - 0x4
    "00001000", -- 2744 - 0xab8  :    8 - 0x8 -- Background 0x57
    "01010101", -- 2745 - 0xab9  :   85 - 0x55
    "00101010", -- 2746 - 0xaba  :   42 - 0x2a
    "01010101", -- 2747 - 0xabb  :   85 - 0x55
    "00101010", -- 2748 - 0xabc  :   42 - 0x2a
    "01000101", -- 2749 - 0xabd  :   69 - 0x45
    "00001010", -- 2750 - 0xabe  :   10 - 0xa
    "00010000", -- 2751 - 0xabf  :   16 - 0x10
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Background 0x58
    "00111111", -- 2753 - 0xac1  :   63 - 0x3f
    "01011111", -- 2754 - 0xac2  :   95 - 0x5f
    "01101111", -- 2755 - 0xac3  :  111 - 0x6f
    "01110000", -- 2756 - 0xac4  :  112 - 0x70
    "01110111", -- 2757 - 0xac5  :  119 - 0x77
    "01110111", -- 2758 - 0xac6  :  119 - 0x77
    "01110111", -- 2759 - 0xac7  :  119 - 0x77
    "01110111", -- 2760 - 0xac8  :  119 - 0x77 -- Background 0x59
    "01110111", -- 2761 - 0xac9  :  119 - 0x77
    "01110111", -- 2762 - 0xaca  :  119 - 0x77
    "01110000", -- 2763 - 0xacb  :  112 - 0x70
    "01101111", -- 2764 - 0xacc  :  111 - 0x6f
    "01011111", -- 2765 - 0xacd  :   95 - 0x5f
    "00010101", -- 2766 - 0xace  :   21 - 0x15
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Background 0x5a
    "11111100", -- 2769 - 0xad1  :  252 - 0xfc
    "11111000", -- 2770 - 0xad2  :  248 - 0xf8
    "11110110", -- 2771 - 0xad3  :  246 - 0xf6
    "00001100", -- 2772 - 0xad4  :   12 - 0xc
    "11101110", -- 2773 - 0xad5  :  238 - 0xee
    "11101100", -- 2774 - 0xad6  :  236 - 0xec
    "11101110", -- 2775 - 0xad7  :  238 - 0xee
    "11101100", -- 2776 - 0xad8  :  236 - 0xec -- Background 0x5b
    "11101110", -- 2777 - 0xad9  :  238 - 0xee
    "11101100", -- 2778 - 0xada  :  236 - 0xec
    "00001110", -- 2779 - 0xadb  :   14 - 0xe
    "11110100", -- 2780 - 0xadc  :  244 - 0xf4
    "11111010", -- 2781 - 0xadd  :  250 - 0xfa
    "01010100", -- 2782 - 0xade  :   84 - 0x54
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Background 0x5c
    "00011100", -- 2785 - 0xae1  :   28 - 0x1c
    "00111110", -- 2786 - 0xae2  :   62 - 0x3e
    "00111110", -- 2787 - 0xae3  :   62 - 0x3e
    "00111110", -- 2788 - 0xae4  :   62 - 0x3e
    "00011100", -- 2789 - 0xae5  :   28 - 0x1c
    "00011100", -- 2790 - 0xae6  :   28 - 0x1c
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0x5e
    "00010100", -- 2801 - 0xaf1  :   20 - 0x14
    "00110110", -- 2802 - 0xaf2  :   54 - 0x36
    "00111110", -- 2803 - 0xaf3  :   62 - 0x3e
    "00111110", -- 2804 - 0xaf4  :   62 - 0x3e
    "00011100", -- 2805 - 0xaf5  :   28 - 0x1c
    "00001000", -- 2806 - 0xaf6  :    8 - 0x8
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- Background 0x5f
    "00010100", -- 2809 - 0xaf9  :   20 - 0x14
    "00011100", -- 2810 - 0xafa  :   28 - 0x1c
    "00011100", -- 2811 - 0xafb  :   28 - 0x1c
    "00011100", -- 2812 - 0xafc  :   28 - 0x1c
    "00011100", -- 2813 - 0xafd  :   28 - 0x1c
    "00011100", -- 2814 - 0xafe  :   28 - 0x1c
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Background 0x60
    "01111111", -- 2817 - 0xb01  :  127 - 0x7f
    "01111111", -- 2818 - 0xb02  :  127 - 0x7f
    "01111111", -- 2819 - 0xb03  :  127 - 0x7f
    "01111111", -- 2820 - 0xb04  :  127 - 0x7f
    "01111111", -- 2821 - 0xb05  :  127 - 0x7f
    "00101010", -- 2822 - 0xb06  :   42 - 0x2a
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- Background 0x61
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11111111", -- 2826 - 0xb0a  :  255 - 0xff
    "11111111", -- 2827 - 0xb0b  :  255 - 0xff
    "11111111", -- 2828 - 0xb0c  :  255 - 0xff
    "11111111", -- 2829 - 0xb0d  :  255 - 0xff
    "10101010", -- 2830 - 0xb0e  :  170 - 0xaa
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Background 0x62
    "11111110", -- 2833 - 0xb11  :  254 - 0xfe
    "11111110", -- 2834 - 0xb12  :  254 - 0xfe
    "11111110", -- 2835 - 0xb13  :  254 - 0xfe
    "11111110", -- 2836 - 0xb14  :  254 - 0xfe
    "11111110", -- 2837 - 0xb15  :  254 - 0xfe
    "10101010", -- 2838 - 0xb16  :  170 - 0xaa
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00000000", -- 2840 - 0xb18  :    0 - 0x0 -- Background 0x63
    "00000000", -- 2841 - 0xb19  :    0 - 0x0
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "00000000", -- 2845 - 0xb1d  :    0 - 0x0
    "00000000", -- 2846 - 0xb1e  :    0 - 0x0
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0x64
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000001", -- 2850 - 0xb22  :    1 - 0x1
    "00000001", -- 2851 - 0xb23  :    1 - 0x1
    "00000011", -- 2852 - 0xb24  :    3 - 0x3
    "00000011", -- 2853 - 0xb25  :    3 - 0x3
    "00000111", -- 2854 - 0xb26  :    7 - 0x7
    "00000111", -- 2855 - 0xb27  :    7 - 0x7
    "00001111", -- 2856 - 0xb28  :   15 - 0xf -- Background 0x65
    "00001111", -- 2857 - 0xb29  :   15 - 0xf
    "00011111", -- 2858 - 0xb2a  :   31 - 0x1f
    "00011111", -- 2859 - 0xb2b  :   31 - 0x1f
    "00111111", -- 2860 - 0xb2c  :   63 - 0x3f
    "00111111", -- 2861 - 0xb2d  :   63 - 0x3f
    "01010101", -- 2862 - 0xb2e  :   85 - 0x55
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00000000", -- 2864 - 0xb30  :    0 - 0x0 -- Background 0x66
    "00000000", -- 2865 - 0xb31  :    0 - 0x0
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "10000000", -- 2867 - 0xb33  :  128 - 0x80
    "01000000", -- 2868 - 0xb34  :   64 - 0x40
    "10000000", -- 2869 - 0xb35  :  128 - 0x80
    "11000000", -- 2870 - 0xb36  :  192 - 0xc0
    "11100000", -- 2871 - 0xb37  :  224 - 0xe0
    "11010000", -- 2872 - 0xb38  :  208 - 0xd0 -- Background 0x67
    "11100000", -- 2873 - 0xb39  :  224 - 0xe0
    "11110000", -- 2874 - 0xb3a  :  240 - 0xf0
    "11101000", -- 2875 - 0xb3b  :  232 - 0xe8
    "11110100", -- 2876 - 0xb3c  :  244 - 0xf4
    "11111000", -- 2877 - 0xb3d  :  248 - 0xf8
    "01010100", -- 2878 - 0xb3e  :   84 - 0x54
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Background 0x68
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000000", -- 2883 - 0xb43  :    0 - 0x0
    "00000000", -- 2884 - 0xb44  :    0 - 0x0
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- Background 0x69
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00000000", -- 2890 - 0xb4a  :    0 - 0x0
    "00000000", -- 2891 - 0xb4b  :    0 - 0x0
    "00000000", -- 2892 - 0xb4c  :    0 - 0x0
    "00000000", -- 2893 - 0xb4d  :    0 - 0x0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00000000", -- 2904 - 0xb58  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "00000000", -- 2906 - 0xb5a  :    0 - 0x0
    "00000000", -- 2907 - 0xb5b  :    0 - 0x0
    "00000000", -- 2908 - 0xb5c  :    0 - 0x0
    "00000000", -- 2909 - 0xb5d  :    0 - 0x0
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "00000000", -- 2915 - 0xb63  :    0 - 0x0
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00000000", -- 2936 - 0xb78  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 2937 - 0xb79  :    0 - 0x0
    "00000000", -- 2938 - 0xb7a  :    0 - 0x0
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0x70
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000000", -- 2946 - 0xb82  :    0 - 0x0
    "00000000", -- 2947 - 0xb83  :    0 - 0x0
    "00000000", -- 2948 - 0xb84  :    0 - 0x0
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- Background 0x71
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "00000000", -- 2957 - 0xb8d  :    0 - 0x0
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Background 0x72
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "00000000", -- 2962 - 0xb92  :    0 - 0x0
    "00000000", -- 2963 - 0xb93  :    0 - 0x0
    "00000000", -- 2964 - 0xb94  :    0 - 0x0
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- Background 0x73
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Background 0x74
    "00000000", -- 2977 - 0xba1  :    0 - 0x0
    "00000000", -- 2978 - 0xba2  :    0 - 0x0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00000000", -- 2980 - 0xba4  :    0 - 0x0
    "00000000", -- 2981 - 0xba5  :    0 - 0x0
    "00000000", -- 2982 - 0xba6  :    0 - 0x0
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- Background 0x75
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000000", -- 2992 - 0xbb0  :    0 - 0x0 -- Background 0x76
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0 -- Background 0x77
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- Background 0x79
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Background 0x7c
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "00000000", -- 3042 - 0xbe2  :    0 - 0x0
    "00000000", -- 3043 - 0xbe3  :    0 - 0x0
    "00000000", -- 3044 - 0xbe4  :    0 - 0x0
    "00000000", -- 3045 - 0xbe5  :    0 - 0x0
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0x80
    "00000011", -- 3073 - 0xc01  :    3 - 0x3
    "00001111", -- 3074 - 0xc02  :   15 - 0xf
    "00011111", -- 3075 - 0xc03  :   31 - 0x1f
    "00011111", -- 3076 - 0xc04  :   31 - 0x1f
    "00111111", -- 3077 - 0xc05  :   63 - 0x3f
    "00111111", -- 3078 - 0xc06  :   63 - 0x3f
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- Background 0x81
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Background 0x82
    "11000000", -- 3089 - 0xc11  :  192 - 0xc0
    "11110000", -- 3090 - 0xc12  :  240 - 0xf0
    "11110000", -- 3091 - 0xc13  :  240 - 0xf0
    "11101100", -- 3092 - 0xc14  :  236 - 0xec
    "11100000", -- 3093 - 0xc15  :  224 - 0xe0
    "11111100", -- 3094 - 0xc16  :  252 - 0xfc
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0 -- Background 0x83
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "11100000", -- 3102 - 0xc1e  :  224 - 0xe0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0x84
    "00000011", -- 3105 - 0xc21  :    3 - 0x3
    "00001111", -- 3106 - 0xc22  :   15 - 0xf
    "00011111", -- 3107 - 0xc23  :   31 - 0x1f
    "00011111", -- 3108 - 0xc24  :   31 - 0x1f
    "00111111", -- 3109 - 0xc25  :   63 - 0x3f
    "00111111", -- 3110 - 0xc26  :   63 - 0x3f
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- Background 0x85
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00001000", -- 3117 - 0xc2d  :    8 - 0x8
    "00001110", -- 3118 - 0xc2e  :   14 - 0xe
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0x86
    "11000000", -- 3121 - 0xc31  :  192 - 0xc0
    "11110000", -- 3122 - 0xc32  :  240 - 0xf0
    "11110000", -- 3123 - 0xc33  :  240 - 0xf0
    "11101100", -- 3124 - 0xc34  :  236 - 0xec
    "11100000", -- 3125 - 0xc35  :  224 - 0xe0
    "11111100", -- 3126 - 0xc36  :  252 - 0xfc
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- Background 0x87
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000110", -- 3133 - 0xc3d  :    6 - 0x6
    "00001100", -- 3134 - 0xc3e  :   12 - 0xc
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0x88
    "00000011", -- 3137 - 0xc41  :    3 - 0x3
    "00000011", -- 3138 - 0xc42  :    3 - 0x3
    "00000100", -- 3139 - 0xc43  :    4 - 0x4
    "00001111", -- 3140 - 0xc44  :   15 - 0xf
    "00011111", -- 3141 - 0xc45  :   31 - 0x1f
    "01101111", -- 3142 - 0xc46  :  111 - 0x6f
    "01101111", -- 3143 - 0xc47  :  111 - 0x6f
    "01101111", -- 3144 - 0xc48  :  111 - 0x6f -- Background 0x89
    "01101111", -- 3145 - 0xc49  :  111 - 0x6f
    "00011111", -- 3146 - 0xc4a  :   31 - 0x1f
    "00001111", -- 3147 - 0xc4b  :   15 - 0xf
    "00000100", -- 3148 - 0xc4c  :    4 - 0x4
    "00000011", -- 3149 - 0xc4d  :    3 - 0x3
    "00000011", -- 3150 - 0xc4e  :    3 - 0x3
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00011000", -- 3154 - 0xc52  :   24 - 0x18
    "00110111", -- 3155 - 0xc53  :   55 - 0x37
    "00101111", -- 3156 - 0xc54  :   47 - 0x2f
    "00011111", -- 3157 - 0xc55  :   31 - 0x1f
    "00011111", -- 3158 - 0xc56  :   31 - 0x1f
    "00011111", -- 3159 - 0xc57  :   31 - 0x1f
    "00011111", -- 3160 - 0xc58  :   31 - 0x1f -- Background 0x8b
    "00011111", -- 3161 - 0xc59  :   31 - 0x1f
    "00011111", -- 3162 - 0xc5a  :   31 - 0x1f
    "00101111", -- 3163 - 0xc5b  :   47 - 0x2f
    "00110111", -- 3164 - 0xc5c  :   55 - 0x37
    "00011000", -- 3165 - 0xc5d  :   24 - 0x18
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Background 0x8c
    "00000011", -- 3169 - 0xc61  :    3 - 0x3
    "00000001", -- 3170 - 0xc62  :    1 - 0x1
    "00011001", -- 3171 - 0xc63  :   25 - 0x19
    "00111001", -- 3172 - 0xc64  :   57 - 0x39
    "00011011", -- 3173 - 0xc65  :   27 - 0x1b
    "00001111", -- 3174 - 0xc66  :   15 - 0xf
    "00001111", -- 3175 - 0xc67  :   15 - 0xf
    "01111111", -- 3176 - 0xc68  :  127 - 0x7f -- Background 0x8d
    "01111111", -- 3177 - 0xc69  :  127 - 0x7f
    "00111111", -- 3178 - 0xc6a  :   63 - 0x3f
    "00010111", -- 3179 - 0xc6b  :   23 - 0x17
    "00000110", -- 3180 - 0xc6c  :    6 - 0x6
    "00000100", -- 3181 - 0xc6d  :    4 - 0x4
    "00000111", -- 3182 - 0xc6e  :    7 - 0x7
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000000", -- 3184 - 0xc70  :    0 - 0x0 -- Background 0x8e
    "11000000", -- 3185 - 0xc71  :  192 - 0xc0
    "11110000", -- 3186 - 0xc72  :  240 - 0xf0
    "10111000", -- 3187 - 0xc73  :  184 - 0xb8
    "10011100", -- 3188 - 0xc74  :  156 - 0x9c
    "11111100", -- 3189 - 0xc75  :  252 - 0xfc
    "11111110", -- 3190 - 0xc76  :  254 - 0xfe
    "11000000", -- 3191 - 0xc77  :  192 - 0xc0
    "11111110", -- 3192 - 0xc78  :  254 - 0xfe -- Background 0x8f
    "11111110", -- 3193 - 0xc79  :  254 - 0xfe
    "11111000", -- 3194 - 0xc7a  :  248 - 0xf8
    "11110000", -- 3195 - 0xc7b  :  240 - 0xf0
    "11000000", -- 3196 - 0xc7c  :  192 - 0xc0
    "00000000", -- 3197 - 0xc7d  :    0 - 0x0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "10000000", -- 3199 - 0xc7f  :  128 - 0x80
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000001", -- 3201 - 0xc81  :    1 - 0x1
    "00001001", -- 3202 - 0xc82  :    9 - 0x9
    "00011001", -- 3203 - 0xc83  :   25 - 0x19
    "00011100", -- 3204 - 0xc84  :   28 - 0x1c
    "00001101", -- 3205 - 0xc85  :   13 - 0xd
    "00001111", -- 3206 - 0xc86  :   15 - 0xf
    "00101111", -- 3207 - 0xc87  :   47 - 0x2f
    "01111111", -- 3208 - 0xc88  :  127 - 0x7f -- Background 0x91
    "01111111", -- 3209 - 0xc89  :  127 - 0x7f
    "00111111", -- 3210 - 0xc8a  :   63 - 0x3f
    "00011011", -- 3211 - 0xc8b  :   27 - 0x1b
    "00000011", -- 3212 - 0xc8c  :    3 - 0x3
    "00000011", -- 3213 - 0xc8d  :    3 - 0x3
    "00000001", -- 3214 - 0xc8e  :    1 - 0x1
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0 -- Background 0x92
    "11000000", -- 3217 - 0xc91  :  192 - 0xc0
    "11110000", -- 3218 - 0xc92  :  240 - 0xf0
    "11011000", -- 3219 - 0xc93  :  216 - 0xd8
    "11001100", -- 3220 - 0xc94  :  204 - 0xcc
    "11111100", -- 3221 - 0xc95  :  252 - 0xfc
    "11111110", -- 3222 - 0xc96  :  254 - 0xfe
    "11100000", -- 3223 - 0xc97  :  224 - 0xe0
    "11111110", -- 3224 - 0xc98  :  254 - 0xfe -- Background 0x93
    "11111110", -- 3225 - 0xc99  :  254 - 0xfe
    "11111000", -- 3226 - 0xc9a  :  248 - 0xf8
    "01110000", -- 3227 - 0xc9b  :  112 - 0x70
    "01000000", -- 3228 - 0xc9c  :   64 - 0x40
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "11000000", -- 3230 - 0xc9e  :  192 - 0xc0
    "00100000", -- 3231 - 0xc9f  :   32 - 0x20
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00001100", -- 3234 - 0xca2  :   12 - 0xc
    "00001110", -- 3235 - 0xca3  :   14 - 0xe
    "00000110", -- 3236 - 0xca4  :    6 - 0x6
    "00100110", -- 3237 - 0xca5  :   38 - 0x26
    "00110111", -- 3238 - 0xca6  :   55 - 0x37
    "00110011", -- 3239 - 0xca7  :   51 - 0x33
    "01111111", -- 3240 - 0xca8  :  127 - 0x7f -- Background 0x95
    "01111111", -- 3241 - 0xca9  :  127 - 0x7f
    "00111111", -- 3242 - 0xcaa  :   63 - 0x3f
    "00011111", -- 3243 - 0xcab  :   31 - 0x1f
    "00001110", -- 3244 - 0xcac  :   14 - 0xe
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Background 0x96
    "11000000", -- 3249 - 0xcb1  :  192 - 0xc0
    "11110000", -- 3250 - 0xcb2  :  240 - 0xf0
    "01101000", -- 3251 - 0xcb3  :  104 - 0x68
    "01100100", -- 3252 - 0xcb4  :  100 - 0x64
    "11111100", -- 3253 - 0xcb5  :  252 - 0xfc
    "11111110", -- 3254 - 0xcb6  :  254 - 0xfe
    "11110000", -- 3255 - 0xcb7  :  240 - 0xf0
    "11111111", -- 3256 - 0xcb8  :  255 - 0xff -- Background 0x97
    "11111110", -- 3257 - 0xcb9  :  254 - 0xfe
    "11111100", -- 3258 - 0xcba  :  252 - 0xfc
    "10110000", -- 3259 - 0xcbb  :  176 - 0xb0
    "11000000", -- 3260 - 0xcbc  :  192 - 0xc0
    "11000000", -- 3261 - 0xcbd  :  192 - 0xc0
    "01110000", -- 3262 - 0xcbe  :  112 - 0x70
    "00001000", -- 3263 - 0xcbf  :    8 - 0x8
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Background 0x98
    "00000001", -- 3265 - 0xcc1  :    1 - 0x1
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000001", -- 3270 - 0xcc6  :    1 - 0x1
    "00000011", -- 3271 - 0xcc7  :    3 - 0x3
    "00000111", -- 3272 - 0xcc8  :    7 - 0x7 -- Background 0x99
    "00010111", -- 3273 - 0xcc9  :   23 - 0x17
    "00101111", -- 3274 - 0xcca  :   47 - 0x2f
    "00011110", -- 3275 - 0xccb  :   30 - 0x1e
    "00010001", -- 3276 - 0xccc  :   17 - 0x11
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000001", -- 3278 - 0xcce  :    1 - 0x1
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0x9a
    "00010000", -- 3281 - 0xcd1  :   16 - 0x10
    "01111000", -- 3282 - 0xcd2  :  120 - 0x78
    "01110100", -- 3283 - 0xcd3  :  116 - 0x74
    "11111110", -- 3284 - 0xcd4  :  254 - 0xfe
    "11111000", -- 3285 - 0xcd5  :  248 - 0xf8
    "11111100", -- 3286 - 0xcd6  :  252 - 0xfc
    "11111000", -- 3287 - 0xcd7  :  248 - 0xf8
    "11111000", -- 3288 - 0xcd8  :  248 - 0xf8 -- Background 0x9b
    "11010000", -- 3289 - 0xcd9  :  208 - 0xd0
    "00110000", -- 3290 - 0xcda  :   48 - 0x30
    "01100000", -- 3291 - 0xcdb  :   96 - 0x60
    "10000000", -- 3292 - 0xcdc  :  128 - 0x80
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0x9c
    "00000001", -- 3297 - 0xce1  :    1 - 0x1
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000001", -- 3302 - 0xce6  :    1 - 0x1
    "00000011", -- 3303 - 0xce7  :    3 - 0x3
    "00000111", -- 3304 - 0xce8  :    7 - 0x7 -- Background 0x9d
    "00010111", -- 3305 - 0xce9  :   23 - 0x17
    "00101111", -- 3306 - 0xcea  :   47 - 0x2f
    "00011110", -- 3307 - 0xceb  :   30 - 0x1e
    "00010000", -- 3308 - 0xcec  :   16 - 0x10
    "00000100", -- 3309 - 0xced  :    4 - 0x4
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Background 0x9e
    "00010000", -- 3313 - 0xcf1  :   16 - 0x10
    "01111000", -- 3314 - 0xcf2  :  120 - 0x78
    "01110100", -- 3315 - 0xcf3  :  116 - 0x74
    "11111110", -- 3316 - 0xcf4  :  254 - 0xfe
    "11111000", -- 3317 - 0xcf5  :  248 - 0xf8
    "11111100", -- 3318 - 0xcf6  :  252 - 0xfc
    "11111000", -- 3319 - 0xcf7  :  248 - 0xf8
    "11111000", -- 3320 - 0xcf8  :  248 - 0xf8 -- Background 0x9f
    "11010000", -- 3321 - 0xcf9  :  208 - 0xd0
    "00110000", -- 3322 - 0xcfa  :   48 - 0x30
    "11000000", -- 3323 - 0xcfb  :  192 - 0xc0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Background 0xa0
    "00000011", -- 3329 - 0xd01  :    3 - 0x3
    "00001111", -- 3330 - 0xd02  :   15 - 0xf
    "00011111", -- 3331 - 0xd03  :   31 - 0x1f
    "00111111", -- 3332 - 0xd04  :   63 - 0x3f
    "00111111", -- 3333 - 0xd05  :   63 - 0x3f
    "01111111", -- 3334 - 0xd06  :  127 - 0x7f
    "01111111", -- 3335 - 0xd07  :  127 - 0x7f
    "01111111", -- 3336 - 0xd08  :  127 - 0x7f -- Background 0xa1
    "01111111", -- 3337 - 0xd09  :  127 - 0x7f
    "00111111", -- 3338 - 0xd0a  :   63 - 0x3f
    "00111111", -- 3339 - 0xd0b  :   63 - 0x3f
    "00011111", -- 3340 - 0xd0c  :   31 - 0x1f
    "00000101", -- 3341 - 0xd0d  :    5 - 0x5
    "00000010", -- 3342 - 0xd0e  :    2 - 0x2
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00000000", -- 3344 - 0xd10  :    0 - 0x0 -- Background 0xa2
    "11000000", -- 3345 - 0xd11  :  192 - 0xc0
    "11110000", -- 3346 - 0xd12  :  240 - 0xf0
    "11111000", -- 3347 - 0xd13  :  248 - 0xf8
    "11111000", -- 3348 - 0xd14  :  248 - 0xf8
    "11111100", -- 3349 - 0xd15  :  252 - 0xfc
    "11111010", -- 3350 - 0xd16  :  250 - 0xfa
    "11111100", -- 3351 - 0xd17  :  252 - 0xfc
    "11111010", -- 3352 - 0xd18  :  250 - 0xfa -- Background 0xa3
    "11110100", -- 3353 - 0xd19  :  244 - 0xf4
    "11101000", -- 3354 - 0xd1a  :  232 - 0xe8
    "11010100", -- 3355 - 0xd1b  :  212 - 0xd4
    "10101000", -- 3356 - 0xd1c  :  168 - 0xa8
    "01010000", -- 3357 - 0xd1d  :   80 - 0x50
    "10000000", -- 3358 - 0xd1e  :  128 - 0x80
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xa4
    "00000000", -- 3361 - 0xd21  :    0 - 0x0
    "00000000", -- 3362 - 0xd22  :    0 - 0x0
    "00001110", -- 3363 - 0xd23  :   14 - 0xe
    "00000000", -- 3364 - 0xd24  :    0 - 0x0
    "00001010", -- 3365 - 0xd25  :   10 - 0xa
    "01001010", -- 3366 - 0xd26  :   74 - 0x4a
    "01100000", -- 3367 - 0xd27  :   96 - 0x60
    "01111111", -- 3368 - 0xd28  :  127 - 0x7f -- Background 0xa5
    "01111000", -- 3369 - 0xd29  :  120 - 0x78
    "00110111", -- 3370 - 0xd2a  :   55 - 0x37
    "00111011", -- 3371 - 0xd2b  :   59 - 0x3b
    "00111100", -- 3372 - 0xd2c  :   60 - 0x3c
    "00011111", -- 3373 - 0xd2d  :   31 - 0x1f
    "00000111", -- 3374 - 0xd2e  :    7 - 0x7
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00000000", -- 3376 - 0xd30  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "00000000", -- 3378 - 0xd32  :    0 - 0x0
    "01110000", -- 3379 - 0xd33  :  112 - 0x70
    "00000000", -- 3380 - 0xd34  :    0 - 0x0
    "01010000", -- 3381 - 0xd35  :   80 - 0x50
    "01010010", -- 3382 - 0xd36  :   82 - 0x52
    "00000110", -- 3383 - 0xd37  :    6 - 0x6
    "11111100", -- 3384 - 0xd38  :  252 - 0xfc -- Background 0xa7
    "00011010", -- 3385 - 0xd39  :   26 - 0x1a
    "11101100", -- 3386 - 0xd3a  :  236 - 0xec
    "11011000", -- 3387 - 0xd3b  :  216 - 0xd8
    "00110100", -- 3388 - 0xd3c  :   52 - 0x34
    "11101000", -- 3389 - 0xd3d  :  232 - 0xe8
    "11000000", -- 3390 - 0xd3e  :  192 - 0xc0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xa8
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00001110", -- 3395 - 0xd43  :   14 - 0xe
    "00000000", -- 3396 - 0xd44  :    0 - 0x0
    "00001110", -- 3397 - 0xd45  :   14 - 0xe
    "01001010", -- 3398 - 0xd46  :   74 - 0x4a
    "01100000", -- 3399 - 0xd47  :   96 - 0x60
    "01111111", -- 3400 - 0xd48  :  127 - 0x7f -- Background 0xa9
    "01111100", -- 3401 - 0xd49  :  124 - 0x7c
    "01111011", -- 3402 - 0xd4a  :  123 - 0x7b
    "01110111", -- 3403 - 0xd4b  :  119 - 0x77
    "01111000", -- 3404 - 0xd4c  :  120 - 0x78
    "01111111", -- 3405 - 0xd4d  :  127 - 0x7f
    "01111111", -- 3406 - 0xd4e  :  127 - 0x7f
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Background 0xaa
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "01110000", -- 3411 - 0xd53  :  112 - 0x70
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "01110000", -- 3413 - 0xd55  :  112 - 0x70
    "01010010", -- 3414 - 0xd56  :   82 - 0x52
    "00000110", -- 3415 - 0xd57  :    6 - 0x6
    "11111100", -- 3416 - 0xd58  :  252 - 0xfc -- Background 0xab
    "00111010", -- 3417 - 0xd59  :   58 - 0x3a
    "11011100", -- 3418 - 0xd5a  :  220 - 0xdc
    "11101010", -- 3419 - 0xd5b  :  234 - 0xea
    "00011100", -- 3420 - 0xd5c  :   28 - 0x1c
    "11111010", -- 3421 - 0xd5d  :  250 - 0xfa
    "11110100", -- 3422 - 0xd5e  :  244 - 0xf4
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xac
    "00000011", -- 3425 - 0xd61  :    3 - 0x3
    "00001111", -- 3426 - 0xd62  :   15 - 0xf
    "00001111", -- 3427 - 0xd63  :   15 - 0xf
    "00011111", -- 3428 - 0xd64  :   31 - 0x1f
    "01011111", -- 3429 - 0xd65  :   95 - 0x5f
    "01010000", -- 3430 - 0xd66  :   80 - 0x50
    "00010000", -- 3431 - 0xd67  :   16 - 0x10
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- Background 0xad
    "11111010", -- 3433 - 0xd69  :  250 - 0xfa
    "11111010", -- 3434 - 0xd6a  :  250 - 0xfa
    "11111010", -- 3435 - 0xd6b  :  250 - 0xfa
    "10111010", -- 3436 - 0xd6c  :  186 - 0xba
    "10011010", -- 3437 - 0xd6d  :  154 - 0x9a
    "00001010", -- 3438 - 0xd6e  :   10 - 0xa
    "00000010", -- 3439 - 0xd6f  :    2 - 0x2
    "00000000", -- 3440 - 0xd70  :    0 - 0x0 -- Background 0xae
    "00000011", -- 3441 - 0xd71  :    3 - 0x3
    "00001111", -- 3442 - 0xd72  :   15 - 0xf
    "00001111", -- 3443 - 0xd73  :   15 - 0xf
    "00011111", -- 3444 - 0xd74  :   31 - 0x1f
    "01011111", -- 3445 - 0xd75  :   95 - 0x5f
    "01010000", -- 3446 - 0xd76  :   80 - 0x50
    "00010111", -- 3447 - 0xd77  :   23 - 0x17
    "00000000", -- 3448 - 0xd78  :    0 - 0x0 -- Background 0xaf
    "11111010", -- 3449 - 0xd79  :  250 - 0xfa
    "11111010", -- 3450 - 0xd7a  :  250 - 0xfa
    "11111010", -- 3451 - 0xd7b  :  250 - 0xfa
    "00111010", -- 3452 - 0xd7c  :   58 - 0x3a
    "01011010", -- 3453 - 0xd7d  :   90 - 0x5a
    "01101010", -- 3454 - 0xd7e  :  106 - 0x6a
    "11110010", -- 3455 - 0xd7f  :  242 - 0xf2
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000011", -- 3458 - 0xd82  :    3 - 0x3
    "00001111", -- 3459 - 0xd83  :   15 - 0xf
    "00111011", -- 3460 - 0xd84  :   59 - 0x3b
    "00111111", -- 3461 - 0xd85  :   63 - 0x3f
    "01101111", -- 3462 - 0xd86  :  111 - 0x6f
    "01111101", -- 3463 - 0xd87  :  125 - 0x7d
    "00001111", -- 3464 - 0xd88  :   15 - 0xf -- Background 0xb1
    "01110000", -- 3465 - 0xd89  :  112 - 0x70
    "01111111", -- 3466 - 0xd8a  :  127 - 0x7f
    "00001111", -- 3467 - 0xd8b  :   15 - 0xf
    "01110000", -- 3468 - 0xd8c  :  112 - 0x70
    "01111111", -- 3469 - 0xd8d  :  127 - 0x7f
    "00001111", -- 3470 - 0xd8e  :   15 - 0xf
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00000000", -- 3472 - 0xd90  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 3473 - 0xd91  :    0 - 0x0
    "11000000", -- 3474 - 0xd92  :  192 - 0xc0
    "11110000", -- 3475 - 0xd93  :  240 - 0xf0
    "10111100", -- 3476 - 0xd94  :  188 - 0xbc
    "11110100", -- 3477 - 0xd95  :  244 - 0xf4
    "11111110", -- 3478 - 0xd96  :  254 - 0xfe
    "11011110", -- 3479 - 0xd97  :  222 - 0xde
    "11110000", -- 3480 - 0xd98  :  240 - 0xf0 -- Background 0xb3
    "00001110", -- 3481 - 0xd99  :   14 - 0xe
    "11111110", -- 3482 - 0xd9a  :  254 - 0xfe
    "11110000", -- 3483 - 0xd9b  :  240 - 0xf0
    "00001110", -- 3484 - 0xd9c  :   14 - 0xe
    "11111110", -- 3485 - 0xd9d  :  254 - 0xfe
    "11110000", -- 3486 - 0xd9e  :  240 - 0xf0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Background 0xb4
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000011", -- 3490 - 0xda2  :    3 - 0x3
    "00001111", -- 3491 - 0xda3  :   15 - 0xf
    "00111011", -- 3492 - 0xda4  :   59 - 0x3b
    "00111111", -- 3493 - 0xda5  :   63 - 0x3f
    "01101111", -- 3494 - 0xda6  :  111 - 0x6f
    "01111101", -- 3495 - 0xda7  :  125 - 0x7d
    "00001111", -- 3496 - 0xda8  :   15 - 0xf -- Background 0xb5
    "01110000", -- 3497 - 0xda9  :  112 - 0x70
    "01111111", -- 3498 - 0xdaa  :  127 - 0x7f
    "00001111", -- 3499 - 0xdab  :   15 - 0xf
    "01110000", -- 3500 - 0xdac  :  112 - 0x70
    "01111111", -- 3501 - 0xdad  :  127 - 0x7f
    "00001111", -- 3502 - 0xdae  :   15 - 0xf
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 3505 - 0xdb1  :    0 - 0x0
    "11000000", -- 3506 - 0xdb2  :  192 - 0xc0
    "11110000", -- 3507 - 0xdb3  :  240 - 0xf0
    "10111100", -- 3508 - 0xdb4  :  188 - 0xbc
    "11110100", -- 3509 - 0xdb5  :  244 - 0xf4
    "11111110", -- 3510 - 0xdb6  :  254 - 0xfe
    "11011110", -- 3511 - 0xdb7  :  222 - 0xde
    "11110000", -- 3512 - 0xdb8  :  240 - 0xf0 -- Background 0xb7
    "00001110", -- 3513 - 0xdb9  :   14 - 0xe
    "11111110", -- 3514 - 0xdba  :  254 - 0xfe
    "11110000", -- 3515 - 0xdbb  :  240 - 0xf0
    "00001110", -- 3516 - 0xdbc  :   14 - 0xe
    "11111110", -- 3517 - 0xdbd  :  254 - 0xfe
    "11110000", -- 3518 - 0xdbe  :  240 - 0xf0
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000011", -- 3522 - 0xdc2  :    3 - 0x3
    "00001111", -- 3523 - 0xdc3  :   15 - 0xf
    "00111011", -- 3524 - 0xdc4  :   59 - 0x3b
    "00111111", -- 3525 - 0xdc5  :   63 - 0x3f
    "01101111", -- 3526 - 0xdc6  :  111 - 0x6f
    "01111101", -- 3527 - 0xdc7  :  125 - 0x7d
    "00001111", -- 3528 - 0xdc8  :   15 - 0xf -- Background 0xb9
    "00100000", -- 3529 - 0xdc9  :   32 - 0x20
    "01010101", -- 3530 - 0xdca  :   85 - 0x55
    "00001010", -- 3531 - 0xdcb  :   10 - 0xa
    "01110000", -- 3532 - 0xdcc  :  112 - 0x70
    "01111111", -- 3533 - 0xdcd  :  127 - 0x7f
    "00001111", -- 3534 - 0xdce  :   15 - 0xf
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Background 0xba
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "11000000", -- 3538 - 0xdd2  :  192 - 0xc0
    "11110000", -- 3539 - 0xdd3  :  240 - 0xf0
    "10111100", -- 3540 - 0xdd4  :  188 - 0xbc
    "11110100", -- 3541 - 0xdd5  :  244 - 0xf4
    "11111110", -- 3542 - 0xdd6  :  254 - 0xfe
    "11011110", -- 3543 - 0xdd7  :  222 - 0xde
    "11110000", -- 3544 - 0xdd8  :  240 - 0xf0 -- Background 0xbb
    "00001010", -- 3545 - 0xdd9  :   10 - 0xa
    "01010100", -- 3546 - 0xdda  :   84 - 0x54
    "10100000", -- 3547 - 0xddb  :  160 - 0xa0
    "00001110", -- 3548 - 0xddc  :   14 - 0xe
    "11111110", -- 3549 - 0xddd  :  254 - 0xfe
    "11110000", -- 3550 - 0xdde  :  240 - 0xf0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Background 0xbc
    "01110011", -- 3553 - 0xde1  :  115 - 0x73
    "01111011", -- 3554 - 0xde2  :  123 - 0x7b
    "01111111", -- 3555 - 0xde3  :  127 - 0x7f
    "00111111", -- 3556 - 0xde4  :   63 - 0x3f
    "00011100", -- 3557 - 0xde5  :   28 - 0x1c
    "01111011", -- 3558 - 0xde6  :  123 - 0x7b
    "01111011", -- 3559 - 0xde7  :  123 - 0x7b
    "01111011", -- 3560 - 0xde8  :  123 - 0x7b -- Background 0xbd
    "01111011", -- 3561 - 0xde9  :  123 - 0x7b
    "00011100", -- 3562 - 0xdea  :   28 - 0x1c
    "00111111", -- 3563 - 0xdeb  :   63 - 0x3f
    "01111111", -- 3564 - 0xdec  :  127 - 0x7f
    "01111011", -- 3565 - 0xded  :  123 - 0x7b
    "01110011", -- 3566 - 0xdee  :  115 - 0x73
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0 -- Background 0xbe
    "11001110", -- 3569 - 0xdf1  :  206 - 0xce
    "11011110", -- 3570 - 0xdf2  :  222 - 0xde
    "11111110", -- 3571 - 0xdf3  :  254 - 0xfe
    "11111100", -- 3572 - 0xdf4  :  252 - 0xfc
    "00111000", -- 3573 - 0xdf5  :   56 - 0x38
    "11011110", -- 3574 - 0xdf6  :  222 - 0xde
    "11011110", -- 3575 - 0xdf7  :  222 - 0xde
    "11011110", -- 3576 - 0xdf8  :  222 - 0xde -- Background 0xbf
    "11011110", -- 3577 - 0xdf9  :  222 - 0xde
    "00111000", -- 3578 - 0xdfa  :   56 - 0x38
    "11111100", -- 3579 - 0xdfb  :  252 - 0xfc
    "11111110", -- 3580 - 0xdfc  :  254 - 0xfe
    "11011110", -- 3581 - 0xdfd  :  222 - 0xde
    "11001110", -- 3582 - 0xdfe  :  206 - 0xce
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "01000000", -- 3586 - 0xe02  :   64 - 0x40
    "01100000", -- 3587 - 0xe03  :   96 - 0x60
    "01100001", -- 3588 - 0xe04  :   97 - 0x61
    "00000010", -- 3589 - 0xe05  :    2 - 0x2
    "00000010", -- 3590 - 0xe06  :    2 - 0x2
    "00000111", -- 3591 - 0xe07  :    7 - 0x7
    "00000111", -- 3592 - 0xe08  :    7 - 0x7 -- Background 0xc1
    "00000100", -- 3593 - 0xe09  :    4 - 0x4
    "00000111", -- 3594 - 0xe0a  :    7 - 0x7
    "00000001", -- 3595 - 0xe0b  :    1 - 0x1
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00010000", -- 3597 - 0xe0d  :   16 - 0x10
    "00101000", -- 3598 - 0xe0e  :   40 - 0x28
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000010", -- 3602 - 0xe12  :    2 - 0x2
    "00000110", -- 3603 - 0xe13  :    6 - 0x6
    "11100110", -- 3604 - 0xe14  :  230 - 0xe6
    "10100000", -- 3605 - 0xe15  :  160 - 0xa0
    "10100000", -- 3606 - 0xe16  :  160 - 0xa0
    "11110000", -- 3607 - 0xe17  :  240 - 0xf0
    "11110000", -- 3608 - 0xe18  :  240 - 0xf0 -- Background 0xc3
    "00110000", -- 3609 - 0xe19  :   48 - 0x30
    "11000000", -- 3610 - 0xe1a  :  192 - 0xc0
    "10000000", -- 3611 - 0xe1b  :  128 - 0x80
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00001000", -- 3613 - 0xe1d  :    8 - 0x8
    "00010100", -- 3614 - 0xe1e  :   20 - 0x14
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xc4
    "00000101", -- 3617 - 0xe21  :    5 - 0x5
    "00000111", -- 3618 - 0xe22  :    7 - 0x7
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000001", -- 3623 - 0xe27  :    1 - 0x1
    "00000010", -- 3624 - 0xe28  :    2 - 0x2 -- Background 0xc5
    "00000111", -- 3625 - 0xe29  :    7 - 0x7
    "00100111", -- 3626 - 0xe2a  :   39 - 0x27
    "01010011", -- 3627 - 0xe2b  :   83 - 0x53
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000010", -- 3629 - 0xe2d  :    2 - 0x2
    "00000101", -- 3630 - 0xe2e  :    5 - 0x5
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00000000", -- 3632 - 0xe30  :    0 - 0x0 -- Background 0xc6
    "00000000", -- 3633 - 0xe31  :    0 - 0x0
    "00000000", -- 3634 - 0xe32  :    0 - 0x0
    "00000000", -- 3635 - 0xe33  :    0 - 0x0
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "01100000", -- 3637 - 0xe35  :   96 - 0x60
    "11011000", -- 3638 - 0xe36  :  216 - 0xd8
    "10110000", -- 3639 - 0xe37  :  176 - 0xb0
    "11101000", -- 3640 - 0xe38  :  232 - 0xe8 -- Background 0xc7
    "01111000", -- 3641 - 0xe39  :  120 - 0x78
    "10110110", -- 3642 - 0xe3a  :  182 - 0xb6
    "11100100", -- 3643 - 0xe3b  :  228 - 0xe4
    "00000110", -- 3644 - 0xe3c  :    6 - 0x6
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xc8
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "01000000", -- 3650 - 0xe42  :   64 - 0x40
    "00100000", -- 3651 - 0xe43  :   32 - 0x20
    "01000000", -- 3652 - 0xe44  :   64 - 0x40
    "00000111", -- 3653 - 0xe45  :    7 - 0x7
    "00000101", -- 3654 - 0xe46  :    5 - 0x5
    "00001101", -- 3655 - 0xe47  :   13 - 0xd
    "00001101", -- 3656 - 0xe48  :   13 - 0xd -- Background 0xc9
    "00000101", -- 3657 - 0xe49  :    5 - 0x5
    "00000011", -- 3658 - 0xe4a  :    3 - 0x3
    "01000011", -- 3659 - 0xe4b  :   67 - 0x43
    "00100000", -- 3660 - 0xe4c  :   32 - 0x20
    "01000000", -- 3661 - 0xe4d  :   64 - 0x40
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Background 0xca
    "00011100", -- 3665 - 0xe51  :   28 - 0x1c
    "00011000", -- 3666 - 0xe52  :   24 - 0x18
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "10000000", -- 3669 - 0xe55  :  128 - 0x80
    "11100000", -- 3670 - 0xe56  :  224 - 0xe0
    "10010000", -- 3671 - 0xe57  :  144 - 0x90
    "11110000", -- 3672 - 0xe58  :  240 - 0xf0 -- Background 0xcb
    "10010000", -- 3673 - 0xe59  :  144 - 0x90
    "11110000", -- 3674 - 0xe5a  :  240 - 0xf0
    "10000000", -- 3675 - 0xe5b  :  128 - 0x80
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00011000", -- 3677 - 0xe5d  :   24 - 0x18
    "00011100", -- 3678 - 0xe5e  :   28 - 0x1c
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xcc
    "00001000", -- 3681 - 0xe61  :    8 - 0x8
    "00000100", -- 3682 - 0xe62  :    4 - 0x4
    "00001000", -- 3683 - 0xe63  :    8 - 0x8
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "01000110", -- 3685 - 0xe65  :   70 - 0x46
    "00101111", -- 3686 - 0xe66  :   47 - 0x2f
    "01001110", -- 3687 - 0xe67  :   78 - 0x4e
    "00001101", -- 3688 - 0xe68  :   13 - 0xd -- Background 0xcd
    "00001011", -- 3689 - 0xe69  :   11 - 0xb
    "00001111", -- 3690 - 0xe6a  :   15 - 0xf
    "00000110", -- 3691 - 0xe6b  :    6 - 0x6
    "00000011", -- 3692 - 0xe6c  :    3 - 0x3
    "00011100", -- 3693 - 0xe6d  :   28 - 0x1c
    "00010100", -- 3694 - 0xe6e  :   20 - 0x14
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000110", -- 3701 - 0xe75  :    6 - 0x6
    "00000100", -- 3702 - 0xe76  :    4 - 0x4
    "10000110", -- 3703 - 0xe77  :  134 - 0x86
    "11000000", -- 3704 - 0xe78  :  192 - 0xc0 -- Background 0xcf
    "01100000", -- 3705 - 0xe79  :   96 - 0x60
    "10100000", -- 3706 - 0xe7a  :  160 - 0xa0
    "11000000", -- 3707 - 0xe7b  :  192 - 0xc0
    "01000000", -- 3708 - 0xe7c  :   64 - 0x40
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000100", -- 3716 - 0xe84  :    4 - 0x4
    "00001110", -- 3717 - 0xe85  :   14 - 0xe
    "00111111", -- 3718 - 0xe86  :   63 - 0x3f
    "00111001", -- 3719 - 0xe87  :   57 - 0x39
    "01110000", -- 3720 - 0xe88  :  112 - 0x70 -- Background 0xd1
    "01111000", -- 3721 - 0xe89  :  120 - 0x78
    "00111111", -- 3722 - 0xe8a  :   63 - 0x3f
    "00111111", -- 3723 - 0xe8b  :   63 - 0x3f
    "00000011", -- 3724 - 0xe8c  :    3 - 0x3
    "00001100", -- 3725 - 0xe8d  :   12 - 0xc
    "00001110", -- 3726 - 0xe8e  :   14 - 0xe
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000000", -- 3728 - 0xe90  :    0 - 0x0 -- Background 0xd2
    "00000000", -- 3729 - 0xe91  :    0 - 0x0
    "00000000", -- 3730 - 0xe92  :    0 - 0x0
    "00001000", -- 3731 - 0xe93  :    8 - 0x8
    "11011000", -- 3732 - 0xe94  :  216 - 0xd8
    "11111100", -- 3733 - 0xe95  :  252 - 0xfc
    "11111100", -- 3734 - 0xe96  :  252 - 0xfc
    "10011100", -- 3735 - 0xe97  :  156 - 0x9c
    "00001100", -- 3736 - 0xe98  :   12 - 0xc -- Background 0xd3
    "10011100", -- 3737 - 0xe99  :  156 - 0x9c
    "11111000", -- 3738 - 0xe9a  :  248 - 0xf8
    "01111000", -- 3739 - 0xe9b  :  120 - 0x78
    "10001000", -- 3740 - 0xe9c  :  136 - 0x88
    "00110000", -- 3741 - 0xe9d  :   48 - 0x30
    "00111000", -- 3742 - 0xe9e  :   56 - 0x38
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000001", -- 3748 - 0xea4  :    1 - 0x1
    "00001011", -- 3749 - 0xea5  :   11 - 0xb
    "00011111", -- 3750 - 0xea6  :   31 - 0x1f
    "00111001", -- 3751 - 0xea7  :   57 - 0x39
    "01110000", -- 3752 - 0xea8  :  112 - 0x70 -- Background 0xd5
    "01111000", -- 3753 - 0xea9  :  120 - 0x78
    "00111111", -- 3754 - 0xeaa  :   63 - 0x3f
    "00111111", -- 3755 - 0xeab  :   63 - 0x3f
    "00000011", -- 3756 - 0xeac  :    3 - 0x3
    "00111000", -- 3757 - 0xead  :   56 - 0x38
    "00011100", -- 3758 - 0xeae  :   28 - 0x1c
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "11000000", -- 3763 - 0xeb3  :  192 - 0xc0
    "11001000", -- 3764 - 0xeb4  :  200 - 0xc8
    "11111000", -- 3765 - 0xeb5  :  248 - 0xf8
    "11111100", -- 3766 - 0xeb6  :  252 - 0xfc
    "10011100", -- 3767 - 0xeb7  :  156 - 0x9c
    "00001100", -- 3768 - 0xeb8  :   12 - 0xc -- Background 0xd7
    "10011100", -- 3769 - 0xeb9  :  156 - 0x9c
    "11111000", -- 3770 - 0xeba  :  248 - 0xf8
    "01111000", -- 3771 - 0xebb  :  120 - 0x78
    "11100010", -- 3772 - 0xebc  :  226 - 0xe2
    "00011110", -- 3773 - 0xebd  :   30 - 0x1e
    "00001100", -- 3774 - 0xebe  :   12 - 0xc
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xd8
    "00110000", -- 3777 - 0xec1  :   48 - 0x30
    "00111100", -- 3778 - 0xec2  :   60 - 0x3c
    "01111100", -- 3779 - 0xec3  :  124 - 0x7c
    "01111100", -- 3780 - 0xec4  :  124 - 0x7c
    "00111110", -- 3781 - 0xec5  :   62 - 0x3e
    "00011100", -- 3782 - 0xec6  :   28 - 0x1c
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- Background 0xd9
    "00001110", -- 3785 - 0xec9  :   14 - 0xe
    "00111110", -- 3786 - 0xeca  :   62 - 0x3e
    "01111110", -- 3787 - 0xecb  :  126 - 0x7e
    "01111110", -- 3788 - 0xecc  :  126 - 0x7e
    "00111100", -- 3789 - 0xecd  :   60 - 0x3c
    "00001100", -- 3790 - 0xece  :   12 - 0xc
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Background 0xda
    "00100000", -- 3793 - 0xed1  :   32 - 0x20
    "01111110", -- 3794 - 0xed2  :  126 - 0x7e
    "01111110", -- 3795 - 0xed3  :  126 - 0x7e
    "01111110", -- 3796 - 0xed4  :  126 - 0x7e
    "00111100", -- 3797 - 0xed5  :   60 - 0x3c
    "00111000", -- 3798 - 0xed6  :   56 - 0x38
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0 -- Background 0xdb
    "00011100", -- 3801 - 0xed9  :   28 - 0x1c
    "00111110", -- 3802 - 0xeda  :   62 - 0x3e
    "01111110", -- 3803 - 0xedb  :  126 - 0x7e
    "01111110", -- 3804 - 0xedc  :  126 - 0x7e
    "00111100", -- 3805 - 0xedd  :   60 - 0x3c
    "00010000", -- 3806 - 0xede  :   16 - 0x10
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000001", -- 3811 - 0xee3  :    1 - 0x1
    "00000011", -- 3812 - 0xee4  :    3 - 0x3
    "00000001", -- 3813 - 0xee5  :    1 - 0x1
    "00000001", -- 3814 - 0xee6  :    1 - 0x1
    "00001111", -- 3815 - 0xee7  :   15 - 0xf
    "00000111", -- 3816 - 0xee8  :    7 - 0x7 -- Background 0xdd
    "00000111", -- 3817 - 0xee9  :    7 - 0x7
    "00000111", -- 3818 - 0xeea  :    7 - 0x7
    "00011111", -- 3819 - 0xeeb  :   31 - 0x1f
    "00001111", -- 3820 - 0xeec  :   15 - 0xf
    "00000111", -- 3821 - 0xeed  :    7 - 0x7
    "00000011", -- 3822 - 0xeee  :    3 - 0x3
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Background 0xde
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "10000000", -- 3828 - 0xef4  :  128 - 0x80
    "10000000", -- 3829 - 0xef5  :  128 - 0x80
    "10010000", -- 3830 - 0xef6  :  144 - 0x90
    "11110000", -- 3831 - 0xef7  :  240 - 0xf0
    "11100000", -- 3832 - 0xef8  :  224 - 0xe0 -- Background 0xdf
    "11100000", -- 3833 - 0xef9  :  224 - 0xe0
    "11110000", -- 3834 - 0xefa  :  240 - 0xf0
    "11110000", -- 3835 - 0xefb  :  240 - 0xf0
    "11100000", -- 3836 - 0xefc  :  224 - 0xe0
    "11000000", -- 3837 - 0xefd  :  192 - 0xc0
    "11000000", -- 3838 - 0xefe  :  192 - 0xc0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00001111", -- 3840 - 0xf00  :   15 - 0xf -- Background 0xe0
    "00011111", -- 3841 - 0xf01  :   31 - 0x1f
    "00011111", -- 3842 - 0xf02  :   31 - 0x1f
    "00111111", -- 3843 - 0xf03  :   63 - 0x3f
    "01111111", -- 3844 - 0xf04  :  127 - 0x7f
    "11111111", -- 3845 - 0xf05  :  255 - 0xff
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11111111", -- 3848 - 0xf08  :  255 - 0xff -- Background 0xe1
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "01111111", -- 3850 - 0xf0a  :  127 - 0x7f
    "00111111", -- 3851 - 0xf0b  :   63 - 0x3f
    "00111111", -- 3852 - 0xf0c  :   63 - 0x3f
    "00011111", -- 3853 - 0xf0d  :   31 - 0x1f
    "00001111", -- 3854 - 0xf0e  :   15 - 0xf
    "00000111", -- 3855 - 0xf0f  :    7 - 0x7
    "11111110", -- 3856 - 0xf10  :  254 - 0xfe -- Background 0xe2
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "00001111", -- 3859 - 0xf13  :   15 - 0xf
    "10111111", -- 3860 - 0xf14  :  191 - 0xbf
    "10100011", -- 3861 - 0xf15  :  163 - 0xa3
    "11110111", -- 3862 - 0xf16  :  247 - 0xf7
    "11110111", -- 3863 - 0xf17  :  247 - 0xf7
    "11111111", -- 3864 - 0xf18  :  255 - 0xff -- Background 0xe3
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "00111111", -- 3866 - 0xf1a  :   63 - 0x3f
    "00011111", -- 3867 - 0xf1b  :   31 - 0x1f
    "11111110", -- 3868 - 0xf1c  :  254 - 0xfe
    "11111100", -- 3869 - 0xf1d  :  252 - 0xfc
    "11111000", -- 3870 - 0xf1e  :  248 - 0xf8
    "11110000", -- 3871 - 0xf1f  :  240 - 0xf0
    "00001111", -- 3872 - 0xf20  :   15 - 0xf -- Background 0xe4
    "00011111", -- 3873 - 0xf21  :   31 - 0x1f
    "00011111", -- 3874 - 0xf22  :   31 - 0x1f
    "00111111", -- 3875 - 0xf23  :   63 - 0x3f
    "01111111", -- 3876 - 0xf24  :  127 - 0x7f
    "11111111", -- 3877 - 0xf25  :  255 - 0xff
    "11111111", -- 3878 - 0xf26  :  255 - 0xff
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff -- Background 0xe5
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "01111110", -- 3882 - 0xf2a  :  126 - 0x7e
    "00111111", -- 3883 - 0xf2b  :   63 - 0x3f
    "00111111", -- 3884 - 0xf2c  :   63 - 0x3f
    "00011111", -- 3885 - 0xf2d  :   31 - 0x1f
    "00001111", -- 3886 - 0xf2e  :   15 - 0xf
    "00000111", -- 3887 - 0xf2f  :    7 - 0x7
    "11111110", -- 3888 - 0xf30  :  254 - 0xfe -- Background 0xe6
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "11100011", -- 3891 - 0xf33  :  227 - 0xe3
    "00010111", -- 3892 - 0xf34  :   23 - 0x17
    "10110111", -- 3893 - 0xf35  :  183 - 0xb7
    "10111111", -- 3894 - 0xf36  :  191 - 0xbf
    "11111111", -- 3895 - 0xf37  :  255 - 0xff
    "11111111", -- 3896 - 0xf38  :  255 - 0xff -- Background 0xe7
    "11111111", -- 3897 - 0xf39  :  255 - 0xff
    "00111111", -- 3898 - 0xf3a  :   63 - 0x3f
    "00001111", -- 3899 - 0xf3b  :   15 - 0xf
    "00001110", -- 3900 - 0xf3c  :   14 - 0xe
    "11111100", -- 3901 - 0xf3d  :  252 - 0xfc
    "11111000", -- 3902 - 0xf3e  :  248 - 0xf8
    "11110000", -- 3903 - 0xf3f  :  240 - 0xf0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xe8
    "00000101", -- 3905 - 0xf41  :    5 - 0x5
    "00000111", -- 3906 - 0xf42  :    7 - 0x7
    "00000011", -- 3907 - 0xf43  :    3 - 0x3
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "00000000", -- 3915 - 0xf4b  :    0 - 0x0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000011", -- 3920 - 0xf50  :    3 - 0x3 -- Background 0xea
    "10011110", -- 3921 - 0xf51  :  158 - 0x9e
    "00001110", -- 3922 - 0xf52  :   14 - 0xe
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 3929 - 0xf59  :    0 - 0x0
    "00000000", -- 3930 - 0xf5a  :    0 - 0x0
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000100", -- 3940 - 0xf64  :    4 - 0x4
    "00001110", -- 3941 - 0xf65  :   14 - 0xe
    "00001111", -- 3942 - 0xf66  :   15 - 0xf
    "00001011", -- 3943 - 0xf67  :   11 - 0xb
    "00001111", -- 3944 - 0xf68  :   15 - 0xf -- Background 0xed
    "00001100", -- 3945 - 0xf69  :   12 - 0xc
    "00001111", -- 3946 - 0xf6a  :   15 - 0xf
    "00001111", -- 3947 - 0xf6b  :   15 - 0xf
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "01111111", -- 3949 - 0xf6d  :  127 - 0x7f
    "11010101", -- 3950 - 0xf6e  :  213 - 0xd5
    "01111111", -- 3951 - 0xf6f  :  127 - 0x7f
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00100000", -- 3956 - 0xf74  :   32 - 0x20
    "01110000", -- 3957 - 0xf75  :  112 - 0x70
    "11110000", -- 3958 - 0xf76  :  240 - 0xf0
    "11100000", -- 3959 - 0xf77  :  224 - 0xe0
    "11110000", -- 3960 - 0xf78  :  240 - 0xf0 -- Background 0xef
    "00110000", -- 3961 - 0xf79  :   48 - 0x30
    "11110000", -- 3962 - 0xf7a  :  240 - 0xf0
    "11110000", -- 3963 - 0xf7b  :  240 - 0xf0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "11111110", -- 3965 - 0xf7d  :  254 - 0xfe
    "01010101", -- 3966 - 0xf7e  :   85 - 0x55
    "11111110", -- 3967 - 0xf7f  :  254 - 0xfe
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000100", -- 3972 - 0xf84  :    4 - 0x4
    "00001110", -- 3973 - 0xf85  :   14 - 0xe
    "00001111", -- 3974 - 0xf86  :   15 - 0xf
    "00001011", -- 3975 - 0xf87  :   11 - 0xb
    "00001111", -- 3976 - 0xf88  :   15 - 0xf -- Background 0xf1
    "00001100", -- 3977 - 0xf89  :   12 - 0xc
    "00001111", -- 3978 - 0xf8a  :   15 - 0xf
    "00001111", -- 3979 - 0xf8b  :   15 - 0xf
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "01111111", -- 3981 - 0xf8d  :  127 - 0x7f
    "10101010", -- 3982 - 0xf8e  :  170 - 0xaa
    "01111111", -- 3983 - 0xf8f  :  127 - 0x7f
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00100000", -- 3988 - 0xf94  :   32 - 0x20
    "01110000", -- 3989 - 0xf95  :  112 - 0x70
    "11110000", -- 3990 - 0xf96  :  240 - 0xf0
    "11100000", -- 3991 - 0xf97  :  224 - 0xe0
    "11110000", -- 3992 - 0xf98  :  240 - 0xf0 -- Background 0xf3
    "00110000", -- 3993 - 0xf99  :   48 - 0x30
    "11110000", -- 3994 - 0xf9a  :  240 - 0xf0
    "11110000", -- 3995 - 0xf9b  :  240 - 0xf0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "11111110", -- 3997 - 0xf9d  :  254 - 0xfe
    "10101011", -- 3998 - 0xf9e  :  171 - 0xab
    "11111110", -- 3999 - 0xf9f  :  254 - 0xfe
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Background 0xf4
    "00010101", -- 4001 - 0xfa1  :   21 - 0x15
    "00001010", -- 4002 - 0xfa2  :   10 - 0xa
    "00000101", -- 4003 - 0xfa3  :    5 - 0x5
    "00000010", -- 4004 - 0xfa4  :    2 - 0x2
    "00000101", -- 4005 - 0xfa5  :    5 - 0x5
    "00000111", -- 4006 - 0xfa6  :    7 - 0x7
    "00000111", -- 4007 - 0xfa7  :    7 - 0x7
    "00111100", -- 4008 - 0xfa8  :   60 - 0x3c -- Background 0xf5
    "01111011", -- 4009 - 0xfa9  :  123 - 0x7b
    "01111011", -- 4010 - 0xfaa  :  123 - 0x7b
    "01111111", -- 4011 - 0xfab  :  127 - 0x7f
    "01111110", -- 4012 - 0xfac  :  126 - 0x7e
    "01111111", -- 4013 - 0xfad  :  127 - 0x7f
    "00111110", -- 4014 - 0xfae  :   62 - 0x3e
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Background 0xf6
    "01010000", -- 4017 - 0xfb1  :   80 - 0x50
    "10100000", -- 4018 - 0xfb2  :  160 - 0xa0
    "01000000", -- 4019 - 0xfb3  :   64 - 0x40
    "10100000", -- 4020 - 0xfb4  :  160 - 0xa0
    "01000000", -- 4021 - 0xfb5  :   64 - 0x40
    "11100000", -- 4022 - 0xfb6  :  224 - 0xe0
    "11100000", -- 4023 - 0xfb7  :  224 - 0xe0
    "01111000", -- 4024 - 0xfb8  :  120 - 0x78 -- Background 0xf7
    "10111100", -- 4025 - 0xfb9  :  188 - 0xbc
    "10111000", -- 4026 - 0xfba  :  184 - 0xb8
    "10111110", -- 4027 - 0xfbb  :  190 - 0xbe
    "01111100", -- 4028 - 0xfbc  :  124 - 0x7c
    "11111110", -- 4029 - 0xfbd  :  254 - 0xfe
    "01111000", -- 4030 - 0xfbe  :  120 - 0x78
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000011", -- 4032 - 0xfc0  :    3 - 0x3 -- Background 0xf8
    "00000011", -- 4033 - 0xfc1  :    3 - 0x3
    "00000000", -- 4034 - 0xfc2  :    0 - 0x0
    "00000011", -- 4035 - 0xfc3  :    3 - 0x3
    "00000111", -- 4036 - 0xfc4  :    7 - 0x7
    "00000110", -- 4037 - 0xfc5  :    6 - 0x6
    "00000111", -- 4038 - 0xfc6  :    7 - 0x7
    "00000000", -- 4039 - 0xfc7  :    0 - 0x0
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0 -- Background 0xf9
    "00011111", -- 4041 - 0xfc9  :   31 - 0x1f
    "00011111", -- 4042 - 0xfca  :   31 - 0x1f
    "00001111", -- 4043 - 0xfcb  :   15 - 0xf
    "00000011", -- 4044 - 0xfcc  :    3 - 0x3
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "11100000", -- 4048 - 0xfd0  :  224 - 0xe0 -- Background 0xfa
    "11100000", -- 4049 - 0xfd1  :  224 - 0xe0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00110000", -- 4051 - 0xfd3  :   48 - 0x30
    "01110000", -- 4052 - 0xfd4  :  112 - 0x70
    "01100000", -- 4053 - 0xfd5  :   96 - 0x60
    "01110000", -- 4054 - 0xfd6  :  112 - 0x70
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0 -- Background 0xfb
    "11111000", -- 4057 - 0xfd9  :  248 - 0xf8
    "11111000", -- 4058 - 0xfda  :  248 - 0xf8
    "11110000", -- 4059 - 0xfdb  :  240 - 0xf0
    "11000000", -- 4060 - 0xfdc  :  192 - 0xc0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00111000", -- 4064 - 0xfe0  :   56 - 0x38 -- Background 0xfc
    "00111000", -- 4065 - 0xfe1  :   56 - 0x38
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "01111100", -- 4067 - 0xfe3  :  124 - 0x7c
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "00111000", -- 4069 - 0xfe5  :   56 - 0x38
    "00111000", -- 4070 - 0xfe6  :   56 - 0x38
    "01111100", -- 4071 - 0xfe7  :  124 - 0x7c
    "01111100", -- 4072 - 0xfe8  :  124 - 0x7c -- Background 0xfd
    "01111100", -- 4073 - 0xfe9  :  124 - 0x7c
    "01111100", -- 4074 - 0xfea  :  124 - 0x7c
    "00111000", -- 4075 - 0xfeb  :   56 - 0x38
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "01111100", -- 4077 - 0xfed  :  124 - 0x7c
    "01111100", -- 4078 - 0xfee  :  124 - 0x7c
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "00010001", -- 4082 - 0xff2  :   17 - 0x11
    "11010111", -- 4083 - 0xff3  :  215 - 0xd7
    "11010111", -- 4084 - 0xff4  :  215 - 0xd7
    "11010111", -- 4085 - 0xff5  :  215 - 0xd7
    "00010001", -- 4086 - 0xff6  :   17 - 0x11
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "11100110", -- 4090 - 0xffa  :  230 - 0xe6
    "11110110", -- 4091 - 0xffb  :  246 - 0xf6
    "11110110", -- 4092 - 0xffc  :  246 - 0xf6
    "11110110", -- 4093 - 0xffd  :  246 - 0xf6
    "11100110", -- 4094 - 0xffe  :  230 - 0xe6
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
