------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : random_256x256_gray.ppm 
--- Filas    : 256 
--- Columnas : 256 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 8 bits
--- De cada palabra hay 3 bits para rojo y verde y 2 para azul: "RRRGGGBB" 256 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_8b_random_256x256_gray is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(16-1 downto 0);
    dout : out std_logic_vector(8-1 downto 0) 
  );
end ROM_RGB_8b_random_256x256_gray;


architecture BEHAVIORAL of ROM_RGB_8b_random_256x256_gray is
  signal addr_int  : natural range 0 to 2**16-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBB"
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "11111111",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10110110",
       "10110110",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10010010",
       "10010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11011011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

