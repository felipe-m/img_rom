//-   Background Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_LAWN_BG
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table both color planes
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      12'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      12'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      12'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout  = 8'b00000101; //    8 :   5 - 0x5 -- plane 1
      12'h9: dout  = 8'b01010101; //    9 :  85 - 0x55
      12'hA: dout  = 8'b01010101; //   10 :  85 - 0x55
      12'hB: dout  = 8'b01010000; //   11 :  80 - 0x50
      12'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout  = 8'b00000101; //   16 :   5 - 0x5 -- Background 0x1
      12'h11: dout  = 8'b01010101; //   17 :  85 - 0x55
      12'h12: dout  = 8'b01010101; //   18 :  85 - 0x55
      12'h13: dout  = 8'b01010000; //   19 :  80 - 0x50
      12'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      12'h15: dout  = 8'b00000000; //   21 :   0 - 0x0
      12'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      12'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout  = 8'b00000101; //   24 :   5 - 0x5 -- plane 1
      12'h19: dout  = 8'b01010101; //   25 :  85 - 0x55
      12'h1A: dout  = 8'b01010101; //   26 :  85 - 0x55
      12'h1B: dout  = 8'b01010000; //   27 :  80 - 0x50
      12'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout  = 8'b00000101; //   32 :   5 - 0x5 -- Background 0x2
      12'h21: dout  = 8'b01010000; //   33 :  80 - 0x50
      12'h22: dout  = 8'b00000101; //   34 :   5 - 0x5
      12'h23: dout  = 8'b01010000; //   35 :  80 - 0x50
      12'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      12'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      12'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout  = 8'b00000101; //   40 :   5 - 0x5 -- plane 1
      12'h29: dout  = 8'b01010000; //   41 :  80 - 0x50
      12'h2A: dout  = 8'b00000101; //   42 :   5 - 0x5
      12'h2B: dout  = 8'b01010000; //   43 :  80 - 0x50
      12'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout  = 8'b00000101; //   48 :   5 - 0x5 -- Background 0x3
      12'h31: dout  = 8'b01010000; //   49 :  80 - 0x50
      12'h32: dout  = 8'b00000101; //   50 :   5 - 0x5
      12'h33: dout  = 8'b01010000; //   51 :  80 - 0x50
      12'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      12'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      12'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      12'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout  = 8'b00000101; //   56 :   5 - 0x5 -- plane 1
      12'h39: dout  = 8'b01010101; //   57 :  85 - 0x55
      12'h3A: dout  = 8'b01010101; //   58 :  85 - 0x55
      12'h3B: dout  = 8'b01010000; //   59 :  80 - 0x50
      12'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00000101; //   64 :   5 - 0x5 -- Background 0x4
      12'h41: dout  = 8'b01010101; //   65 :  85 - 0x55
      12'h42: dout  = 8'b01010101; //   66 :  85 - 0x55
      12'h43: dout  = 8'b01010000; //   67 :  80 - 0x50
      12'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      12'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout  = 8'b00000101; //   72 :   5 - 0x5 -- plane 1
      12'h49: dout  = 8'b01010101; //   73 :  85 - 0x55
      12'h4A: dout  = 8'b01010101; //   74 :  85 - 0x55
      12'h4B: dout  = 8'b01010000; //   75 :  80 - 0x50
      12'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Background 0x5
      12'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      12'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      12'h53: dout  = 8'b00000000; //   83 :   0 - 0x0
      12'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      12'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      12'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout  = 8'b00001110; //   88 :  14 - 0xe -- plane 1
      12'h59: dout  = 8'b00000111; //   89 :   7 - 0x7
      12'h5A: dout  = 8'b00001000; //   90 :   8 - 0x8
      12'h5B: dout  = 8'b01100000; //   91 :  96 - 0x60
      12'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout  = 8'b00001010; //   93 :  10 - 0xa
      12'h5E: dout  = 8'b00000001; //   94 :   1 - 0x1
      12'h5F: dout  = 8'b00010101; //   95 :  21 - 0x15
      12'h60: dout  = 8'b01010101; //   96 :  85 - 0x55 -- Background 0x6
      12'h61: dout  = 8'b01010101; //   97 :  85 - 0x55
      12'h62: dout  = 8'b01010100; //   98 :  84 - 0x54
      12'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      12'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      12'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout  = 8'b00010101; //  103 :  21 - 0x15
      12'h68: dout  = 8'b01010101; //  104 :  85 - 0x55 -- plane 1
      12'h69: dout  = 8'b01010101; //  105 :  85 - 0x55
      12'h6A: dout  = 8'b01010100; //  106 :  84 - 0x54
      12'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout  = 8'b00010110; //  111 :  22 - 0x16
      12'h70: dout  = 8'b10101010; //  112 : 170 - 0xaa -- Background 0x7
      12'h71: dout  = 8'b10011010; //  113 : 154 - 0x9a
      12'h72: dout  = 8'b10010100; //  114 : 148 - 0x94
      12'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      12'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      12'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      12'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      12'h77: dout  = 8'b00010110; //  119 :  22 - 0x16
      12'h78: dout  = 8'b01010101; //  120 :  85 - 0x55 -- plane 1
      12'h79: dout  = 8'b01010101; //  121 :  85 - 0x55
      12'h7A: dout  = 8'b10010100; //  122 : 148 - 0x94
      12'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout  = 8'b00010110; //  127 :  22 - 0x16
      12'h80: dout  = 8'b01010000; //  128 :  80 - 0x50 -- Background 0x8
      12'h81: dout  = 8'b00000101; //  129 :   5 - 0x5
      12'h82: dout  = 8'b10010100; //  130 : 148 - 0x94
      12'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout  = 8'b00000000; //  133 :   0 - 0x0
      12'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout  = 8'b00010101; //  135 :  21 - 0x15
      12'h88: dout  = 8'b01010000; //  136 :  80 - 0x50 -- plane 1
      12'h89: dout  = 8'b00000101; //  137 :   5 - 0x5
      12'h8A: dout  = 8'b01010100; //  138 :  84 - 0x54
      12'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout  = 8'b00010110; //  143 :  22 - 0x16
      12'h90: dout  = 8'b01010000; //  144 :  80 - 0x50 -- Background 0x9
      12'h91: dout  = 8'b00000101; //  145 :   5 - 0x5
      12'h92: dout  = 8'b10010100; //  146 : 148 - 0x94
      12'h93: dout  = 8'b00000000; //  147 :   0 - 0x0
      12'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      12'h95: dout  = 8'b00000000; //  149 :   0 - 0x0
      12'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout  = 8'b00010110; //  151 :  22 - 0x16
      12'h98: dout  = 8'b01010101; //  152 :  85 - 0x55 -- plane 1
      12'h99: dout  = 8'b01010101; //  153 :  85 - 0x55
      12'h9A: dout  = 8'b10010100; //  154 : 148 - 0x94
      12'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout  = 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout  = 8'b00010110; //  159 :  22 - 0x16
      12'hA0: dout  = 8'b10100110; //  160 : 166 - 0xa6 -- Background 0xa
      12'hA1: dout  = 8'b10101010; //  161 : 170 - 0xaa
      12'hA2: dout  = 8'b10010100; //  162 : 148 - 0x94
      12'hA3: dout  = 8'b00000000; //  163 :   0 - 0x0
      12'hA4: dout  = 8'b00000000; //  164 :   0 - 0x0
      12'hA5: dout  = 8'b00000000; //  165 :   0 - 0x0
      12'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout  = 8'b00010101; //  167 :  21 - 0x15
      12'hA8: dout  = 8'b01010101; //  168 :  85 - 0x55 -- plane 1
      12'hA9: dout  = 8'b01010101; //  169 :  85 - 0x55
      12'hAA: dout  = 8'b01010100; //  170 :  84 - 0x54
      12'hAB: dout  = 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout  = 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout  = 8'b00010101; //  175 :  21 - 0x15
      12'hB0: dout  = 8'b01010101; //  176 :  85 - 0x55 -- Background 0xb
      12'hB1: dout  = 8'b01010101; //  177 :  85 - 0x55
      12'hB2: dout  = 8'b01010100; //  178 :  84 - 0x54
      12'hB3: dout  = 8'b00000000; //  179 :   0 - 0x0
      12'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout  = 8'b00001110; //  183 :  14 - 0xe
      12'hB8: dout  = 8'b00000111; //  184 :   7 - 0x7 -- plane 1
      12'hB9: dout  = 8'b00001000; //  185 :   8 - 0x8
      12'hBA: dout  = 8'b01110100; //  186 : 116 - 0x74
      12'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout  = 8'b11011100; //  188 : 220 - 0xdc
      12'hBD: dout  = 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout  = 8'b00010101; //  190 :  21 - 0x15
      12'hBF: dout  = 8'b01010101; //  191 :  85 - 0x55
      12'hC0: dout  = 8'b01010101; //  192 :  85 - 0x55 -- Background 0xc
      12'hC1: dout  = 8'b01010100; //  193 :  84 - 0x54
      12'hC2: dout  = 8'b00000000; //  194 :   0 - 0x0
      12'hC3: dout  = 8'b00000000; //  195 :   0 - 0x0
      12'hC4: dout  = 8'b00000000; //  196 :   0 - 0x0
      12'hC5: dout  = 8'b00000000; //  197 :   0 - 0x0
      12'hC6: dout  = 8'b00011010; //  198 :  26 - 0x1a
      12'hC7: dout  = 8'b10011101; //  199 : 157 - 0x9d
      12'hC8: dout  = 8'b01110110; //  200 : 118 - 0x76 -- plane 1
      12'hC9: dout  = 8'b10100100; //  201 : 164 - 0xa4
      12'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout  = 8'b00000000; //  204 :   0 - 0x0
      12'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout  = 8'b00010101; //  206 :  21 - 0x15
      12'hCF: dout  = 8'b01010101; //  207 :  85 - 0x55
      12'hD0: dout  = 8'b01010101; //  208 :  85 - 0x55 -- Background 0xd
      12'hD1: dout  = 8'b01010100; //  209 :  84 - 0x54
      12'hD2: dout  = 8'b00000000; //  210 :   0 - 0x0
      12'hD3: dout  = 8'b00000000; //  211 :   0 - 0x0
      12'hD4: dout  = 8'b00000000; //  212 :   0 - 0x0
      12'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout  = 8'b00010111; //  214 :  23 - 0x17
      12'hD7: dout  = 8'b01010101; //  215 :  85 - 0x55
      12'hD8: dout  = 8'b01010101; //  216 :  85 - 0x55 -- plane 1
      12'hD9: dout  = 8'b11010100; //  217 : 212 - 0xd4
      12'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout  = 8'b00000000; //  219 :   0 - 0x0
      12'hDC: dout  = 8'b00000000; //  220 :   0 - 0x0
      12'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout  = 8'b00010101; //  222 :  21 - 0x15
      12'hDF: dout  = 8'b01010000; //  223 :  80 - 0x50
      12'hE0: dout  = 8'b00000101; //  224 :   5 - 0x5 -- Background 0xe
      12'hE1: dout  = 8'b01010100; //  225 :  84 - 0x54
      12'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      12'hE3: dout  = 8'b00000000; //  227 :   0 - 0x0
      12'hE4: dout  = 8'b00000000; //  228 :   0 - 0x0
      12'hE5: dout  = 8'b00000000; //  229 :   0 - 0x0
      12'hE6: dout  = 8'b00010101; //  230 :  21 - 0x15
      12'hE7: dout  = 8'b01010000; //  231 :  80 - 0x50
      12'hE8: dout  = 8'b00000101; //  232 :   5 - 0x5 -- plane 1
      12'hE9: dout  = 8'b01010100; //  233 :  84 - 0x54
      12'hEA: dout  = 8'b00000000; //  234 :   0 - 0x0
      12'hEB: dout  = 8'b00000000; //  235 :   0 - 0x0
      12'hEC: dout  = 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout  = 8'b00010101; //  238 :  21 - 0x15
      12'hEF: dout  = 8'b01010000; //  239 :  80 - 0x50
      12'hF0: dout  = 8'b00000101; //  240 :   5 - 0x5 -- Background 0xf
      12'hF1: dout  = 8'b01010100; //  241 :  84 - 0x54
      12'hF2: dout  = 8'b00000000; //  242 :   0 - 0x0
      12'hF3: dout  = 8'b00000000; //  243 :   0 - 0x0
      12'hF4: dout  = 8'b00000000; //  244 :   0 - 0x0
      12'hF5: dout  = 8'b00000000; //  245 :   0 - 0x0
      12'hF6: dout  = 8'b00010111; //  246 :  23 - 0x17
      12'hF7: dout  = 8'b01010101; //  247 :  85 - 0x55
      12'hF8: dout  = 8'b01010101; //  248 :  85 - 0x55 -- plane 1
      12'hF9: dout  = 8'b11010100; //  249 : 212 - 0xd4
      12'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout  = 8'b00010101; //  254 :  21 - 0x15
      12'hFF: dout  = 8'b01010101; //  255 :  85 - 0x55
      12'h100: dout  = 8'b01010101; //  256 :  85 - 0x55 -- Background 0x10
      12'h101: dout  = 8'b01010100; //  257 :  84 - 0x54
      12'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      12'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      12'h106: dout  = 8'b00011010; //  262 :  26 - 0x1a
      12'h107: dout  = 8'b10011101; //  263 : 157 - 0x9d
      12'h108: dout  = 8'b01110110; //  264 : 118 - 0x76 -- plane 1
      12'h109: dout  = 8'b10100100; //  265 : 164 - 0xa4
      12'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout  = 8'b00010101; //  270 :  21 - 0x15
      12'h10F: dout  = 8'b01010101; //  271 :  85 - 0x55
      12'h110: dout  = 8'b01010101; //  272 :  85 - 0x55 -- Background 0x11
      12'h111: dout  = 8'b01010100; //  273 :  84 - 0x54
      12'h112: dout  = 8'b00000000; //  274 :   0 - 0x0
      12'h113: dout  = 8'b00000000; //  275 :   0 - 0x0
      12'h114: dout  = 8'b00000000; //  276 :   0 - 0x0
      12'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      12'h116: dout  = 8'b00001110; //  278 :  14 - 0xe
      12'h117: dout  = 8'b00000111; //  279 :   7 - 0x7
      12'h118: dout  = 8'b00001000; //  280 :   8 - 0x8 -- plane 1
      12'h119: dout  = 8'b01111010; //  281 : 122 - 0x7a
      12'h11A: dout  = 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout  = 8'b11010001; //  283 : 209 - 0xd1
      12'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout  = 8'b00010101; //  285 :  21 - 0x15
      12'h11E: dout  = 8'b01010101; //  286 :  85 - 0x55
      12'h11F: dout  = 8'b01010101; //  287 :  85 - 0x55
      12'h120: dout  = 8'b01010101; //  288 :  85 - 0x55 -- Background 0x12
      12'h121: dout  = 8'b01010101; //  289 :  85 - 0x55
      12'h122: dout  = 8'b01000000; //  290 :  64 - 0x40
      12'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout  = 8'b00010101; //  293 :  21 - 0x15
      12'h126: dout  = 8'b01010101; //  294 :  85 - 0x55
      12'h127: dout  = 8'b01010101; //  295 :  85 - 0x55
      12'h128: dout  = 8'b01010101; //  296 :  85 - 0x55 -- plane 1
      12'h129: dout  = 8'b01010101; //  297 :  85 - 0x55
      12'h12A: dout  = 8'b01000000; //  298 :  64 - 0x40
      12'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout  = 8'b00010110; //  301 :  22 - 0x16
      12'h12E: dout  = 8'b10100101; //  302 : 165 - 0xa5
      12'h12F: dout  = 8'b01010101; //  303 :  85 - 0x55
      12'h130: dout  = 8'b01010101; //  304 :  85 - 0x55 -- Background 0x13
      12'h131: dout  = 8'b10101001; //  305 : 169 - 0xa9
      12'h132: dout  = 8'b01000000; //  306 :  64 - 0x40
      12'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout  = 8'b00010110; //  309 :  22 - 0x16
      12'h136: dout  = 8'b01010101; //  310 :  85 - 0x55
      12'h137: dout  = 8'b01101010; //  311 : 106 - 0x6a
      12'h138: dout  = 8'b10010101; //  312 : 149 - 0x95 -- plane 1
      12'h139: dout  = 8'b01011001; //  313 :  89 - 0x59
      12'h13A: dout  = 8'b01000000; //  314 :  64 - 0x40
      12'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00010110; //  317 :  22 - 0x16
      12'h13E: dout  = 8'b01000000; //  318 :  64 - 0x40
      12'h13F: dout  = 8'b01010101; //  319 :  85 - 0x55
      12'h140: dout  = 8'b01010101; //  320 :  85 - 0x55 -- Background 0x14
      12'h141: dout  = 8'b01011001; //  321 :  89 - 0x59
      12'h142: dout  = 8'b01000000; //  322 :  64 - 0x40
      12'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      12'h145: dout  = 8'b00010101; //  325 :  21 - 0x15
      12'h146: dout  = 8'b01000000; //  326 :  64 - 0x40
      12'h147: dout  = 8'b01010101; //  327 :  85 - 0x55
      12'h148: dout  = 8'b01010101; //  328 :  85 - 0x55 -- plane 1
      12'h149: dout  = 8'b01010101; //  329 :  85 - 0x55
      12'h14A: dout  = 8'b01000000; //  330 :  64 - 0x40
      12'h14B: dout  = 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout  = 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout  = 8'b00010110; //  333 :  22 - 0x16
      12'h14E: dout  = 8'b01000000; //  334 :  64 - 0x40
      12'h14F: dout  = 8'b01010101; //  335 :  85 - 0x55
      12'h150: dout  = 8'b01010101; //  336 :  85 - 0x55 -- Background 0x15
      12'h151: dout  = 8'b01011001; //  337 :  89 - 0x59
      12'h152: dout  = 8'b01000000; //  338 :  64 - 0x40
      12'h153: dout  = 8'b00000000; //  339 :   0 - 0x0
      12'h154: dout  = 8'b00000000; //  340 :   0 - 0x0
      12'h155: dout  = 8'b00010110; //  341 :  22 - 0x16
      12'h156: dout  = 8'b01010101; //  342 :  85 - 0x55
      12'h157: dout  = 8'b01101010; //  343 : 106 - 0x6a
      12'h158: dout  = 8'b10010101; //  344 : 149 - 0x95 -- plane 1
      12'h159: dout  = 8'b01011001; //  345 :  89 - 0x59
      12'h15A: dout  = 8'b01000000; //  346 :  64 - 0x40
      12'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout  = 8'b00010110; //  349 :  22 - 0x16
      12'h15E: dout  = 8'b10100101; //  350 : 165 - 0xa5
      12'h15F: dout  = 8'b01010101; //  351 :  85 - 0x55
      12'h160: dout  = 8'b01010101; //  352 :  85 - 0x55 -- Background 0x16
      12'h161: dout  = 8'b10101001; //  353 : 169 - 0xa9
      12'h162: dout  = 8'b01000000; //  354 :  64 - 0x40
      12'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout  = 8'b00010101; //  357 :  21 - 0x15
      12'h166: dout  = 8'b01010101; //  358 :  85 - 0x55
      12'h167: dout  = 8'b01010101; //  359 :  85 - 0x55
      12'h168: dout  = 8'b01010101; //  360 :  85 - 0x55 -- plane 1
      12'h169: dout  = 8'b01010101; //  361 :  85 - 0x55
      12'h16A: dout  = 8'b01000000; //  362 :  64 - 0x40
      12'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout  = 8'b00010101; //  365 :  21 - 0x15
      12'h16E: dout  = 8'b01010101; //  366 :  85 - 0x55
      12'h16F: dout  = 8'b01010101; //  367 :  85 - 0x55
      12'h170: dout  = 8'b01010101; //  368 :  85 - 0x55 -- Background 0x17
      12'h171: dout  = 8'b01010101; //  369 :  85 - 0x55
      12'h172: dout  = 8'b01000000; //  370 :  64 - 0x40
      12'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      12'h175: dout  = 8'b00010100; //  373 :  20 - 0x14
      12'h176: dout  = 8'b00000110; //  374 :   6 - 0x6
      12'h177: dout  = 8'b00001000; //  375 :   8 - 0x8
      12'h178: dout  = 8'b10110111; //  376 : 183 - 0xb7 -- plane 1
      12'h179: dout  = 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout  = 8'b10001011; //  378 : 139 - 0x8b
      12'h17B: dout  = 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout  = 8'b00010101; //  380 :  21 - 0x15
      12'h17D: dout  = 8'b01010101; //  381 :  85 - 0x55
      12'h17E: dout  = 8'b01010101; //  382 :  85 - 0x55
      12'h17F: dout  = 8'b01010101; //  383 :  85 - 0x55
      12'h180: dout  = 8'b01010101; //  384 :  85 - 0x55 -- Background 0x18
      12'h181: dout  = 8'b01000000; //  385 :  64 - 0x40
      12'h182: dout  = 8'b00000000; //  386 :   0 - 0x0
      12'h183: dout  = 8'b00000000; //  387 :   0 - 0x0
      12'h184: dout  = 8'b00011010; //  388 :  26 - 0x1a
      12'h185: dout  = 8'b01010111; //  389 :  87 - 0x57
      12'h186: dout  = 8'b01010101; //  390 :  85 - 0x55
      12'h187: dout  = 8'b01011101; //  391 :  93 - 0x5d
      12'h188: dout  = 8'b01011010; //  392 :  90 - 0x5a -- plane 1
      12'h189: dout  = 8'b01000000; //  393 :  64 - 0x40
      12'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout  = 8'b00011010; //  396 :  26 - 0x1a
      12'h18D: dout  = 8'b01010111; //  397 :  87 - 0x57
      12'h18E: dout  = 8'b01010101; //  398 :  85 - 0x55
      12'h18F: dout  = 8'b01011101; //  399 :  93 - 0x5d
      12'h190: dout  = 8'b01011010; //  400 :  90 - 0x5a -- Background 0x19
      12'h191: dout  = 8'b01000000; //  401 :  64 - 0x40
      12'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      12'h193: dout  = 8'b00000000; //  403 :   0 - 0x0
      12'h194: dout  = 8'b00010101; //  404 :  21 - 0x15
      12'h195: dout  = 8'b01010111; //  405 :  87 - 0x57
      12'h196: dout  = 8'b01011010; //  406 :  90 - 0x5a
      12'h197: dout  = 8'b01011101; //  407 :  93 - 0x5d
      12'h198: dout  = 8'b01010101; //  408 :  85 - 0x55 -- plane 1
      12'h199: dout  = 8'b01000000; //  409 :  64 - 0x40
      12'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout  = 8'b00010000; //  412 :  16 - 0x10
      12'h19D: dout  = 8'b00010101; //  413 :  21 - 0x15
      12'h19E: dout  = 8'b01011010; //  414 :  90 - 0x5a
      12'h19F: dout  = 8'b01010101; //  415 :  85 - 0x55
      12'h1A0: dout  = 8'b01010101; //  416 :  85 - 0x55 -- Background 0x1a
      12'h1A1: dout  = 8'b01000000; //  417 :  64 - 0x40
      12'h1A2: dout  = 8'b00000000; //  418 :   0 - 0x0
      12'h1A3: dout  = 8'b00000000; //  419 :   0 - 0x0
      12'h1A4: dout  = 8'b00010000; //  420 :  16 - 0x10
      12'h1A5: dout  = 8'b00010101; //  421 :  21 - 0x15
      12'h1A6: dout  = 8'b01011010; //  422 :  90 - 0x5a
      12'h1A7: dout  = 8'b01010101; //  423 :  85 - 0x55
      12'h1A8: dout  = 8'b01010101; //  424 :  85 - 0x55 -- plane 1
      12'h1A9: dout  = 8'b01000000; //  425 :  64 - 0x40
      12'h1AA: dout  = 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout  = 8'b00010000; //  428 :  16 - 0x10
      12'h1AD: dout  = 8'b00010101; //  429 :  21 - 0x15
      12'h1AE: dout  = 8'b01011010; //  430 :  90 - 0x5a
      12'h1AF: dout  = 8'b01010101; //  431 :  85 - 0x55
      12'h1B0: dout  = 8'b01010101; //  432 :  85 - 0x55 -- Background 0x1b
      12'h1B1: dout  = 8'b01000000; //  433 :  64 - 0x40
      12'h1B2: dout  = 8'b00000000; //  434 :   0 - 0x0
      12'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      12'h1B4: dout  = 8'b00010101; //  436 :  21 - 0x15
      12'h1B5: dout  = 8'b01010111; //  437 :  87 - 0x57
      12'h1B6: dout  = 8'b01011010; //  438 :  90 - 0x5a
      12'h1B7: dout  = 8'b01011101; //  439 :  93 - 0x5d
      12'h1B8: dout  = 8'b01010101; //  440 :  85 - 0x55 -- plane 1
      12'h1B9: dout  = 8'b01000000; //  441 :  64 - 0x40
      12'h1BA: dout  = 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout  = 8'b00011010; //  444 :  26 - 0x1a
      12'h1BD: dout  = 8'b01010111; //  445 :  87 - 0x57
      12'h1BE: dout  = 8'b01010101; //  446 :  85 - 0x55
      12'h1BF: dout  = 8'b01011101; //  447 :  93 - 0x5d
      12'h1C0: dout  = 8'b01011010; //  448 :  90 - 0x5a -- Background 0x1c
      12'h1C1: dout  = 8'b01000000; //  449 :  64 - 0x40
      12'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout  = 8'b00011010; //  452 :  26 - 0x1a
      12'h1C5: dout  = 8'b01010111; //  453 :  87 - 0x57
      12'h1C6: dout  = 8'b01010101; //  454 :  85 - 0x55
      12'h1C7: dout  = 8'b01011101; //  455 :  93 - 0x5d
      12'h1C8: dout  = 8'b01011010; //  456 :  90 - 0x5a -- plane 1
      12'h1C9: dout  = 8'b01000000; //  457 :  64 - 0x40
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout  = 8'b00010101; //  460 :  21 - 0x15
      12'h1CD: dout  = 8'b01010101; //  461 :  85 - 0x55
      12'h1CE: dout  = 8'b01010101; //  462 :  85 - 0x55
      12'h1CF: dout  = 8'b01010101; //  463 :  85 - 0x55
      12'h1D0: dout  = 8'b01010101; //  464 :  85 - 0x55 -- Background 0x1d
      12'h1D1: dout  = 8'b01000000; //  465 :  64 - 0x40
      12'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      12'h1D4: dout  = 8'b00010100; //  468 :  20 - 0x14
      12'h1D5: dout  = 8'b00000011; //  469 :   3 - 0x3
      12'h1D6: dout  = 8'b00001000; //  470 :   8 - 0x8
      12'h1D7: dout  = 8'b10101101; //  471 : 173 - 0xad
      12'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- plane 1
      12'h1D9: dout  = 8'b10010011; //  473 : 147 - 0x93
      12'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout  = 8'b00010101; //  475 :  21 - 0x15
      12'h1DC: dout  = 8'b01010101; //  476 :  85 - 0x55
      12'h1DD: dout  = 8'b01010101; //  477 :  85 - 0x55
      12'h1DE: dout  = 8'b01010101; //  478 :  85 - 0x55
      12'h1DF: dout  = 8'b01010101; //  479 :  85 - 0x55
      12'h1E0: dout  = 8'b01010101; //  480 :  85 - 0x55 -- Background 0x1e
      12'h1E1: dout  = 8'b01010000; //  481 :  80 - 0x50
      12'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout  = 8'b00010101; //  483 :  21 - 0x15
      12'h1E4: dout  = 8'b01110101; //  484 : 117 - 0x75
      12'h1E5: dout  = 8'b01010101; //  485 :  85 - 0x55
      12'h1E6: dout  = 8'b01010111; //  486 :  87 - 0x57
      12'h1E7: dout  = 8'b01010101; //  487 :  85 - 0x55
      12'h1E8: dout  = 8'b01010111; //  488 :  87 - 0x57 -- plane 1
      12'h1E9: dout  = 8'b01010000; //  489 :  80 - 0x50
      12'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout  = 8'b00011101; //  491 :  29 - 0x1d
      12'h1EC: dout  = 8'b01010101; //  492 :  85 - 0x55
      12'h1ED: dout  = 8'b01110101; //  493 : 117 - 0x75
      12'h1EE: dout  = 8'b01010101; //  494 :  85 - 0x55
      12'h1EF: dout  = 8'b01011101; //  495 :  93 - 0x5d
      12'h1F0: dout  = 8'b01010101; //  496 :  85 - 0x55 -- Background 0x1f
      12'h1F1: dout  = 8'b01010000; //  497 :  80 - 0x50
      12'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      12'h1F3: dout  = 8'b00010101; //  499 :  21 - 0x15
      12'h1F4: dout  = 8'b01010111; //  500 :  87 - 0x57
      12'h1F5: dout  = 8'b01010101; //  501 :  85 - 0x55
      12'h1F6: dout  = 8'b01010101; //  502 :  85 - 0x55
      12'h1F7: dout  = 8'b01010101; //  503 :  85 - 0x55
      12'h1F8: dout  = 8'b01110101; //  504 : 117 - 0x75 -- plane 1
      12'h1F9: dout  = 8'b01010000; //  505 :  80 - 0x50
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00010101; //  507 :  21 - 0x15
      12'h1FC: dout  = 8'b01010101; //  508 :  85 - 0x55
      12'h1FD: dout  = 8'b01010101; //  509 :  85 - 0x55
      12'h1FE: dout  = 8'b00000001; //  510 :   1 - 0x1
      12'h1FF: dout  = 8'b01010101; //  511 :  85 - 0x55
      12'h200: dout  = 8'b01010101; //  512 :  85 - 0x55 -- Background 0x20
      12'h201: dout  = 8'b11010000; //  513 : 208 - 0xd0
      12'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout  = 8'b00010111; //  515 :  23 - 0x17
      12'h204: dout  = 8'b01010101; //  516 :  85 - 0x55
      12'h205: dout  = 8'b01010101; //  517 :  85 - 0x55
      12'h206: dout  = 8'b00000001; //  518 :   1 - 0x1
      12'h207: dout  = 8'b01010111; //  519 :  87 - 0x57
      12'h208: dout  = 8'b01010101; //  520 :  85 - 0x55 -- plane 1
      12'h209: dout  = 8'b01010000; //  521 :  80 - 0x50
      12'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout  = 8'b00010101; //  523 :  21 - 0x15
      12'h20C: dout  = 8'b01011101; //  524 :  93 - 0x5d
      12'h20D: dout  = 8'b01010101; //  525 :  85 - 0x55
      12'h20E: dout  = 8'b00000001; //  526 :   1 - 0x1
      12'h20F: dout  = 8'b01010101; //  527 :  85 - 0x55
      12'h210: dout  = 8'b01010101; //  528 :  85 - 0x55 -- Background 0x21
      12'h211: dout  = 8'b01010000; //  529 :  80 - 0x50
      12'h212: dout  = 8'b00000000; //  530 :   0 - 0x0
      12'h213: dout  = 8'b00010101; //  531 :  21 - 0x15
      12'h214: dout  = 8'b01010101; //  532 :  85 - 0x55
      12'h215: dout  = 8'b01110101; //  533 : 117 - 0x75
      12'h216: dout  = 8'b01010101; //  534 :  85 - 0x55
      12'h217: dout  = 8'b01010101; //  535 :  85 - 0x55
      12'h218: dout  = 8'b01110101; //  536 : 117 - 0x75 -- plane 1
      12'h219: dout  = 8'b01010000; //  537 :  80 - 0x50
      12'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout  = 8'b00011101; //  539 :  29 - 0x1d
      12'h21C: dout  = 8'b01010101; //  540 :  85 - 0x55
      12'h21D: dout  = 8'b01010101; //  541 :  85 - 0x55
      12'h21E: dout  = 8'b01010101; //  542 :  85 - 0x55
      12'h21F: dout  = 8'b01110101; //  543 : 117 - 0x75
      12'h220: dout  = 8'b01010101; //  544 :  85 - 0x55 -- Background 0x22
      12'h221: dout  = 8'b01010000; //  545 :  80 - 0x50
      12'h222: dout  = 8'b00000000; //  546 :   0 - 0x0
      12'h223: dout  = 8'b00010101; //  547 :  21 - 0x15
      12'h224: dout  = 8'b01110101; //  548 : 117 - 0x75
      12'h225: dout  = 8'b01010101; //  549 :  85 - 0x55
      12'h226: dout  = 8'b11010101; //  550 : 213 - 0xd5
      12'h227: dout  = 8'b01010101; //  551 :  85 - 0x55
      12'h228: dout  = 8'b01010111; //  552 :  87 - 0x57 -- plane 1
      12'h229: dout  = 8'b01010000; //  553 :  80 - 0x50
      12'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      12'h22B: dout  = 8'b00010101; //  555 :  21 - 0x15
      12'h22C: dout  = 8'b01010101; //  556 :  85 - 0x55
      12'h22D: dout  = 8'b01010101; //  557 :  85 - 0x55
      12'h22E: dout  = 8'b01010101; //  558 :  85 - 0x55
      12'h22F: dout  = 8'b01010101; //  559 :  85 - 0x55
      12'h230: dout  = 8'b01010101; //  560 :  85 - 0x55 -- Background 0x23
      12'h231: dout  = 8'b01010000; //  561 :  80 - 0x50
      12'h232: dout  = 8'b00000000; //  562 :   0 - 0x0
      12'h233: dout  = 8'b00011001; //  563 :  25 - 0x19
      12'h234: dout  = 8'b00001101; //  564 :  13 - 0xd
      12'h235: dout  = 8'b00001000; //  565 :   8 - 0x8
      12'h236: dout  = 8'b11110111; //  566 : 247 - 0xf7
      12'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout  = 8'b01100111; //  568 : 103 - 0x67 -- plane 1
      12'h239: dout  = 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout  = 8'b00010101; //  570 :  21 - 0x15
      12'h23B: dout  = 8'b01010101; //  571 :  85 - 0x55
      12'h23C: dout  = 8'b01010101; //  572 :  85 - 0x55
      12'h23D: dout  = 8'b01010101; //  573 :  85 - 0x55
      12'h23E: dout  = 8'b01010101; //  574 :  85 - 0x55
      12'h23F: dout  = 8'b01010101; //  575 :  85 - 0x55
      12'h240: dout  = 8'b01010000; //  576 :  80 - 0x50 -- Background 0x24
      12'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout  = 8'b00011010; //  578 :  26 - 0x1a
      12'h243: dout  = 8'b10101001; //  579 : 169 - 0xa9
      12'h244: dout  = 8'b10101010; //  580 : 170 - 0xaa
      12'h245: dout  = 8'b10011001; //  581 : 153 - 0x99
      12'h246: dout  = 8'b01011001; //  582 :  89 - 0x59
      12'h247: dout  = 8'b10101010; //  583 : 170 - 0xaa
      12'h248: dout  = 8'b10010000; //  584 : 144 - 0x90 -- plane 1
      12'h249: dout  = 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout  = 8'b00011001; //  586 :  25 - 0x19
      12'h24B: dout  = 8'b01011001; //  587 :  89 - 0x59
      12'h24C: dout  = 8'b10010101; //  588 : 149 - 0x95
      12'h24D: dout  = 8'b10011001; //  589 : 153 - 0x99
      12'h24E: dout  = 8'b01011001; //  590 :  89 - 0x59
      12'h24F: dout  = 8'b10010101; //  591 : 149 - 0x95
      12'h250: dout  = 8'b10010000; //  592 : 144 - 0x90 -- Background 0x25
      12'h251: dout  = 8'b00000000; //  593 :   0 - 0x0
      12'h252: dout  = 8'b00010101; //  594 :  21 - 0x15
      12'h253: dout  = 8'b01011001; //  595 :  89 - 0x59
      12'h254: dout  = 8'b10010101; //  596 : 149 - 0x95
      12'h255: dout  = 8'b10011001; //  597 : 153 - 0x99
      12'h256: dout  = 8'b01011001; //  598 :  89 - 0x59
      12'h257: dout  = 8'b10010101; //  599 : 149 - 0x95
      12'h258: dout  = 8'b01010000; //  600 :  80 - 0x50 -- plane 1
      12'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout  = 8'b00010000; //  602 :  16 - 0x10
      12'h25B: dout  = 8'b00010101; //  603 :  21 - 0x15
      12'h25C: dout  = 8'b10010101; //  604 : 149 - 0x95
      12'h25D: dout  = 8'b10011010; //  605 : 154 - 0x9a
      12'h25E: dout  = 8'b10101001; //  606 : 169 - 0xa9
      12'h25F: dout  = 8'b01010101; //  607 :  85 - 0x55
      12'h260: dout  = 8'b01010000; //  608 :  80 - 0x50 -- Background 0x26
      12'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout  = 8'b00010000; //  610 :  16 - 0x10
      12'h263: dout  = 8'b00010101; //  611 :  21 - 0x15
      12'h264: dout  = 8'b01010101; //  612 :  85 - 0x55
      12'h265: dout  = 8'b01010101; //  613 :  85 - 0x55
      12'h266: dout  = 8'b01010101; //  614 :  85 - 0x55
      12'h267: dout  = 8'b01010101; //  615 :  85 - 0x55
      12'h268: dout  = 8'b01010000; //  616 :  80 - 0x50 -- plane 1
      12'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout  = 8'b00010000; //  618 :  16 - 0x10
      12'h26B: dout  = 8'b00010101; //  619 :  21 - 0x15
      12'h26C: dout  = 8'b10101010; //  620 : 170 - 0xaa
      12'h26D: dout  = 8'b10011001; //  621 : 153 - 0x99
      12'h26E: dout  = 8'b01011001; //  622 :  89 - 0x59
      12'h26F: dout  = 8'b01010101; //  623 :  85 - 0x55
      12'h270: dout  = 8'b01010000; //  624 :  80 - 0x50 -- Background 0x27
      12'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      12'h272: dout  = 8'b00010101; //  626 :  21 - 0x15
      12'h273: dout  = 8'b01011001; //  627 :  89 - 0x59
      12'h274: dout  = 8'b10010101; //  628 : 149 - 0x95
      12'h275: dout  = 8'b10011001; //  629 : 153 - 0x99
      12'h276: dout  = 8'b01011001; //  630 :  89 - 0x59
      12'h277: dout  = 8'b10010101; //  631 : 149 - 0x95
      12'h278: dout  = 8'b01010000; //  632 :  80 - 0x50 -- plane 1
      12'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout  = 8'b00011001; //  634 :  25 - 0x19
      12'h27B: dout  = 8'b01011001; //  635 :  89 - 0x59
      12'h27C: dout  = 8'b10010101; //  636 : 149 - 0x95
      12'h27D: dout  = 8'b10011001; //  637 : 153 - 0x99
      12'h27E: dout  = 8'b01011001; //  638 :  89 - 0x59
      12'h27F: dout  = 8'b10010101; //  639 : 149 - 0x95
      12'h280: dout  = 8'b10010000; //  640 : 144 - 0x90 -- Background 0x28
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00011010; //  642 :  26 - 0x1a
      12'h283: dout  = 8'b10101001; //  643 : 169 - 0xa9
      12'h284: dout  = 8'b10010101; //  644 : 149 - 0x95
      12'h285: dout  = 8'b10011010; //  645 : 154 - 0x9a
      12'h286: dout  = 8'b10101001; //  646 : 169 - 0xa9
      12'h287: dout  = 8'b10101010; //  647 : 170 - 0xaa
      12'h288: dout  = 8'b10010000; //  648 : 144 - 0x90 -- plane 1
      12'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout  = 8'b00010101; //  650 :  21 - 0x15
      12'h28B: dout  = 8'b01010101; //  651 :  85 - 0x55
      12'h28C: dout  = 8'b01010101; //  652 :  85 - 0x55
      12'h28D: dout  = 8'b01010101; //  653 :  85 - 0x55
      12'h28E: dout  = 8'b01010101; //  654 :  85 - 0x55
      12'h28F: dout  = 8'b01010101; //  655 :  85 - 0x55
      12'h290: dout  = 8'b01010000; //  656 :  80 - 0x50 -- Background 0x29
      12'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout  = 8'b00011001; //  658 :  25 - 0x19
      12'h293: dout  = 8'b00000011; //  659 :   3 - 0x3
      12'h294: dout  = 8'b00001000; //  660 :   8 - 0x8
      12'h295: dout  = 8'b10111110; //  661 : 190 - 0xbe
      12'h296: dout  = 8'b00000000; //  662 :   0 - 0x0
      12'h297: dout  = 8'b10000110; //  663 : 134 - 0x86
      12'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- plane 1
      12'h299: dout  = 8'b00010101; //  665 :  21 - 0x15
      12'h29A: dout  = 8'b01010111; //  666 :  87 - 0x57
      12'h29B: dout  = 8'b01010101; //  667 :  85 - 0x55
      12'h29C: dout  = 8'b01010101; //  668 :  85 - 0x55
      12'h29D: dout  = 8'b01010111; //  669 :  87 - 0x57
      12'h29E: dout  = 8'b01010101; //  670 :  85 - 0x55
      12'h29F: dout  = 8'b01010000; //  671 :  80 - 0x50
      12'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Background 0x2a
      12'h2A1: dout  = 8'b00010101; //  673 :  21 - 0x15
      12'h2A2: dout  = 8'b01010111; //  674 :  87 - 0x57
      12'h2A3: dout  = 8'b01101010; //  675 : 106 - 0x6a
      12'h2A4: dout  = 8'b01010110; //  676 :  86 - 0x56
      12'h2A5: dout  = 8'b10100111; //  677 : 167 - 0xa7
      12'h2A6: dout  = 8'b01010101; //  678 :  85 - 0x55
      12'h2A7: dout  = 8'b01010000; //  679 :  80 - 0x50
      12'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- plane 1
      12'h2A9: dout  = 8'b00010101; //  681 :  21 - 0x15
      12'h2AA: dout  = 8'b01010111; //  682 :  87 - 0x57
      12'h2AB: dout  = 8'b01101010; //  683 : 106 - 0x6a
      12'h2AC: dout  = 8'b01010110; //  684 :  86 - 0x56
      12'h2AD: dout  = 8'b10100111; //  685 : 167 - 0xa7
      12'h2AE: dout  = 8'b01010101; //  686 :  85 - 0x55
      12'h2AF: dout  = 8'b01010000; //  687 :  80 - 0x50
      12'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Background 0x2b
      12'h2B1: dout  = 8'b00010101; //  689 :  21 - 0x15
      12'h2B2: dout  = 8'b01010111; //  690 :  87 - 0x57
      12'h2B3: dout  = 8'b01010101; //  691 :  85 - 0x55
      12'h2B4: dout  = 8'b01110101; //  692 : 117 - 0x75
      12'h2B5: dout  = 8'b01010111; //  693 :  87 - 0x57
      12'h2B6: dout  = 8'b01010101; //  694 :  85 - 0x55
      12'h2B7: dout  = 8'b01010000; //  695 :  80 - 0x50
      12'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- plane 1
      12'h2B9: dout  = 8'b00010000; //  697 :  16 - 0x10
      12'h2BA: dout  = 8'b00010101; //  698 :  21 - 0x15
      12'h2BB: dout  = 8'b01010101; //  699 :  85 - 0x55
      12'h2BC: dout  = 8'b01110101; //  700 : 117 - 0x75
      12'h2BD: dout  = 8'b01010101; //  701 :  85 - 0x55
      12'h2BE: dout  = 8'b01010101; //  702 :  85 - 0x55
      12'h2BF: dout  = 8'b01010000; //  703 :  80 - 0x50
      12'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Background 0x2c
      12'h2C1: dout  = 8'b00010000; //  705 :  16 - 0x10
      12'h2C2: dout  = 8'b00010101; //  706 :  21 - 0x15
      12'h2C3: dout  = 8'b01010101; //  707 :  85 - 0x55
      12'h2C4: dout  = 8'b01110101; //  708 : 117 - 0x75
      12'h2C5: dout  = 8'b01010101; //  709 :  85 - 0x55
      12'h2C6: dout  = 8'b01010101; //  710 :  85 - 0x55
      12'h2C7: dout  = 8'b01010000; //  711 :  80 - 0x50
      12'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout  = 8'b00010000; //  713 :  16 - 0x10
      12'h2CA: dout  = 8'b00010101; //  714 :  21 - 0x15
      12'h2CB: dout  = 8'b01010101; //  715 :  85 - 0x55
      12'h2CC: dout  = 8'b01110101; //  716 : 117 - 0x75
      12'h2CD: dout  = 8'b01010101; //  717 :  85 - 0x55
      12'h2CE: dout  = 8'b01010101; //  718 :  85 - 0x55
      12'h2CF: dout  = 8'b01010000; //  719 :  80 - 0x50
      12'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Background 0x2d
      12'h2D1: dout  = 8'b00010101; //  721 :  21 - 0x15
      12'h2D2: dout  = 8'b01010111; //  722 :  87 - 0x57
      12'h2D3: dout  = 8'b01010101; //  723 :  85 - 0x55
      12'h2D4: dout  = 8'b01110101; //  724 : 117 - 0x75
      12'h2D5: dout  = 8'b01010111; //  725 :  87 - 0x57
      12'h2D6: dout  = 8'b01010101; //  726 :  85 - 0x55
      12'h2D7: dout  = 8'b01010000; //  727 :  80 - 0x50
      12'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- plane 1
      12'h2D9: dout  = 8'b00010101; //  729 :  21 - 0x15
      12'h2DA: dout  = 8'b01010111; //  730 :  87 - 0x57
      12'h2DB: dout  = 8'b01101010; //  731 : 106 - 0x6a
      12'h2DC: dout  = 8'b01010110; //  732 :  86 - 0x56
      12'h2DD: dout  = 8'b10100111; //  733 : 167 - 0xa7
      12'h2DE: dout  = 8'b01010101; //  734 :  85 - 0x55
      12'h2DF: dout  = 8'b01010000; //  735 :  80 - 0x50
      12'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Background 0x2e
      12'h2E1: dout  = 8'b00010101; //  737 :  21 - 0x15
      12'h2E2: dout  = 8'b01010111; //  738 :  87 - 0x57
      12'h2E3: dout  = 8'b01101010; //  739 : 106 - 0x6a
      12'h2E4: dout  = 8'b01010110; //  740 :  86 - 0x56
      12'h2E5: dout  = 8'b10100111; //  741 : 167 - 0xa7
      12'h2E6: dout  = 8'b01010101; //  742 :  85 - 0x55
      12'h2E7: dout  = 8'b01010000; //  743 :  80 - 0x50
      12'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout  = 8'b00010101; //  745 :  21 - 0x15
      12'h2EA: dout  = 8'b01010111; //  746 :  87 - 0x57
      12'h2EB: dout  = 8'b01010101; //  747 :  85 - 0x55
      12'h2EC: dout  = 8'b01010101; //  748 :  85 - 0x55
      12'h2ED: dout  = 8'b01010111; //  749 :  87 - 0x57
      12'h2EE: dout  = 8'b01010101; //  750 :  85 - 0x55
      12'h2EF: dout  = 8'b01010000; //  751 :  80 - 0x50
      12'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Background 0x2f
      12'h2F1: dout  = 8'b00011001; //  753 :  25 - 0x19
      12'h2F2: dout  = 8'b00000011; //  754 :   3 - 0x3
      12'h2F3: dout  = 8'b00001000; //  755 :   8 - 0x8
      12'h2F4: dout  = 8'b11011101; //  756 : 221 - 0xdd
      12'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout  = 8'b01110011; //  758 : 115 - 0x73
      12'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout  = 8'b00010101; //  760 :  21 - 0x15 -- plane 1
      12'h2F9: dout  = 8'b01010101; //  761 :  85 - 0x55
      12'h2FA: dout  = 8'b01010101; //  762 :  85 - 0x55
      12'h2FB: dout  = 8'b01010101; //  763 :  85 - 0x55
      12'h2FC: dout  = 8'b01010101; //  764 :  85 - 0x55
      12'h2FD: dout  = 8'b01010101; //  765 :  85 - 0x55
      12'h2FE: dout  = 8'b01010101; //  766 :  85 - 0x55
      12'h2FF: dout  = 8'b01010100; //  767 :  84 - 0x54
      12'h300: dout  = 8'b00011001; //  768 :  25 - 0x19 -- Background 0x30
      12'h301: dout  = 8'b01100101; //  769 : 101 - 0x65
      12'h302: dout  = 8'b10010110; //  770 : 150 - 0x96
      12'h303: dout  = 8'b10100101; //  771 : 165 - 0xa5
      12'h304: dout  = 8'b01011010; //  772 :  90 - 0x5a
      12'h305: dout  = 8'b10010110; //  773 : 150 - 0x96
      12'h306: dout  = 8'b01011001; //  774 :  89 - 0x59
      12'h307: dout  = 8'b01100100; //  775 : 100 - 0x64
      12'h308: dout  = 8'b00011001; //  776 :  25 - 0x19 -- plane 1
      12'h309: dout  = 8'b01100101; //  777 : 101 - 0x65
      12'h30A: dout  = 8'b10010101; //  778 : 149 - 0x95
      12'h30B: dout  = 8'b01010101; //  779 :  85 - 0x55
      12'h30C: dout  = 8'b01010101; //  780 :  85 - 0x55
      12'h30D: dout  = 8'b01010110; //  781 :  86 - 0x56
      12'h30E: dout  = 8'b01011001; //  782 :  89 - 0x59
      12'h30F: dout  = 8'b01100100; //  783 : 100 - 0x64
      12'h310: dout  = 8'b00011001; //  784 :  25 - 0x19 -- Background 0x31
      12'h311: dout  = 8'b01100101; //  785 : 101 - 0x65
      12'h312: dout  = 8'b10010110; //  786 : 150 - 0x96
      12'h313: dout  = 8'b10100101; //  787 : 165 - 0xa5
      12'h314: dout  = 8'b01011010; //  788 :  90 - 0x5a
      12'h315: dout  = 8'b10010110; //  789 : 150 - 0x96
      12'h316: dout  = 8'b01011001; //  790 :  89 - 0x59
      12'h317: dout  = 8'b01100100; //  791 : 100 - 0x64
      12'h318: dout  = 8'b00010101; //  792 :  21 - 0x15 -- plane 1
      12'h319: dout  = 8'b01010101; //  793 :  85 - 0x55
      12'h31A: dout  = 8'b01010101; //  794 :  85 - 0x55
      12'h31B: dout  = 8'b01010000; //  795 :  80 - 0x50
      12'h31C: dout  = 8'b00000101; //  796 :   5 - 0x5
      12'h31D: dout  = 8'b01010101; //  797 :  85 - 0x55
      12'h31E: dout  = 8'b01010101; //  798 :  85 - 0x55
      12'h31F: dout  = 8'b01010100; //  799 :  84 - 0x54
      12'h320: dout  = 8'b00011111; //  800 :  31 - 0x1f -- Background 0x32
      12'h321: dout  = 8'b01111101; //  801 : 125 - 0x7d
      12'h322: dout  = 8'b11010101; //  802 : 213 - 0xd5
      12'h323: dout  = 8'b01010000; //  803 :  80 - 0x50
      12'h324: dout  = 8'b00000101; //  804 :   5 - 0x5
      12'h325: dout  = 8'b01010111; //  805 :  87 - 0x57
      12'h326: dout  = 8'b11111111; //  806 : 255 - 0xff
      12'h327: dout  = 8'b01110100; //  807 : 116 - 0x74
      12'h328: dout  = 8'b00010101; //  808 :  21 - 0x15 -- plane 1
      12'h329: dout  = 8'b01010101; //  809 :  85 - 0x55
      12'h32A: dout  = 8'b01010101; //  810 :  85 - 0x55
      12'h32B: dout  = 8'b01010000; //  811 :  80 - 0x50
      12'h32C: dout  = 8'b00000101; //  812 :   5 - 0x5
      12'h32D: dout  = 8'b01010101; //  813 :  85 - 0x55
      12'h32E: dout  = 8'b01010101; //  814 :  85 - 0x55
      12'h32F: dout  = 8'b01010100; //  815 :  84 - 0x54
      12'h330: dout  = 8'b00011001; //  816 :  25 - 0x19 -- Background 0x33
      12'h331: dout  = 8'b01100101; //  817 : 101 - 0x65
      12'h332: dout  = 8'b10010110; //  818 : 150 - 0x96
      12'h333: dout  = 8'b10100101; //  819 : 165 - 0xa5
      12'h334: dout  = 8'b01011010; //  820 :  90 - 0x5a
      12'h335: dout  = 8'b10010110; //  821 : 150 - 0x96
      12'h336: dout  = 8'b01011001; //  822 :  89 - 0x59
      12'h337: dout  = 8'b01100100; //  823 : 100 - 0x64
      12'h338: dout  = 8'b00011001; //  824 :  25 - 0x19 -- plane 1
      12'h339: dout  = 8'b01100101; //  825 : 101 - 0x65
      12'h33A: dout  = 8'b10010101; //  826 : 149 - 0x95
      12'h33B: dout  = 8'b01010101; //  827 :  85 - 0x55
      12'h33C: dout  = 8'b01010101; //  828 :  85 - 0x55
      12'h33D: dout  = 8'b01010110; //  829 :  86 - 0x56
      12'h33E: dout  = 8'b01011001; //  830 :  89 - 0x59
      12'h33F: dout  = 8'b01100100; //  831 : 100 - 0x64
      12'h340: dout  = 8'b00011001; //  832 :  25 - 0x19 -- Background 0x34
      12'h341: dout  = 8'b01100101; //  833 : 101 - 0x65
      12'h342: dout  = 8'b10010110; //  834 : 150 - 0x96
      12'h343: dout  = 8'b10100101; //  835 : 165 - 0xa5
      12'h344: dout  = 8'b01011010; //  836 :  90 - 0x5a
      12'h345: dout  = 8'b10010110; //  837 : 150 - 0x96
      12'h346: dout  = 8'b01011001; //  838 :  89 - 0x59
      12'h347: dout  = 8'b01100100; //  839 : 100 - 0x64
      12'h348: dout  = 8'b00010101; //  840 :  21 - 0x15 -- plane 1
      12'h349: dout  = 8'b01010101; //  841 :  85 - 0x55
      12'h34A: dout  = 8'b01010101; //  842 :  85 - 0x55
      12'h34B: dout  = 8'b01010101; //  843 :  85 - 0x55
      12'h34C: dout  = 8'b01010101; //  844 :  85 - 0x55
      12'h34D: dout  = 8'b01010101; //  845 :  85 - 0x55
      12'h34E: dout  = 8'b01010101; //  846 :  85 - 0x55
      12'h34F: dout  = 8'b01010100; //  847 :  84 - 0x54
      12'h350: dout  = 8'b00011110; //  848 :  30 - 0x1e -- Background 0x35
      12'h351: dout  = 8'b00001111; //  849 :  15 - 0xf
      12'h352: dout  = 8'b00001000; //  850 :   8 - 0x8
      12'h353: dout  = 8'b11110111; //  851 : 247 - 0xf7
      12'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout  = 8'b01100111; //  853 : 103 - 0x67
      12'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout  = 8'b00010101; //  855 :  21 - 0x15
      12'h358: dout  = 8'b01010101; //  856 :  85 - 0x55 -- plane 1
      12'h359: dout  = 8'b01010101; //  857 :  85 - 0x55
      12'h35A: dout  = 8'b01010101; //  858 :  85 - 0x55
      12'h35B: dout  = 8'b01010101; //  859 :  85 - 0x55
      12'h35C: dout  = 8'b01010101; //  860 :  85 - 0x55
      12'h35D: dout  = 8'b01010101; //  861 :  85 - 0x55
      12'h35E: dout  = 8'b01010100; //  862 :  84 - 0x54
      12'h35F: dout  = 8'b00010111; //  863 :  23 - 0x17
      12'h360: dout  = 8'b01110101; //  864 : 117 - 0x75 -- Background 0x36
      12'h361: dout  = 8'b01010110; //  865 :  86 - 0x56
      12'h362: dout  = 8'b10100101; //  866 : 165 - 0xa5
      12'h363: dout  = 8'b01011010; //  867 :  90 - 0x5a
      12'h364: dout  = 8'b10010101; //  868 : 149 - 0x95
      12'h365: dout  = 8'b01011101; //  869 :  93 - 0x5d
      12'h366: dout  = 8'b11010100; //  870 : 212 - 0xd4
      12'h367: dout  = 8'b00010101; //  871 :  21 - 0x15
      12'h368: dout  = 8'b01010101; //  872 :  85 - 0x55 -- plane 1
      12'h369: dout  = 8'b01110110; //  873 : 118 - 0x76
      12'h36A: dout  = 8'b10100101; //  874 : 165 - 0xa5
      12'h36B: dout  = 8'b01011010; //  875 :  90 - 0x5a
      12'h36C: dout  = 8'b10011101; //  876 : 157 - 0x9d
      12'h36D: dout  = 8'b01010101; //  877 :  85 - 0x55
      12'h36E: dout  = 8'b01010100; //  878 :  84 - 0x54
      12'h36F: dout  = 8'b00010111; //  879 :  23 - 0x17
      12'h370: dout  = 8'b01010101; //  880 :  85 - 0x55 -- Background 0x37
      12'h371: dout  = 8'b01110101; //  881 : 117 - 0x75
      12'h372: dout  = 8'b01010101; //  882 :  85 - 0x55
      12'h373: dout  = 8'b01010101; //  883 :  85 - 0x55
      12'h374: dout  = 8'b01011101; //  884 :  93 - 0x5d
      12'h375: dout  = 8'b01010101; //  885 :  85 - 0x55
      12'h376: dout  = 8'b11010100; //  886 : 212 - 0xd4
      12'h377: dout  = 8'b00010101; //  887 :  21 - 0x15
      12'h378: dout  = 8'b01101010; //  888 : 106 - 0x6a -- plane 1
      12'h379: dout  = 8'b01110101; //  889 : 117 - 0x75
      12'h37A: dout  = 8'b01010000; //  890 :  80 - 0x50
      12'h37B: dout  = 8'b00000101; //  891 :   5 - 0x5
      12'h37C: dout  = 8'b01011101; //  892 :  93 - 0x5d
      12'h37D: dout  = 8'b10101001; //  893 : 169 - 0xa9
      12'h37E: dout  = 8'b01010100; //  894 :  84 - 0x54
      12'h37F: dout  = 8'b00010101; //  895 :  21 - 0x15
      12'h380: dout  = 8'b01101110; //  896 : 110 - 0x6e -- Background 0x38
      12'h381: dout  = 8'b01110101; //  897 : 117 - 0x75
      12'h382: dout  = 8'b01010000; //  898 :  80 - 0x50
      12'h383: dout  = 8'b00000101; //  899 :   5 - 0x5
      12'h384: dout  = 8'b01011101; //  900 :  93 - 0x5d
      12'h385: dout  = 8'b10111001; //  901 : 185 - 0xb9
      12'h386: dout  = 8'b01010100; //  902 :  84 - 0x54
      12'h387: dout  = 8'b00010101; //  903 :  21 - 0x15
      12'h388: dout  = 8'b01101010; //  904 : 106 - 0x6a -- plane 1
      12'h389: dout  = 8'b01110101; //  905 : 117 - 0x75
      12'h38A: dout  = 8'b01010000; //  906 :  80 - 0x50
      12'h38B: dout  = 8'b00000101; //  907 :   5 - 0x5
      12'h38C: dout  = 8'b01011101; //  908 :  93 - 0x5d
      12'h38D: dout  = 8'b10101001; //  909 : 169 - 0xa9
      12'h38E: dout  = 8'b01010100; //  910 :  84 - 0x54
      12'h38F: dout  = 8'b00010111; //  911 :  23 - 0x17
      12'h390: dout  = 8'b01010101; //  912 :  85 - 0x55 -- Background 0x39
      12'h391: dout  = 8'b01110101; //  913 : 117 - 0x75
      12'h392: dout  = 8'b01010101; //  914 :  85 - 0x55
      12'h393: dout  = 8'b01010101; //  915 :  85 - 0x55
      12'h394: dout  = 8'b01011101; //  916 :  93 - 0x5d
      12'h395: dout  = 8'b01010101; //  917 :  85 - 0x55
      12'h396: dout  = 8'b11010100; //  918 : 212 - 0xd4
      12'h397: dout  = 8'b00010101; //  919 :  21 - 0x15
      12'h398: dout  = 8'b01010101; //  920 :  85 - 0x55 -- plane 1
      12'h399: dout  = 8'b01110101; //  921 : 117 - 0x75
      12'h39A: dout  = 8'b10101010; //  922 : 170 - 0xaa
      12'h39B: dout  = 8'b10101010; //  923 : 170 - 0xaa
      12'h39C: dout  = 8'b01011101; //  924 :  93 - 0x5d
      12'h39D: dout  = 8'b01010101; //  925 :  85 - 0x55
      12'h39E: dout  = 8'b01010100; //  926 :  84 - 0x54
      12'h39F: dout  = 8'b00010111; //  927 :  23 - 0x17
      12'h3A0: dout  = 8'b01110101; //  928 : 117 - 0x75 -- Background 0x3a
      12'h3A1: dout  = 8'b01010101; //  929 :  85 - 0x55
      12'h3A2: dout  = 8'b01101010; //  930 : 106 - 0x6a
      12'h3A3: dout  = 8'b10101001; //  931 : 169 - 0xa9
      12'h3A4: dout  = 8'b01010101; //  932 :  85 - 0x55
      12'h3A5: dout  = 8'b01011101; //  933 :  93 - 0x5d
      12'h3A6: dout  = 8'b11010100; //  934 : 212 - 0xd4
      12'h3A7: dout  = 8'b00010101; //  935 :  21 - 0x15
      12'h3A8: dout  = 8'b01010101; //  936 :  85 - 0x55 -- plane 1
      12'h3A9: dout  = 8'b01010101; //  937 :  85 - 0x55
      12'h3AA: dout  = 8'b01010101; //  938 :  85 - 0x55
      12'h3AB: dout  = 8'b01010101; //  939 :  85 - 0x55
      12'h3AC: dout  = 8'b01010101; //  940 :  85 - 0x55
      12'h3AD: dout  = 8'b01010101; //  941 :  85 - 0x55
      12'h3AE: dout  = 8'b01010100; //  942 :  84 - 0x54
      12'h3AF: dout  = 8'b00011110; //  943 :  30 - 0x1e
      12'h3B0: dout  = 8'b00001111; //  944 :  15 - 0xf -- Background 0x3b
      12'h3B1: dout  = 8'b00001000; //  945 :   8 - 0x8
      12'h3B2: dout  = 8'b11111000; //  946 : 248 - 0xf8
      12'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout  = 8'b01100111; //  948 : 103 - 0x67
      12'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Background 0x3c
      12'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Background 0x3d
      12'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Background 0x3e
      12'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x3f
      12'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- plane 1
      12'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Background 0x40
      12'h401: dout  = 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout  = 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout  = 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout  = 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout  = 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout  = 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- plane 1
      12'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x41
      12'h411: dout  = 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout  = 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout  = 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout  = 8'b00000000; // 1044 :   0 - 0x0
      12'h415: dout  = 8'b00000000; // 1045 :   0 - 0x0
      12'h416: dout  = 8'b00000000; // 1046 :   0 - 0x0
      12'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Background 0x42
      12'h421: dout  = 8'b00000000; // 1057 :   0 - 0x0
      12'h422: dout  = 8'b00000000; // 1058 :   0 - 0x0
      12'h423: dout  = 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout  = 8'b00000000; // 1060 :   0 - 0x0
      12'h425: dout  = 8'b00000000; // 1061 :   0 - 0x0
      12'h426: dout  = 8'b00000000; // 1062 :   0 - 0x0
      12'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- plane 1
      12'h429: dout  = 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout  = 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout  = 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout  = 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout  = 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x43
      12'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout  = 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout  = 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout  = 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout  = 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- plane 1
      12'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout  = 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x44
      12'h441: dout  = 8'b00000000; // 1089 :   0 - 0x0
      12'h442: dout  = 8'b00000000; // 1090 :   0 - 0x0
      12'h443: dout  = 8'b00000000; // 1091 :   0 - 0x0
      12'h444: dout  = 8'b00000000; // 1092 :   0 - 0x0
      12'h445: dout  = 8'b00000000; // 1093 :   0 - 0x0
      12'h446: dout  = 8'b00000000; // 1094 :   0 - 0x0
      12'h447: dout  = 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout  = 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout  = 8'b00000000; // 1097 :   0 - 0x0
      12'h44A: dout  = 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout  = 8'b00000000; // 1099 :   0 - 0x0
      12'h44C: dout  = 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout  = 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout  = 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x45
      12'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      12'h452: dout  = 8'b00000000; // 1106 :   0 - 0x0
      12'h453: dout  = 8'b00000000; // 1107 :   0 - 0x0
      12'h454: dout  = 8'b00000000; // 1108 :   0 - 0x0
      12'h455: dout  = 8'b00000000; // 1109 :   0 - 0x0
      12'h456: dout  = 8'b00000000; // 1110 :   0 - 0x0
      12'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout  = 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout  = 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout  = 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout  = 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout  = 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout  = 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x46
      12'h461: dout  = 8'b00000000; // 1121 :   0 - 0x0
      12'h462: dout  = 8'b00000000; // 1122 :   0 - 0x0
      12'h463: dout  = 8'b00000000; // 1123 :   0 - 0x0
      12'h464: dout  = 8'b00000000; // 1124 :   0 - 0x0
      12'h465: dout  = 8'b00000000; // 1125 :   0 - 0x0
      12'h466: dout  = 8'b00000000; // 1126 :   0 - 0x0
      12'h467: dout  = 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout  = 8'b00000000; // 1128 :   0 - 0x0 -- plane 1
      12'h469: dout  = 8'b00000000; // 1129 :   0 - 0x0
      12'h46A: dout  = 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout  = 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout  = 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout  = 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout  = 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Background 0x47
      12'h471: dout  = 8'b00000000; // 1137 :   0 - 0x0
      12'h472: dout  = 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout  = 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout  = 8'b00000000; // 1140 :   0 - 0x0
      12'h475: dout  = 8'b00000000; // 1141 :   0 - 0x0
      12'h476: dout  = 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout  = 8'b00000000; // 1144 :   0 - 0x0 -- plane 1
      12'h479: dout  = 8'b00000000; // 1145 :   0 - 0x0
      12'h47A: dout  = 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout  = 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout  = 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Background 0x48
      12'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout  = 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout  = 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout  = 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout  = 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout  = 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout  = 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Background 0x49
      12'h491: dout  = 8'b00000000; // 1169 :   0 - 0x0
      12'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout  = 8'b00000000; // 1171 :   0 - 0x0
      12'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout  = 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout  = 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout  = 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout  = 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout  = 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Background 0x4a
      12'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout  = 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout  = 8'b00000000; // 1188 :   0 - 0x0
      12'h4A5: dout  = 8'b00000000; // 1189 :   0 - 0x0
      12'h4A6: dout  = 8'b00000000; // 1190 :   0 - 0x0
      12'h4A7: dout  = 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout  = 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout  = 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout  = 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout  = 8'b00000000; // 1195 :   0 - 0x0
      12'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Background 0x4b
      12'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout  = 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout  = 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout  = 8'b00000000; // 1204 :   0 - 0x0
      12'h4B5: dout  = 8'b00000000; // 1205 :   0 - 0x0
      12'h4B6: dout  = 8'b00000000; // 1206 :   0 - 0x0
      12'h4B7: dout  = 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout  = 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout  = 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout  = 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout  = 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Background 0x4c
      12'h4C1: dout  = 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      12'h4C6: dout  = 8'b00000000; // 1222 :   0 - 0x0
      12'h4C7: dout  = 8'b00000000; // 1223 :   0 - 0x0
      12'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout  = 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout  = 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout  = 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x4d
      12'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      12'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout  = 8'b00000000; // 1235 :   0 - 0x0
      12'h4D4: dout  = 8'b00000000; // 1236 :   0 - 0x0
      12'h4D5: dout  = 8'b00000000; // 1237 :   0 - 0x0
      12'h4D6: dout  = 8'b00000000; // 1238 :   0 - 0x0
      12'h4D7: dout  = 8'b00000000; // 1239 :   0 - 0x0
      12'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Background 0x4e
      12'h4E1: dout  = 8'b00000000; // 1249 :   0 - 0x0
      12'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      12'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      12'h4E4: dout  = 8'b00000000; // 1252 :   0 - 0x0
      12'h4E5: dout  = 8'b00000000; // 1253 :   0 - 0x0
      12'h4E6: dout  = 8'b00000000; // 1254 :   0 - 0x0
      12'h4E7: dout  = 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout  = 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout  = 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout  = 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout  = 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Background 0x4f
      12'h4F1: dout  = 8'b00000000; // 1265 :   0 - 0x0
      12'h4F2: dout  = 8'b00000000; // 1266 :   0 - 0x0
      12'h4F3: dout  = 8'b00000000; // 1267 :   0 - 0x0
      12'h4F4: dout  = 8'b00000000; // 1268 :   0 - 0x0
      12'h4F5: dout  = 8'b00000000; // 1269 :   0 - 0x0
      12'h4F6: dout  = 8'b00000000; // 1270 :   0 - 0x0
      12'h4F7: dout  = 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Background 0x50
      12'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      12'h503: dout  = 8'b00000000; // 1283 :   0 - 0x0
      12'h504: dout  = 8'b00000000; // 1284 :   0 - 0x0
      12'h505: dout  = 8'b00000000; // 1285 :   0 - 0x0
      12'h506: dout  = 8'b00000000; // 1286 :   0 - 0x0
      12'h507: dout  = 8'b00000000; // 1287 :   0 - 0x0
      12'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout  = 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout  = 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout  = 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout  = 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Background 0x51
      12'h511: dout  = 8'b00000000; // 1297 :   0 - 0x0
      12'h512: dout  = 8'b00000000; // 1298 :   0 - 0x0
      12'h513: dout  = 8'b00000000; // 1299 :   0 - 0x0
      12'h514: dout  = 8'b00000000; // 1300 :   0 - 0x0
      12'h515: dout  = 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout  = 8'b00000000; // 1302 :   0 - 0x0
      12'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Background 0x52
      12'h521: dout  = 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout  = 8'b00000000; // 1314 :   0 - 0x0
      12'h523: dout  = 8'b00000000; // 1315 :   0 - 0x0
      12'h524: dout  = 8'b00000000; // 1316 :   0 - 0x0
      12'h525: dout  = 8'b00000000; // 1317 :   0 - 0x0
      12'h526: dout  = 8'b00000000; // 1318 :   0 - 0x0
      12'h527: dout  = 8'b00000000; // 1319 :   0 - 0x0
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout  = 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout  = 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout  = 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout  = 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Background 0x53
      12'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout  = 8'b00000000; // 1331 :   0 - 0x0
      12'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout  = 8'b00000000; // 1333 :   0 - 0x0
      12'h536: dout  = 8'b00000000; // 1334 :   0 - 0x0
      12'h537: dout  = 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout  = 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Background 0x54
      12'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout  = 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout  = 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout  = 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout  = 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout  = 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout  = 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout  = 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Background 0x55
      12'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout  = 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Background 0x56
      12'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout  = 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout  = 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout  = 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout  = 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout  = 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout  = 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Background 0x57
      12'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Background 0x58
      12'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout  = 8'b00000000; // 1410 :   0 - 0x0
      12'h583: dout  = 8'b00000000; // 1411 :   0 - 0x0
      12'h584: dout  = 8'b00000000; // 1412 :   0 - 0x0
      12'h585: dout  = 8'b00000000; // 1413 :   0 - 0x0
      12'h586: dout  = 8'b00000000; // 1414 :   0 - 0x0
      12'h587: dout  = 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout  = 8'b00000000; // 1417 :   0 - 0x0
      12'h58A: dout  = 8'b00000000; // 1418 :   0 - 0x0
      12'h58B: dout  = 8'b00000000; // 1419 :   0 - 0x0
      12'h58C: dout  = 8'b00000000; // 1420 :   0 - 0x0
      12'h58D: dout  = 8'b00000000; // 1421 :   0 - 0x0
      12'h58E: dout  = 8'b00000000; // 1422 :   0 - 0x0
      12'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Background 0x59
      12'h591: dout  = 8'b00000000; // 1425 :   0 - 0x0
      12'h592: dout  = 8'b00000000; // 1426 :   0 - 0x0
      12'h593: dout  = 8'b00000000; // 1427 :   0 - 0x0
      12'h594: dout  = 8'b00000000; // 1428 :   0 - 0x0
      12'h595: dout  = 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout  = 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout  = 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout  = 8'b00000000; // 1433 :   0 - 0x0
      12'h59A: dout  = 8'b00000000; // 1434 :   0 - 0x0
      12'h59B: dout  = 8'b00000000; // 1435 :   0 - 0x0
      12'h59C: dout  = 8'b00000000; // 1436 :   0 - 0x0
      12'h59D: dout  = 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout  = 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Background 0x5a
      12'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout  = 8'b00000000; // 1442 :   0 - 0x0
      12'h5A3: dout  = 8'b00000000; // 1443 :   0 - 0x0
      12'h5A4: dout  = 8'b00000000; // 1444 :   0 - 0x0
      12'h5A5: dout  = 8'b00000000; // 1445 :   0 - 0x0
      12'h5A6: dout  = 8'b00000000; // 1446 :   0 - 0x0
      12'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout  = 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout  = 8'b00000000; // 1450 :   0 - 0x0
      12'h5AB: dout  = 8'b00000000; // 1451 :   0 - 0x0
      12'h5AC: dout  = 8'b00000000; // 1452 :   0 - 0x0
      12'h5AD: dout  = 8'b00000000; // 1453 :   0 - 0x0
      12'h5AE: dout  = 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Background 0x5b
      12'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout  = 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout  = 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout  = 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout  = 8'b00000000; // 1461 :   0 - 0x0
      12'h5B6: dout  = 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout  = 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout  = 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout  = 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout  = 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout  = 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout  = 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Background 0x5c
      12'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      12'h5C2: dout  = 8'b00000000; // 1474 :   0 - 0x0
      12'h5C3: dout  = 8'b00000000; // 1475 :   0 - 0x0
      12'h5C4: dout  = 8'b00000000; // 1476 :   0 - 0x0
      12'h5C5: dout  = 8'b00000000; // 1477 :   0 - 0x0
      12'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout  = 8'b00000000; // 1482 :   0 - 0x0
      12'h5CB: dout  = 8'b00000000; // 1483 :   0 - 0x0
      12'h5CC: dout  = 8'b00000000; // 1484 :   0 - 0x0
      12'h5CD: dout  = 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout  = 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Background 0x5d
      12'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout  = 8'b00000000; // 1490 :   0 - 0x0
      12'h5D3: dout  = 8'b00000000; // 1491 :   0 - 0x0
      12'h5D4: dout  = 8'b00000000; // 1492 :   0 - 0x0
      12'h5D5: dout  = 8'b00000000; // 1493 :   0 - 0x0
      12'h5D6: dout  = 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Background 0x5e
      12'h5E1: dout  = 8'b00000000; // 1505 :   0 - 0x0
      12'h5E2: dout  = 8'b00000000; // 1506 :   0 - 0x0
      12'h5E3: dout  = 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout  = 8'b00000000; // 1508 :   0 - 0x0
      12'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      12'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout  = 8'b00000000; // 1514 :   0 - 0x0
      12'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout  = 8'b00000000; // 1516 :   0 - 0x0
      12'h5ED: dout  = 8'b00000000; // 1517 :   0 - 0x0
      12'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Background 0x5f
      12'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout  = 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout  = 8'b00000000; // 1523 :   0 - 0x0
      12'h5F4: dout  = 8'b00000000; // 1524 :   0 - 0x0
      12'h5F5: dout  = 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Background 0x60
      12'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout  = 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout  = 8'b00000000; // 1542 :   0 - 0x0
      12'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout  = 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout  = 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Background 0x61
      12'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout  = 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout  = 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout  = 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout  = 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout  = 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout  = 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Background 0x62
      12'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout  = 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout  = 8'b00000000; // 1578 :   0 - 0x0
      12'h62B: dout  = 8'b00000000; // 1579 :   0 - 0x0
      12'h62C: dout  = 8'b00000000; // 1580 :   0 - 0x0
      12'h62D: dout  = 8'b00000000; // 1581 :   0 - 0x0
      12'h62E: dout  = 8'b00000000; // 1582 :   0 - 0x0
      12'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Background 0x63
      12'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout  = 8'b00000000; // 1589 :   0 - 0x0
      12'h636: dout  = 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- plane 1
      12'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Background 0x64
      12'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout  = 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout  = 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout  = 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout  = 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout  = 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Background 0x65
      12'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout  = 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout  = 8'b00000000; // 1622 :   0 - 0x0
      12'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Background 0x66
      12'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout  = 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout  = 8'b00000000; // 1638 :   0 - 0x0
      12'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout  = 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout  = 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout  = 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout  = 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Background 0x67
      12'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      12'h676: dout  = 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Background 0x68
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout  = 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout  = 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout  = 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Background 0x69
      12'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout  = 8'b00000000; // 1685 :   0 - 0x0
      12'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout  = 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout  = 8'b00000000; // 1690 :   0 - 0x0
      12'h69B: dout  = 8'b00000000; // 1691 :   0 - 0x0
      12'h69C: dout  = 8'b00000000; // 1692 :   0 - 0x0
      12'h69D: dout  = 8'b00000000; // 1693 :   0 - 0x0
      12'h69E: dout  = 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Background 0x6a
      12'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout  = 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout  = 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout  = 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout  = 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Background 0x6b
      12'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      12'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0 -- plane 1
      12'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      12'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      12'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      12'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      12'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Background 0x6c
      12'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout  = 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout  = 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- plane 1
      12'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Background 0x6d
      12'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout  = 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout  = 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout  = 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout  = 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Background 0x6e
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout  = 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Background 0x6f
      12'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout  = 8'b00000000; // 1781 :   0 - 0x0
      12'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout  = 8'b00000000; // 1784 :   0 - 0x0 -- plane 1
      12'h6F9: dout  = 8'b00000000; // 1785 :   0 - 0x0
      12'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout  = 8'b00000000; // 1787 :   0 - 0x0
      12'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout  = 8'b00000000; // 1789 :   0 - 0x0
      12'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Background 0x70
      12'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Background 0x71
      12'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout  = 8'b00000000; // 1816 :   0 - 0x0 -- plane 1
      12'h719: dout  = 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout  = 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout  = 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Background 0x72
      12'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout  = 8'b00000000; // 1829 :   0 - 0x0
      12'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout  = 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout  = 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Background 0x73
      12'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout  = 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout  = 8'b00000000; // 1845 :   0 - 0x0
      12'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- plane 1
      12'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Background 0x74
      12'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Background 0x75
      12'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- plane 1
      12'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Background 0x76
      12'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0 -- plane 1
      12'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Background 0x77
      12'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- plane 1
      12'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Background 0x78
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Background 0x79
      12'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0 -- plane 1
      12'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Background 0x7a
      12'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout  = 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout  = 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0 -- plane 1
      12'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Background 0x7b
      12'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- plane 1
      12'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Background 0x7c
      12'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Background 0x7d
      12'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Background 0x7e
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- plane 1
      12'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Background 0x7f
      12'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- plane 1
      12'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      12'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
      12'h800: dout  = 8'b10111111; // 2048 : 191 - 0xbf -- Background 0x80
      12'h801: dout  = 8'b11110111; // 2049 : 247 - 0xf7
      12'h802: dout  = 8'b11111101; // 2050 : 253 - 0xfd
      12'h803: dout  = 8'b11011111; // 2051 : 223 - 0xdf
      12'h804: dout  = 8'b11111011; // 2052 : 251 - 0xfb
      12'h805: dout  = 8'b10111111; // 2053 : 191 - 0xbf
      12'h806: dout  = 8'b11111110; // 2054 : 254 - 0xfe
      12'h807: dout  = 8'b11101111; // 2055 : 239 - 0xef
      12'h808: dout  = 8'b01000000; // 2056 :  64 - 0x40 -- plane 1
      12'h809: dout  = 8'b00001000; // 2057 :   8 - 0x8
      12'h80A: dout  = 8'b00000010; // 2058 :   2 - 0x2
      12'h80B: dout  = 8'b00100000; // 2059 :  32 - 0x20
      12'h80C: dout  = 8'b00000100; // 2060 :   4 - 0x4
      12'h80D: dout  = 8'b01000000; // 2061 :  64 - 0x40
      12'h80E: dout  = 8'b00000001; // 2062 :   1 - 0x1
      12'h80F: dout  = 8'b00010000; // 2063 :  16 - 0x10
      12'h810: dout  = 8'b11111111; // 2064 : 255 - 0xff -- Background 0x81
      12'h811: dout  = 8'b11101110; // 2065 : 238 - 0xee
      12'h812: dout  = 8'b11111111; // 2066 : 255 - 0xff
      12'h813: dout  = 8'b11011111; // 2067 : 223 - 0xdf
      12'h814: dout  = 8'b01110111; // 2068 : 119 - 0x77
      12'h815: dout  = 8'b11111101; // 2069 : 253 - 0xfd
      12'h816: dout  = 8'b11011111; // 2070 : 223 - 0xdf
      12'h817: dout  = 8'b10111111; // 2071 : 191 - 0xbf
      12'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout  = 8'b00010001; // 2073 :  17 - 0x11
      12'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout  = 8'b00100000; // 2075 :  32 - 0x20
      12'h81C: dout  = 8'b10001000; // 2076 : 136 - 0x88
      12'h81D: dout  = 8'b00000010; // 2077 :   2 - 0x2
      12'h81E: dout  = 8'b00100000; // 2078 :  32 - 0x20
      12'h81F: dout  = 8'b01000000; // 2079 :  64 - 0x40
      12'h820: dout  = 8'b11111110; // 2080 : 254 - 0xfe -- Background 0x82
      12'h821: dout  = 8'b11101111; // 2081 : 239 - 0xef
      12'h822: dout  = 8'b10111111; // 2082 : 191 - 0xbf
      12'h823: dout  = 8'b11110111; // 2083 : 247 - 0xf7
      12'h824: dout  = 8'b11111101; // 2084 : 253 - 0xfd
      12'h825: dout  = 8'b11011111; // 2085 : 223 - 0xdf
      12'h826: dout  = 8'b11111011; // 2086 : 251 - 0xfb
      12'h827: dout  = 8'b10111111; // 2087 : 191 - 0xbf
      12'h828: dout  = 8'b00000001; // 2088 :   1 - 0x1 -- plane 1
      12'h829: dout  = 8'b00010000; // 2089 :  16 - 0x10
      12'h82A: dout  = 8'b01000000; // 2090 :  64 - 0x40
      12'h82B: dout  = 8'b00001000; // 2091 :   8 - 0x8
      12'h82C: dout  = 8'b00000010; // 2092 :   2 - 0x2
      12'h82D: dout  = 8'b00100000; // 2093 :  32 - 0x20
      12'h82E: dout  = 8'b00000100; // 2094 :   4 - 0x4
      12'h82F: dout  = 8'b01000000; // 2095 :  64 - 0x40
      12'h830: dout  = 8'b11101111; // 2096 : 239 - 0xef -- Background 0x83
      12'h831: dout  = 8'b11111111; // 2097 : 255 - 0xff
      12'h832: dout  = 8'b10111011; // 2098 : 187 - 0xbb
      12'h833: dout  = 8'b11111111; // 2099 : 255 - 0xff
      12'h834: dout  = 8'b11110111; // 2100 : 247 - 0xf7
      12'h835: dout  = 8'b11011101; // 2101 : 221 - 0xdd
      12'h836: dout  = 8'b01111111; // 2102 : 127 - 0x7f
      12'h837: dout  = 8'b11110111; // 2103 : 247 - 0xf7
      12'h838: dout  = 8'b00010000; // 2104 :  16 - 0x10 -- plane 1
      12'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout  = 8'b01000100; // 2106 :  68 - 0x44
      12'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout  = 8'b00001000; // 2108 :   8 - 0x8
      12'h83D: dout  = 8'b00100010; // 2109 :  34 - 0x22
      12'h83E: dout  = 8'b10000000; // 2110 : 128 - 0x80
      12'h83F: dout  = 8'b00001000; // 2111 :   8 - 0x8
      12'h840: dout  = 8'b11111111; // 2112 : 255 - 0xff -- Background 0x84
      12'h841: dout  = 8'b11101110; // 2113 : 238 - 0xee
      12'h842: dout  = 8'b11111011; // 2114 : 251 - 0xfb
      12'h843: dout  = 8'b10111111; // 2115 : 191 - 0xbf
      12'h844: dout  = 8'b01111111; // 2116 : 127 - 0x7f
      12'h845: dout  = 8'b11101101; // 2117 : 237 - 0xed
      12'h846: dout  = 8'b11111111; // 2118 : 255 - 0xff
      12'h847: dout  = 8'b10111111; // 2119 : 191 - 0xbf
      12'h848: dout  = 8'b00010100; // 2120 :  20 - 0x14 -- plane 1
      12'h849: dout  = 8'b10110101; // 2121 : 181 - 0xb5
      12'h84A: dout  = 8'b01000100; // 2122 :  68 - 0x44
      12'h84B: dout  = 8'b01001010; // 2123 :  74 - 0x4a
      12'h84C: dout  = 8'b10010010; // 2124 : 146 - 0x92
      12'h84D: dout  = 8'b10010010; // 2125 : 146 - 0x92
      12'h84E: dout  = 8'b01000100; // 2126 :  68 - 0x44
      12'h84F: dout  = 8'b01001001; // 2127 :  73 - 0x49
      12'h850: dout  = 8'b11111111; // 2128 : 255 - 0xff -- Background 0x85
      12'h851: dout  = 8'b10111111; // 2129 : 191 - 0xbf
      12'h852: dout  = 8'b01111101; // 2130 : 125 - 0x7d
      12'h853: dout  = 8'b11110111; // 2131 : 247 - 0xf7
      12'h854: dout  = 8'b11011011; // 2132 : 219 - 0xdb
      12'h855: dout  = 8'b11111101; // 2133 : 253 - 0xfd
      12'h856: dout  = 8'b01111110; // 2134 : 126 - 0x7e
      12'h857: dout  = 8'b11111011; // 2135 : 251 - 0xfb
      12'h858: dout  = 8'b01000010; // 2136 :  66 - 0x42 -- plane 1
      12'h859: dout  = 8'b01001010; // 2137 :  74 - 0x4a
      12'h85A: dout  = 8'b11001010; // 2138 : 202 - 0xca
      12'h85B: dout  = 8'b00101001; // 2139 :  41 - 0x29
      12'h85C: dout  = 8'b10100110; // 2140 : 166 - 0xa6
      12'h85D: dout  = 8'b10010010; // 2141 : 146 - 0x92
      12'h85E: dout  = 8'b10001001; // 2142 : 137 - 0x89
      12'h85F: dout  = 8'b00101101; // 2143 :  45 - 0x2d
      12'h860: dout  = 8'b11111111; // 2144 : 255 - 0xff -- Background 0x86
      12'h861: dout  = 8'b11110111; // 2145 : 247 - 0xf7
      12'h862: dout  = 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout  = 8'b11011101; // 2147 : 221 - 0xdd
      12'h864: dout  = 8'b01111111; // 2148 : 127 - 0x7f
      12'h865: dout  = 8'b11110111; // 2149 : 247 - 0xf7
      12'h866: dout  = 8'b11101111; // 2150 : 239 - 0xef
      12'h867: dout  = 8'b10111101; // 2151 : 189 - 0xbd
      12'h868: dout  = 8'b10001000; // 2152 : 136 - 0x88 -- plane 1
      12'h869: dout  = 8'b00101001; // 2153 :  41 - 0x29
      12'h86A: dout  = 8'b10000010; // 2154 : 130 - 0x82
      12'h86B: dout  = 8'b10110110; // 2155 : 182 - 0xb6
      12'h86C: dout  = 8'b10001000; // 2156 : 136 - 0x88
      12'h86D: dout  = 8'b01001001; // 2157 :  73 - 0x49
      12'h86E: dout  = 8'b01010010; // 2158 :  82 - 0x52
      12'h86F: dout  = 8'b01010010; // 2159 :  82 - 0x52
      12'h870: dout  = 8'b01011111; // 2160 :  95 - 0x5f -- Background 0x87
      12'h871: dout  = 8'b11111101; // 2161 : 253 - 0xfd
      12'h872: dout  = 8'b11110110; // 2162 : 246 - 0xf6
      12'h873: dout  = 8'b01111111; // 2163 : 127 - 0x7f
      12'h874: dout  = 8'b10011111; // 2164 : 159 - 0x9f
      12'h875: dout  = 8'b11111110; // 2165 : 254 - 0xfe
      12'h876: dout  = 8'b11111111; // 2166 : 255 - 0xff
      12'h877: dout  = 8'b11101111; // 2167 : 239 - 0xef
      12'h878: dout  = 8'b10110010; // 2168 : 178 - 0xb2 -- plane 1
      12'h879: dout  = 8'b01001010; // 2169 :  74 - 0x4a
      12'h87A: dout  = 8'b10101001; // 2170 : 169 - 0xa9
      12'h87B: dout  = 8'b10100100; // 2171 : 164 - 0xa4
      12'h87C: dout  = 8'b01100010; // 2172 :  98 - 0x62
      12'h87D: dout  = 8'b01001011; // 2173 :  75 - 0x4b
      12'h87E: dout  = 8'b10010000; // 2174 : 144 - 0x90
      12'h87F: dout  = 8'b10010010; // 2175 : 146 - 0x92
      12'h880: dout  = 8'b11111111; // 2176 : 255 - 0xff -- Background 0x88
      12'h881: dout  = 8'b10011111; // 2177 : 159 - 0x9f
      12'h882: dout  = 8'b10111111; // 2178 : 191 - 0xbf
      12'h883: dout  = 8'b11111111; // 2179 : 255 - 0xff
      12'h884: dout  = 8'b11110011; // 2180 : 243 - 0xf3
      12'h885: dout  = 8'b11110011; // 2181 : 243 - 0xf3
      12'h886: dout  = 8'b11111111; // 2182 : 255 - 0xff
      12'h887: dout  = 8'b11111111; // 2183 : 255 - 0xff
      12'h888: dout  = 8'b01100000; // 2184 :  96 - 0x60 -- plane 1
      12'h889: dout  = 8'b11110000; // 2185 : 240 - 0xf0
      12'h88A: dout  = 8'b11110000; // 2186 : 240 - 0xf0
      12'h88B: dout  = 8'b01101110; // 2187 : 110 - 0x6e
      12'h88C: dout  = 8'b00011111; // 2188 :  31 - 0x1f
      12'h88D: dout  = 8'b00011111; // 2189 :  31 - 0x1f
      12'h88E: dout  = 8'b00011111; // 2190 :  31 - 0x1f
      12'h88F: dout  = 8'b00001110; // 2191 :  14 - 0xe
      12'h890: dout  = 8'b11111111; // 2192 : 255 - 0xff -- Background 0x89
      12'h891: dout  = 8'b10011111; // 2193 : 159 - 0x9f
      12'h892: dout  = 8'b10111111; // 2194 : 191 - 0xbf
      12'h893: dout  = 8'b11110011; // 2195 : 243 - 0xf3
      12'h894: dout  = 8'b11110011; // 2196 : 243 - 0xf3
      12'h895: dout  = 8'b11111111; // 2197 : 255 - 0xff
      12'h896: dout  = 8'b11111111; // 2198 : 255 - 0xff
      12'h897: dout  = 8'b11111111; // 2199 : 255 - 0xff
      12'h898: dout  = 8'b01100000; // 2200 :  96 - 0x60 -- plane 1
      12'h899: dout  = 8'b11110000; // 2201 : 240 - 0xf0
      12'h89A: dout  = 8'b11111110; // 2202 : 254 - 0xfe
      12'h89B: dout  = 8'b01111111; // 2203 : 127 - 0x7f
      12'h89C: dout  = 8'b00011111; // 2204 :  31 - 0x1f
      12'h89D: dout  = 8'b00011111; // 2205 :  31 - 0x1f
      12'h89E: dout  = 8'b00001110; // 2206 :  14 - 0xe
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b10111111; // 2208 : 191 - 0xbf -- Background 0x8a
      12'h8A1: dout  = 8'b11110111; // 2209 : 247 - 0xf7
      12'h8A2: dout  = 8'b11111101; // 2210 : 253 - 0xfd
      12'h8A3: dout  = 8'b11111111; // 2211 : 255 - 0xff
      12'h8A4: dout  = 8'b11111011; // 2212 : 251 - 0xfb
      12'h8A5: dout  = 8'b10111111; // 2213 : 191 - 0xbf
      12'h8A6: dout  = 8'b11111110; // 2214 : 254 - 0xfe
      12'h8A7: dout  = 8'b11101111; // 2215 : 239 - 0xef
      12'h8A8: dout  = 8'b01000000; // 2216 :  64 - 0x40 -- plane 1
      12'h8A9: dout  = 8'b00001000; // 2217 :   8 - 0x8
      12'h8AA: dout  = 8'b00000010; // 2218 :   2 - 0x2
      12'h8AB: dout  = 8'b00101000; // 2219 :  40 - 0x28
      12'h8AC: dout  = 8'b00010100; // 2220 :  20 - 0x14
      12'h8AD: dout  = 8'b01010100; // 2221 :  84 - 0x54
      12'h8AE: dout  = 8'b00000001; // 2222 :   1 - 0x1
      12'h8AF: dout  = 8'b00010000; // 2223 :  16 - 0x10
      12'h8B0: dout  = 8'b10111111; // 2224 : 191 - 0xbf -- Background 0x8b
      12'h8B1: dout  = 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout  = 8'b11101110; // 2226 : 238 - 0xee
      12'h8B3: dout  = 8'b11111111; // 2227 : 255 - 0xff
      12'h8B4: dout  = 8'b11011111; // 2228 : 223 - 0xdf
      12'h8B5: dout  = 8'b01111101; // 2229 : 125 - 0x7d
      12'h8B6: dout  = 8'b11111111; // 2230 : 255 - 0xff
      12'h8B7: dout  = 8'b11011111; // 2231 : 223 - 0xdf
      12'h8B8: dout  = 8'b01000000; // 2232 :  64 - 0x40 -- plane 1
      12'h8B9: dout  = 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout  = 8'b10010001; // 2234 : 145 - 0x91
      12'h8BB: dout  = 8'b00010100; // 2235 :  20 - 0x14
      12'h8BC: dout  = 8'b00101000; // 2236 :  40 - 0x28
      12'h8BD: dout  = 8'b10001010; // 2237 : 138 - 0x8a
      12'h8BE: dout  = 8'b01000000; // 2238 :  64 - 0x40
      12'h8BF: dout  = 8'b00100000; // 2239 :  32 - 0x20
      12'h8C0: dout  = 8'b11111111; // 2240 : 255 - 0xff -- Background 0x8c
      12'h8C1: dout  = 8'b11111000; // 2241 : 248 - 0xf8
      12'h8C2: dout  = 8'b11100010; // 2242 : 226 - 0xe2
      12'h8C3: dout  = 8'b11010111; // 2243 : 215 - 0xd7
      12'h8C4: dout  = 8'b11001111; // 2244 : 207 - 0xcf
      12'h8C5: dout  = 8'b10011111; // 2245 : 159 - 0x9f
      12'h8C6: dout  = 8'b10111110; // 2246 : 190 - 0xbe
      12'h8C7: dout  = 8'b10011101; // 2247 : 157 - 0x9d
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout  = 8'b00000111; // 2249 :   7 - 0x7
      12'h8CA: dout  = 8'b00011111; // 2250 :  31 - 0x1f
      12'h8CB: dout  = 8'b00111111; // 2251 :  63 - 0x3f
      12'h8CC: dout  = 8'b00111111; // 2252 :  63 - 0x3f
      12'h8CD: dout  = 8'b01111111; // 2253 : 127 - 0x7f
      12'h8CE: dout  = 8'b01111111; // 2254 : 127 - 0x7f
      12'h8CF: dout  = 8'b01111111; // 2255 : 127 - 0x7f
      12'h8D0: dout  = 8'b11111111; // 2256 : 255 - 0xff -- Background 0x8d
      12'h8D1: dout  = 8'b00011111; // 2257 :  31 - 0x1f
      12'h8D2: dout  = 8'b10100111; // 2258 : 167 - 0xa7
      12'h8D3: dout  = 8'b11000011; // 2259 : 195 - 0xc3
      12'h8D4: dout  = 8'b11100011; // 2260 : 227 - 0xe3
      12'h8D5: dout  = 8'b01000001; // 2261 :  65 - 0x41
      12'h8D6: dout  = 8'b10100001; // 2262 : 161 - 0xa1
      12'h8D7: dout  = 8'b00000001; // 2263 :   1 - 0x1
      12'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0 -- plane 1
      12'h8D9: dout  = 8'b11100000; // 2265 : 224 - 0xe0
      12'h8DA: dout  = 8'b11111000; // 2266 : 248 - 0xf8
      12'h8DB: dout  = 8'b11111000; // 2267 : 248 - 0xf8
      12'h8DC: dout  = 8'b11110000; // 2268 : 240 - 0xf0
      12'h8DD: dout  = 8'b11111000; // 2269 : 248 - 0xf8
      12'h8DE: dout  = 8'b11110100; // 2270 : 244 - 0xf4
      12'h8DF: dout  = 8'b11111000; // 2271 : 248 - 0xf8
      12'h8E0: dout  = 8'b10111110; // 2272 : 190 - 0xbe -- Background 0x8e
      12'h8E1: dout  = 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout  = 8'b11011111; // 2274 : 223 - 0xdf
      12'h8E3: dout  = 8'b11111111; // 2275 : 255 - 0xff
      12'h8E4: dout  = 8'b11101111; // 2276 : 239 - 0xef
      12'h8E5: dout  = 8'b11111111; // 2277 : 255 - 0xff
      12'h8E6: dout  = 8'b11110111; // 2278 : 247 - 0xf7
      12'h8E7: dout  = 8'b11111111; // 2279 : 255 - 0xff
      12'h8E8: dout  = 8'b01111111; // 2280 : 127 - 0x7f -- plane 1
      12'h8E9: dout  = 8'b00111111; // 2281 :  63 - 0x3f
      12'h8EA: dout  = 8'b00111111; // 2282 :  63 - 0x3f
      12'h8EB: dout  = 8'b00011111; // 2283 :  31 - 0x1f
      12'h8EC: dout  = 8'b00011111; // 2284 :  31 - 0x1f
      12'h8ED: dout  = 8'b00001111; // 2285 :  15 - 0xf
      12'h8EE: dout  = 8'b00001111; // 2286 :  15 - 0xf
      12'h8EF: dout  = 8'b00000111; // 2287 :   7 - 0x7
      12'h8F0: dout  = 8'b01111101; // 2288 : 125 - 0x7d -- Background 0x8f
      12'h8F1: dout  = 8'b11111111; // 2289 : 255 - 0xff
      12'h8F2: dout  = 8'b11111011; // 2290 : 251 - 0xfb
      12'h8F3: dout  = 8'b11111111; // 2291 : 255 - 0xff
      12'h8F4: dout  = 8'b11110111; // 2292 : 247 - 0xf7
      12'h8F5: dout  = 8'b11111111; // 2293 : 255 - 0xff
      12'h8F6: dout  = 8'b11101111; // 2294 : 239 - 0xef
      12'h8F7: dout  = 8'b11111111; // 2295 : 255 - 0xff
      12'h8F8: dout  = 8'b11111110; // 2296 : 254 - 0xfe -- plane 1
      12'h8F9: dout  = 8'b11111100; // 2297 : 252 - 0xfc
      12'h8FA: dout  = 8'b11111100; // 2298 : 252 - 0xfc
      12'h8FB: dout  = 8'b11111000; // 2299 : 248 - 0xf8
      12'h8FC: dout  = 8'b11111000; // 2300 : 248 - 0xf8
      12'h8FD: dout  = 8'b11110000; // 2301 : 240 - 0xf0
      12'h8FE: dout  = 8'b11110000; // 2302 : 240 - 0xf0
      12'h8FF: dout  = 8'b11100000; // 2303 : 224 - 0xe0
      12'h900: dout  = 8'b10111110; // 2304 : 190 - 0xbe -- Background 0x90
      12'h901: dout  = 8'b11110111; // 2305 : 247 - 0xf7
      12'h902: dout  = 8'b11111111; // 2306 : 255 - 0xff
      12'h903: dout  = 8'b11011111; // 2307 : 223 - 0xdf
      12'h904: dout  = 8'b11111011; // 2308 : 251 - 0xfb
      12'h905: dout  = 8'b11111110; // 2309 : 254 - 0xfe
      12'h906: dout  = 8'b10111111; // 2310 : 191 - 0xbf
      12'h907: dout  = 8'b11110111; // 2311 : 247 - 0xf7
      12'h908: dout  = 8'b01000001; // 2312 :  65 - 0x41 -- plane 1
      12'h909: dout  = 8'b00001000; // 2313 :   8 - 0x8
      12'h90A: dout  = 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout  = 8'b00100000; // 2315 :  32 - 0x20
      12'h90C: dout  = 8'b00000100; // 2316 :   4 - 0x4
      12'h90D: dout  = 8'b00000001; // 2317 :   1 - 0x1
      12'h90E: dout  = 8'b01000000; // 2318 :  64 - 0x40
      12'h90F: dout  = 8'b00001000; // 2319 :   8 - 0x8
      12'h910: dout  = 8'b11101110; // 2320 : 238 - 0xee -- Background 0x91
      12'h911: dout  = 8'b11111111; // 2321 : 255 - 0xff
      12'h912: dout  = 8'b01111011; // 2322 : 123 - 0x7b
      12'h913: dout  = 8'b11111101; // 2323 : 253 - 0xfd
      12'h914: dout  = 8'b11101111; // 2324 : 239 - 0xef
      12'h915: dout  = 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout  = 8'b10111101; // 2326 : 189 - 0xbd
      12'h917: dout  = 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout  = 8'b00010001; // 2328 :  17 - 0x11 -- plane 1
      12'h919: dout  = 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout  = 8'b10000100; // 2330 : 132 - 0x84
      12'h91B: dout  = 8'b00000010; // 2331 :   2 - 0x2
      12'h91C: dout  = 8'b00010000; // 2332 :  16 - 0x10
      12'h91D: dout  = 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout  = 8'b01000010; // 2334 :  66 - 0x42
      12'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout  = 8'b11111011; // 2336 : 251 - 0xfb -- Background 0x92
      12'h921: dout  = 8'b10111111; // 2337 : 191 - 0xbf
      12'h922: dout  = 8'b11101111; // 2338 : 239 - 0xef
      12'h923: dout  = 8'b11111101; // 2339 : 253 - 0xfd
      12'h924: dout  = 8'b11111111; // 2340 : 255 - 0xff
      12'h925: dout  = 8'b10111111; // 2341 : 191 - 0xbf
      12'h926: dout  = 8'b11111011; // 2342 : 251 - 0xfb
      12'h927: dout  = 8'b11011111; // 2343 : 223 - 0xdf
      12'h928: dout  = 8'b00000100; // 2344 :   4 - 0x4 -- plane 1
      12'h929: dout  = 8'b01000000; // 2345 :  64 - 0x40
      12'h92A: dout  = 8'b00010000; // 2346 :  16 - 0x10
      12'h92B: dout  = 8'b00000010; // 2347 :   2 - 0x2
      12'h92C: dout  = 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout  = 8'b01000000; // 2349 :  64 - 0x40
      12'h92E: dout  = 8'b00000100; // 2350 :   4 - 0x4
      12'h92F: dout  = 8'b00100000; // 2351 :  32 - 0x20
      12'h930: dout  = 8'b10111101; // 2352 : 189 - 0xbd -- Background 0x93
      12'h931: dout  = 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout  = 8'b01110111; // 2354 : 119 - 0x77
      12'h933: dout  = 8'b11111110; // 2355 : 254 - 0xfe
      12'h934: dout  = 8'b11011111; // 2356 : 223 - 0xdf
      12'h935: dout  = 8'b11111011; // 2357 : 251 - 0xfb
      12'h936: dout  = 8'b11101111; // 2358 : 239 - 0xef
      12'h937: dout  = 8'b01111111; // 2359 : 127 - 0x7f
      12'h938: dout  = 8'b01000010; // 2360 :  66 - 0x42 -- plane 1
      12'h939: dout  = 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout  = 8'b10001000; // 2362 : 136 - 0x88
      12'h93B: dout  = 8'b00000001; // 2363 :   1 - 0x1
      12'h93C: dout  = 8'b00100000; // 2364 :  32 - 0x20
      12'h93D: dout  = 8'b00000100; // 2365 :   4 - 0x4
      12'h93E: dout  = 8'b00010000; // 2366 :  16 - 0x10
      12'h93F: dout  = 8'b10000000; // 2367 : 128 - 0x80
      12'h940: dout  = 8'b01111111; // 2368 : 127 - 0x7f -- Background 0x94
      12'h941: dout  = 8'b11110111; // 2369 : 247 - 0xf7
      12'h942: dout  = 8'b11011101; // 2370 : 221 - 0xdd
      12'h943: dout  = 8'b01111011; // 2371 : 123 - 0x7b
      12'h944: dout  = 8'b11111111; // 2372 : 255 - 0xff
      12'h945: dout  = 8'b11101110; // 2373 : 238 - 0xee
      12'h946: dout  = 8'b10111011; // 2374 : 187 - 0xbb
      12'h947: dout  = 8'b11111101; // 2375 : 253 - 0xfd
      12'h948: dout  = 8'b11001000; // 2376 : 200 - 0xc8 -- plane 1
      12'h949: dout  = 8'b00101010; // 2377 :  42 - 0x2a
      12'h94A: dout  = 8'b10100010; // 2378 : 162 - 0xa2
      12'h94B: dout  = 8'b10010100; // 2379 : 148 - 0x94
      12'h94C: dout  = 8'b10010001; // 2380 : 145 - 0x91
      12'h94D: dout  = 8'b01010101; // 2381 :  85 - 0x55
      12'h94E: dout  = 8'b01000100; // 2382 :  68 - 0x44
      12'h94F: dout  = 8'b00010010; // 2383 :  18 - 0x12
      12'h950: dout  = 8'b11010111; // 2384 : 215 - 0xd7 -- Background 0x95
      12'h951: dout  = 8'b01111111; // 2385 : 127 - 0x7f
      12'h952: dout  = 8'b11111101; // 2386 : 253 - 0xfd
      12'h953: dout  = 8'b11101110; // 2387 : 238 - 0xee
      12'h954: dout  = 8'b11110111; // 2388 : 247 - 0xf7
      12'h955: dout  = 8'b10111011; // 2389 : 187 - 0xbb
      12'h956: dout  = 8'b11101111; // 2390 : 239 - 0xef
      12'h957: dout  = 8'b11110111; // 2391 : 247 - 0xf7
      12'h958: dout  = 8'b10101010; // 2392 : 170 - 0xaa -- plane 1
      12'h959: dout  = 8'b10100010; // 2393 : 162 - 0xa2
      12'h95A: dout  = 8'b00010010; // 2394 :  18 - 0x12
      12'h95B: dout  = 8'b01010011; // 2395 :  83 - 0x53
      12'h95C: dout  = 8'b01001100; // 2396 :  76 - 0x4c
      12'h95D: dout  = 8'b01010101; // 2397 :  85 - 0x55
      12'h95E: dout  = 8'b10010001; // 2398 : 145 - 0x91
      12'h95F: dout  = 8'b01001000; // 2399 :  72 - 0x48
      12'h960: dout  = 8'b10111111; // 2400 : 191 - 0xbf -- Background 0x96
      12'h961: dout  = 8'b11101110; // 2401 : 238 - 0xee
      12'h962: dout  = 8'b11011011; // 2402 : 219 - 0xdb
      12'h963: dout  = 8'b11111111; // 2403 : 255 - 0xff
      12'h964: dout  = 8'b01110111; // 2404 : 119 - 0x77
      12'h965: dout  = 8'b11011101; // 2405 : 221 - 0xdd
      12'h966: dout  = 8'b11101111; // 2406 : 239 - 0xef
      12'h967: dout  = 8'b11111011; // 2407 : 251 - 0xfb
      12'h968: dout  = 8'b01010001; // 2408 :  81 - 0x51 -- plane 1
      12'h969: dout  = 8'b00010101; // 2409 :  21 - 0x15
      12'h96A: dout  = 8'b10100100; // 2410 : 164 - 0xa4
      12'h96B: dout  = 8'b10001100; // 2411 : 140 - 0x8c
      12'h96C: dout  = 8'b10101010; // 2412 : 170 - 0xaa
      12'h96D: dout  = 8'b00100010; // 2413 :  34 - 0x22
      12'h96E: dout  = 8'b10010000; // 2414 : 144 - 0x90
      12'h96F: dout  = 8'b01000110; // 2415 :  70 - 0x46
      12'h970: dout  = 8'b11111101; // 2416 : 253 - 0xfd -- Background 0x97
      12'h971: dout  = 8'b11101110; // 2417 : 238 - 0xee
      12'h972: dout  = 8'b11111011; // 2418 : 251 - 0xfb
      12'h973: dout  = 8'b11111101; // 2419 : 253 - 0xfd
      12'h974: dout  = 8'b11110101; // 2420 : 245 - 0xf5
      12'h975: dout  = 8'b11011111; // 2421 : 223 - 0xdf
      12'h976: dout  = 8'b01111111; // 2422 : 127 - 0x7f
      12'h977: dout  = 8'b10111011; // 2423 : 187 - 0xbb
      12'h978: dout  = 8'b00010011; // 2424 :  19 - 0x13 -- plane 1
      12'h979: dout  = 8'b01010101; // 2425 :  85 - 0x55
      12'h97A: dout  = 8'b01100100; // 2426 : 100 - 0x64
      12'h97B: dout  = 8'b00010010; // 2427 :  18 - 0x12
      12'h97C: dout  = 8'b10101010; // 2428 : 170 - 0xaa
      12'h97D: dout  = 8'b10101000; // 2429 : 168 - 0xa8
      12'h97E: dout  = 8'b10000100; // 2430 : 132 - 0x84
      12'h97F: dout  = 8'b11010100; // 2431 : 212 - 0xd4
      12'h980: dout  = 8'b11111111; // 2432 : 255 - 0xff -- Background 0x98
      12'h981: dout  = 8'b10011111; // 2433 : 159 - 0x9f
      12'h982: dout  = 8'b10111111; // 2434 : 191 - 0xbf
      12'h983: dout  = 8'b11110011; // 2435 : 243 - 0xf3
      12'h984: dout  = 8'b11110011; // 2436 : 243 - 0xf3
      12'h985: dout  = 8'b11111111; // 2437 : 255 - 0xff
      12'h986: dout  = 8'b11111111; // 2438 : 255 - 0xff
      12'h987: dout  = 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout  = 8'b01100000; // 2440 :  96 - 0x60 -- plane 1
      12'h989: dout  = 8'b11110000; // 2441 : 240 - 0xf0
      12'h98A: dout  = 8'b11111110; // 2442 : 254 - 0xfe
      12'h98B: dout  = 8'b01111111; // 2443 : 127 - 0x7f
      12'h98C: dout  = 8'b00011111; // 2444 :  31 - 0x1f
      12'h98D: dout  = 8'b00011111; // 2445 :  31 - 0x1f
      12'h98E: dout  = 8'b00001110; // 2446 :  14 - 0xe
      12'h98F: dout  = 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout  = 8'b11111111; // 2448 : 255 - 0xff -- Background 0x99
      12'h991: dout  = 8'b10011111; // 2449 : 159 - 0x9f
      12'h992: dout  = 8'b10111111; // 2450 : 191 - 0xbf
      12'h993: dout  = 8'b11111111; // 2451 : 255 - 0xff
      12'h994: dout  = 8'b11110011; // 2452 : 243 - 0xf3
      12'h995: dout  = 8'b11110011; // 2453 : 243 - 0xf3
      12'h996: dout  = 8'b11111111; // 2454 : 255 - 0xff
      12'h997: dout  = 8'b11111111; // 2455 : 255 - 0xff
      12'h998: dout  = 8'b01100000; // 2456 :  96 - 0x60 -- plane 1
      12'h999: dout  = 8'b11110000; // 2457 : 240 - 0xf0
      12'h99A: dout  = 8'b11110000; // 2458 : 240 - 0xf0
      12'h99B: dout  = 8'b01101110; // 2459 : 110 - 0x6e
      12'h99C: dout  = 8'b00011111; // 2460 :  31 - 0x1f
      12'h99D: dout  = 8'b00011111; // 2461 :  31 - 0x1f
      12'h99E: dout  = 8'b00011111; // 2462 :  31 - 0x1f
      12'h99F: dout  = 8'b00001110; // 2463 :  14 - 0xe
      12'h9A0: dout  = 8'b10111111; // 2464 : 191 - 0xbf -- Background 0x9a
      12'h9A1: dout  = 8'b11110111; // 2465 : 247 - 0xf7
      12'h9A2: dout  = 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout  = 8'b11011111; // 2467 : 223 - 0xdf
      12'h9A4: dout  = 8'b11111011; // 2468 : 251 - 0xfb
      12'h9A5: dout  = 8'b11111111; // 2469 : 255 - 0xff
      12'h9A6: dout  = 8'b10111111; // 2470 : 191 - 0xbf
      12'h9A7: dout  = 8'b11110111; // 2471 : 247 - 0xf7
      12'h9A8: dout  = 8'b01000000; // 2472 :  64 - 0x40 -- plane 1
      12'h9A9: dout  = 8'b00001100; // 2473 :  12 - 0xc
      12'h9AA: dout  = 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout  = 8'b00101000; // 2475 :  40 - 0x28
      12'h9AC: dout  = 8'b00101100; // 2476 :  44 - 0x2c
      12'h9AD: dout  = 8'b00010001; // 2477 :  17 - 0x11
      12'h9AE: dout  = 8'b01000000; // 2478 :  64 - 0x40
      12'h9AF: dout  = 8'b00001000; // 2479 :   8 - 0x8
      12'h9B0: dout  = 8'b11011111; // 2480 : 223 - 0xdf -- Background 0x9b
      12'h9B1: dout  = 8'b11111111; // 2481 : 255 - 0xff
      12'h9B2: dout  = 8'b01111011; // 2482 : 123 - 0x7b
      12'h9B3: dout  = 8'b11111111; // 2483 : 255 - 0xff
      12'h9B4: dout  = 8'b11101111; // 2484 : 239 - 0xef
      12'h9B5: dout  = 8'b11111101; // 2485 : 253 - 0xfd
      12'h9B6: dout  = 8'b10111111; // 2486 : 191 - 0xbf
      12'h9B7: dout  = 8'b11111111; // 2487 : 255 - 0xff
      12'h9B8: dout  = 8'b00100000; // 2488 :  32 - 0x20 -- plane 1
      12'h9B9: dout  = 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout  = 8'b10010100; // 2490 : 148 - 0x94
      12'h9BB: dout  = 8'b01001000; // 2491 :  72 - 0x48
      12'h9BC: dout  = 8'b00011000; // 2492 :  24 - 0x18
      12'h9BD: dout  = 8'b00000110; // 2493 :   6 - 0x6
      12'h9BE: dout  = 8'b01000000; // 2494 :  64 - 0x40
      12'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout  = 8'b10111010; // 2496 : 186 - 0xba -- Background 0x9c
      12'h9C1: dout  = 8'b10011100; // 2497 : 156 - 0x9c
      12'h9C2: dout  = 8'b10101010; // 2498 : 170 - 0xaa
      12'h9C3: dout  = 8'b11000000; // 2499 : 192 - 0xc0
      12'h9C4: dout  = 8'b11000000; // 2500 : 192 - 0xc0
      12'h9C5: dout  = 8'b11100000; // 2501 : 224 - 0xe0
      12'h9C6: dout  = 8'b11111000; // 2502 : 248 - 0xf8
      12'h9C7: dout  = 8'b11111111; // 2503 : 255 - 0xff
      12'h9C8: dout  = 8'b01111111; // 2504 : 127 - 0x7f -- plane 1
      12'h9C9: dout  = 8'b01111111; // 2505 : 127 - 0x7f
      12'h9CA: dout  = 8'b01111111; // 2506 : 127 - 0x7f
      12'h9CB: dout  = 8'b00111111; // 2507 :  63 - 0x3f
      12'h9CC: dout  = 8'b00110101; // 2508 :  53 - 0x35
      12'h9CD: dout  = 8'b00000010; // 2509 :   2 - 0x2
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b00000001; // 2512 :   1 - 0x1 -- Background 0x9d
      12'h9D1: dout  = 8'b00000001; // 2513 :   1 - 0x1
      12'h9D2: dout  = 8'b00000001; // 2514 :   1 - 0x1
      12'h9D3: dout  = 8'b00000011; // 2515 :   3 - 0x3
      12'h9D4: dout  = 8'b00000011; // 2516 :   3 - 0x3
      12'h9D5: dout  = 8'b00000111; // 2517 :   7 - 0x7
      12'h9D6: dout  = 8'b00011111; // 2518 :  31 - 0x1f
      12'h9D7: dout  = 8'b11111111; // 2519 : 255 - 0xff
      12'h9D8: dout  = 8'b11110100; // 2520 : 244 - 0xf4 -- plane 1
      12'h9D9: dout  = 8'b11111000; // 2521 : 248 - 0xf8
      12'h9DA: dout  = 8'b11110000; // 2522 : 240 - 0xf0
      12'h9DB: dout  = 8'b11101000; // 2523 : 232 - 0xe8
      12'h9DC: dout  = 8'b01010000; // 2524 :  80 - 0x50
      12'h9DD: dout  = 8'b10000000; // 2525 : 128 - 0x80
      12'h9DE: dout  = 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout  = 8'b01111101; // 2528 : 125 - 0x7d -- Background 0x9e
      12'h9E1: dout  = 8'b11111111; // 2529 : 255 - 0xff
      12'h9E2: dout  = 8'b11111011; // 2530 : 251 - 0xfb
      12'h9E3: dout  = 8'b11111111; // 2531 : 255 - 0xff
      12'h9E4: dout  = 8'b11111111; // 2532 : 255 - 0xff
      12'h9E5: dout  = 8'b11111011; // 2533 : 251 - 0xfb
      12'h9E6: dout  = 8'b11111111; // 2534 : 255 - 0xff
      12'h9E7: dout  = 8'b01111101; // 2535 : 125 - 0x7d
      12'h9E8: dout  = 8'b11111110; // 2536 : 254 - 0xfe -- plane 1
      12'h9E9: dout  = 8'b11111100; // 2537 : 252 - 0xfc
      12'h9EA: dout  = 8'b11111100; // 2538 : 252 - 0xfc
      12'h9EB: dout  = 8'b11111000; // 2539 : 248 - 0xf8
      12'h9EC: dout  = 8'b11111000; // 2540 : 248 - 0xf8
      12'h9ED: dout  = 8'b11111100; // 2541 : 252 - 0xfc
      12'h9EE: dout  = 8'b11111100; // 2542 : 252 - 0xfc
      12'h9EF: dout  = 8'b11111110; // 2543 : 254 - 0xfe
      12'h9F0: dout  = 8'b11111111; // 2544 : 255 - 0xff -- Background 0x9f
      12'h9F1: dout  = 8'b11111111; // 2545 : 255 - 0xff
      12'h9F2: dout  = 8'b10111101; // 2546 : 189 - 0xbd
      12'h9F3: dout  = 8'b11111111; // 2547 : 255 - 0xff
      12'h9F4: dout  = 8'b11111111; // 2548 : 255 - 0xff
      12'h9F5: dout  = 8'b11111111; // 2549 : 255 - 0xff
      12'h9F6: dout  = 8'b11111111; // 2550 : 255 - 0xff
      12'h9F7: dout  = 8'b10111101; // 2551 : 189 - 0xbd
      12'h9F8: dout  = 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout  = 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout  = 8'b01111110; // 2554 : 126 - 0x7e
      12'h9FB: dout  = 8'b01111110; // 2555 : 126 - 0x7e
      12'h9FC: dout  = 8'b01111110; // 2556 : 126 - 0x7e
      12'h9FD: dout  = 8'b01111110; // 2557 : 126 - 0x7e
      12'h9FE: dout  = 8'b01111110; // 2558 : 126 - 0x7e
      12'h9FF: dout  = 8'b01111110; // 2559 : 126 - 0x7e
      12'hA00: dout  = 8'b11101111; // 2560 : 239 - 0xef -- Background 0xa0
      12'hA01: dout  = 8'b11000111; // 2561 : 199 - 0xc7
      12'hA02: dout  = 8'b10000011; // 2562 : 131 - 0x83
      12'hA03: dout  = 8'b00000111; // 2563 :   7 - 0x7
      12'hA04: dout  = 8'b10001111; // 2564 : 143 - 0x8f
      12'hA05: dout  = 8'b11011101; // 2565 : 221 - 0xdd
      12'hA06: dout  = 8'b11111010; // 2566 : 250 - 0xfa
      12'hA07: dout  = 8'b11111101; // 2567 : 253 - 0xfd
      12'hA08: dout  = 8'b00010000; // 2568 :  16 - 0x10 -- plane 1
      12'hA09: dout  = 8'b00111000; // 2569 :  56 - 0x38
      12'hA0A: dout  = 8'b01111100; // 2570 : 124 - 0x7c
      12'hA0B: dout  = 8'b11111000; // 2571 : 248 - 0xf8
      12'hA0C: dout  = 8'b01110000; // 2572 : 112 - 0x70
      12'hA0D: dout  = 8'b00100010; // 2573 :  34 - 0x22
      12'hA0E: dout  = 8'b00000101; // 2574 :   5 - 0x5
      12'hA0F: dout  = 8'b00000010; // 2575 :   2 - 0x2
      12'hA10: dout  = 8'b11101111; // 2576 : 239 - 0xef -- Background 0xa1
      12'hA11: dout  = 8'b11000111; // 2577 : 199 - 0xc7
      12'hA12: dout  = 8'b10000011; // 2578 : 131 - 0x83
      12'hA13: dout  = 8'b00011111; // 2579 :  31 - 0x1f
      12'hA14: dout  = 8'b10010000; // 2580 : 144 - 0x90
      12'hA15: dout  = 8'b11010100; // 2581 : 212 - 0xd4
      12'hA16: dout  = 8'b11110011; // 2582 : 243 - 0xf3
      12'hA17: dout  = 8'b11110010; // 2583 : 242 - 0xf2
      12'hA18: dout  = 8'b00010000; // 2584 :  16 - 0x10 -- plane 1
      12'hA19: dout  = 8'b00111000; // 2585 :  56 - 0x38
      12'hA1A: dout  = 8'b01111100; // 2586 : 124 - 0x7c
      12'hA1B: dout  = 8'b11100000; // 2587 : 224 - 0xe0
      12'hA1C: dout  = 8'b01100000; // 2588 :  96 - 0x60
      12'hA1D: dout  = 8'b00100000; // 2589 :  32 - 0x20
      12'hA1E: dout  = 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout  = 8'b11101111; // 2592 : 239 - 0xef -- Background 0xa2
      12'hA21: dout  = 8'b11000111; // 2593 : 199 - 0xc7
      12'hA22: dout  = 8'b10000011; // 2594 : 131 - 0x83
      12'hA23: dout  = 8'b11111111; // 2595 : 255 - 0xff
      12'hA24: dout  = 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout  = 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout  = 8'b01010101; // 2598 :  85 - 0x55
      12'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout  = 8'b00010000; // 2600 :  16 - 0x10 -- plane 1
      12'hA29: dout  = 8'b00111000; // 2601 :  56 - 0x38
      12'hA2A: dout  = 8'b01111100; // 2602 : 124 - 0x7c
      12'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout  = 8'b11110000; // 2608 : 240 - 0xf0 -- Background 0xa3
      12'hA31: dout  = 8'b11010010; // 2609 : 210 - 0xd2
      12'hA32: dout  = 8'b10010000; // 2610 : 144 - 0x90
      12'hA33: dout  = 8'b00010010; // 2611 :  18 - 0x12
      12'hA34: dout  = 8'b10010000; // 2612 : 144 - 0x90
      12'hA35: dout  = 8'b11010010; // 2613 : 210 - 0xd2
      12'hA36: dout  = 8'b11110000; // 2614 : 240 - 0xf0
      12'hA37: dout  = 8'b11110010; // 2615 : 242 - 0xf2
      12'hA38: dout  = 8'b00000000; // 2616 :   0 - 0x0 -- plane 1
      12'hA39: dout  = 8'b00100000; // 2617 :  32 - 0x20
      12'hA3A: dout  = 8'b01100000; // 2618 :  96 - 0x60
      12'hA3B: dout  = 8'b11100000; // 2619 : 224 - 0xe0
      12'hA3C: dout  = 8'b01100000; // 2620 :  96 - 0x60
      12'hA3D: dout  = 8'b00100000; // 2621 :  32 - 0x20
      12'hA3E: dout  = 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b11110000; // 2624 : 240 - 0xf0 -- Background 0xa4
      12'hA41: dout  = 8'b11010011; // 2625 : 211 - 0xd3
      12'hA42: dout  = 8'b10010100; // 2626 : 148 - 0x94
      12'hA43: dout  = 8'b00011000; // 2627 :  24 - 0x18
      12'hA44: dout  = 8'b10011111; // 2628 : 159 - 0x9f
      12'hA45: dout  = 8'b11011101; // 2629 : 221 - 0xdd
      12'hA46: dout  = 8'b11111010; // 2630 : 250 - 0xfa
      12'hA47: dout  = 8'b11111101; // 2631 : 253 - 0xfd
      12'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout  = 8'b00100000; // 2633 :  32 - 0x20
      12'hA4A: dout  = 8'b01100011; // 2634 :  99 - 0x63
      12'hA4B: dout  = 8'b11100111; // 2635 : 231 - 0xe7
      12'hA4C: dout  = 8'b01100000; // 2636 :  96 - 0x60
      12'hA4D: dout  = 8'b00100010; // 2637 :  34 - 0x22
      12'hA4E: dout  = 8'b00000101; // 2638 :   5 - 0x5
      12'hA4F: dout  = 8'b00000010; // 2639 :   2 - 0x2
      12'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Background 0xa5
      12'hA51: dout  = 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout  = 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout  = 8'b11111111; // 2644 : 255 - 0xff
      12'hA55: dout  = 8'b11011101; // 2645 : 221 - 0xdd
      12'hA56: dout  = 8'b11111010; // 2646 : 250 - 0xfa
      12'hA57: dout  = 8'b11111101; // 2647 : 253 - 0xfd
      12'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout  = 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout  = 8'b11111111; // 2650 : 255 - 0xff
      12'hA5B: dout  = 8'b11111111; // 2651 : 255 - 0xff
      12'hA5C: dout  = 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout  = 8'b00100010; // 2653 :  34 - 0x22
      12'hA5E: dout  = 8'b00000101; // 2654 :   5 - 0x5
      12'hA5F: dout  = 8'b00000010; // 2655 :   2 - 0x2
      12'hA60: dout  = 8'b11101111; // 2656 : 239 - 0xef -- Background 0xa6
      12'hA61: dout  = 8'b11000111; // 2657 : 199 - 0xc7
      12'hA62: dout  = 8'b10000011; // 2658 : 131 - 0x83
      12'hA63: dout  = 8'b11111111; // 2659 : 255 - 0xff
      12'hA64: dout  = 8'b00011111; // 2660 :  31 - 0x1f
      12'hA65: dout  = 8'b00101101; // 2661 :  45 - 0x2d
      12'hA66: dout  = 8'b01001010; // 2662 :  74 - 0x4a
      12'hA67: dout  = 8'b01001101; // 2663 :  77 - 0x4d
      12'hA68: dout  = 8'b00010000; // 2664 :  16 - 0x10 -- plane 1
      12'hA69: dout  = 8'b00111000; // 2665 :  56 - 0x38
      12'hA6A: dout  = 8'b01111100; // 2666 : 124 - 0x7c
      12'hA6B: dout  = 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout  = 8'b00010010; // 2669 :  18 - 0x12
      12'hA6E: dout  = 8'b00110101; // 2670 :  53 - 0x35
      12'hA6F: dout  = 8'b00110010; // 2671 :  50 - 0x32
      12'hA70: dout  = 8'b01001111; // 2672 :  79 - 0x4f -- Background 0xa7
      12'hA71: dout  = 8'b01001111; // 2673 :  79 - 0x4f
      12'hA72: dout  = 8'b01001011; // 2674 :  75 - 0x4b
      12'hA73: dout  = 8'b01001111; // 2675 :  79 - 0x4f
      12'hA74: dout  = 8'b01001111; // 2676 :  79 - 0x4f
      12'hA75: dout  = 8'b01001101; // 2677 :  77 - 0x4d
      12'hA76: dout  = 8'b01001010; // 2678 :  74 - 0x4a
      12'hA77: dout  = 8'b01001101; // 2679 :  77 - 0x4d
      12'hA78: dout  = 8'b00110000; // 2680 :  48 - 0x30 -- plane 1
      12'hA79: dout  = 8'b00110000; // 2681 :  48 - 0x30
      12'hA7A: dout  = 8'b00110100; // 2682 :  52 - 0x34
      12'hA7B: dout  = 8'b00110000; // 2683 :  48 - 0x30
      12'hA7C: dout  = 8'b00110000; // 2684 :  48 - 0x30
      12'hA7D: dout  = 8'b00110010; // 2685 :  50 - 0x32
      12'hA7E: dout  = 8'b00110101; // 2686 :  53 - 0x35
      12'hA7F: dout  = 8'b00110010; // 2687 :  50 - 0x32
      12'hA80: dout  = 8'b01001111; // 2688 :  79 - 0x4f -- Background 0xa8
      12'hA81: dout  = 8'b11001111; // 2689 : 207 - 0xcf
      12'hA82: dout  = 8'b00001011; // 2690 :  11 - 0xb
      12'hA83: dout  = 8'b00001111; // 2691 :  15 - 0xf
      12'hA84: dout  = 8'b11111111; // 2692 : 255 - 0xff
      12'hA85: dout  = 8'b11011101; // 2693 : 221 - 0xdd
      12'hA86: dout  = 8'b11111010; // 2694 : 250 - 0xfa
      12'hA87: dout  = 8'b11111101; // 2695 : 253 - 0xfd
      12'hA88: dout  = 8'b00110000; // 2696 :  48 - 0x30 -- plane 1
      12'hA89: dout  = 8'b00110000; // 2697 :  48 - 0x30
      12'hA8A: dout  = 8'b11110100; // 2698 : 244 - 0xf4
      12'hA8B: dout  = 8'b11110000; // 2699 : 240 - 0xf0
      12'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout  = 8'b00100010; // 2701 :  34 - 0x22
      12'hA8E: dout  = 8'b00000101; // 2702 :   5 - 0x5
      12'hA8F: dout  = 8'b00000010; // 2703 :   2 - 0x2
      12'hA90: dout  = 8'b11111111; // 2704 : 255 - 0xff -- Background 0xa9
      12'hA91: dout  = 8'b11111111; // 2705 : 255 - 0xff
      12'hA92: dout  = 8'b11111111; // 2706 : 255 - 0xff
      12'hA93: dout  = 8'b11111111; // 2707 : 255 - 0xff
      12'hA94: dout  = 8'b11111111; // 2708 : 255 - 0xff
      12'hA95: dout  = 8'b11111111; // 2709 : 255 - 0xff
      12'hA96: dout  = 8'b11111111; // 2710 : 255 - 0xff
      12'hA97: dout  = 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0 -- plane 1
      12'hA99: dout  = 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout  = 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout  = 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout  = 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout  = 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout  = 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout  = 8'b11111111; // 2720 : 255 - 0xff -- Background 0xaa
      12'hAA1: dout  = 8'b11111111; // 2721 : 255 - 0xff
      12'hAA2: dout  = 8'b10101111; // 2722 : 175 - 0xaf
      12'hAA3: dout  = 8'b01010111; // 2723 :  87 - 0x57
      12'hAA4: dout  = 8'b10001111; // 2724 : 143 - 0x8f
      12'hAA5: dout  = 8'b11011101; // 2725 : 221 - 0xdd
      12'hAA6: dout  = 8'b11111010; // 2726 : 250 - 0xfa
      12'hAA7: dout  = 8'b11111101; // 2727 : 253 - 0xfd
      12'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout  = 8'b01010000; // 2730 :  80 - 0x50
      12'hAAB: dout  = 8'b10101000; // 2731 : 168 - 0xa8
      12'hAAC: dout  = 8'b01110000; // 2732 : 112 - 0x70
      12'hAAD: dout  = 8'b00100010; // 2733 :  34 - 0x22
      12'hAAE: dout  = 8'b00000101; // 2734 :   5 - 0x5
      12'hAAF: dout  = 8'b00000010; // 2735 :   2 - 0x2
      12'hAB0: dout  = 8'b11111111; // 2736 : 255 - 0xff -- Background 0xab
      12'hAB1: dout  = 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout  = 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout  = 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout  = 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout  = 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout  = 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout  = 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout  = 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout  = 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout  = 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout  = 8'b00000000; // 2752 :   0 - 0x0 -- Background 0xac
      12'hAC1: dout  = 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout  = 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout  = 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout  = 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout  = 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout  = 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout  = 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout  = 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout  = 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout  = 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout  = 8'b00000000; // 2768 :   0 - 0x0 -- Background 0xad
      12'hAD1: dout  = 8'b11111111; // 2769 : 255 - 0xff
      12'hAD2: dout  = 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout  = 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout  = 8'b11111111; // 2772 : 255 - 0xff
      12'hAD5: dout  = 8'b11111111; // 2773 : 255 - 0xff
      12'hAD6: dout  = 8'b11111111; // 2774 : 255 - 0xff
      12'hAD7: dout  = 8'b11111111; // 2775 : 255 - 0xff
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- plane 1
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b11111111; // 2778 : 255 - 0xff
      12'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout  = 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout  = 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout  = 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout  = 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout  = 8'b11111111; // 2784 : 255 - 0xff -- Background 0xae
      12'hAE1: dout  = 8'b11111111; // 2785 : 255 - 0xff
      12'hAE2: dout  = 8'b11111111; // 2786 : 255 - 0xff
      12'hAE3: dout  = 8'b11111111; // 2787 : 255 - 0xff
      12'hAE4: dout  = 8'b11111111; // 2788 : 255 - 0xff
      12'hAE5: dout  = 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout  = 8'b11111111; // 2790 : 255 - 0xff
      12'hAE7: dout  = 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout  = 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout  = 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout  = 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout  = 8'b11111111; // 2800 : 255 - 0xff -- Background 0xaf
      12'hAF1: dout  = 8'b11111111; // 2801 : 255 - 0xff
      12'hAF2: dout  = 8'b11111111; // 2802 : 255 - 0xff
      12'hAF3: dout  = 8'b11111111; // 2803 : 255 - 0xff
      12'hAF4: dout  = 8'b11111111; // 2804 : 255 - 0xff
      12'hAF5: dout  = 8'b11111111; // 2805 : 255 - 0xff
      12'hAF6: dout  = 8'b11111111; // 2806 : 255 - 0xff
      12'hAF7: dout  = 8'b11111111; // 2807 : 255 - 0xff
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout  = 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout  = 8'b00000000; // 2816 :   0 - 0x0 -- Background 0xb0
      12'hB01: dout  = 8'b00000000; // 2817 :   0 - 0x0
      12'hB02: dout  = 8'b00011111; // 2818 :  31 - 0x1f
      12'hB03: dout  = 8'b00010000; // 2819 :  16 - 0x10
      12'hB04: dout  = 8'b00010000; // 2820 :  16 - 0x10
      12'hB05: dout  = 8'b00010000; // 2821 :  16 - 0x10
      12'hB06: dout  = 8'b00010000; // 2822 :  16 - 0x10
      12'hB07: dout  = 8'b00010000; // 2823 :  16 - 0x10
      12'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout  = 8'b00011111; // 2826 :  31 - 0x1f
      12'hB0B: dout  = 8'b00011111; // 2827 :  31 - 0x1f
      12'hB0C: dout  = 8'b00011111; // 2828 :  31 - 0x1f
      12'hB0D: dout  = 8'b00011111; // 2829 :  31 - 0x1f
      12'hB0E: dout  = 8'b00011111; // 2830 :  31 - 0x1f
      12'hB0F: dout  = 8'b00011111; // 2831 :  31 - 0x1f
      12'hB10: dout  = 8'b00000000; // 2832 :   0 - 0x0 -- Background 0xb1
      12'hB11: dout  = 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout  = 8'b11111000; // 2834 : 248 - 0xf8
      12'hB13: dout  = 8'b00001000; // 2835 :   8 - 0x8
      12'hB14: dout  = 8'b00001000; // 2836 :   8 - 0x8
      12'hB15: dout  = 8'b00001000; // 2837 :   8 - 0x8
      12'hB16: dout  = 8'b00001000; // 2838 :   8 - 0x8
      12'hB17: dout  = 8'b00001000; // 2839 :   8 - 0x8
      12'hB18: dout  = 8'b00000000; // 2840 :   0 - 0x0 -- plane 1
      12'hB19: dout  = 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout  = 8'b11110000; // 2842 : 240 - 0xf0
      12'hB1B: dout  = 8'b11110000; // 2843 : 240 - 0xf0
      12'hB1C: dout  = 8'b11110000; // 2844 : 240 - 0xf0
      12'hB1D: dout  = 8'b11110000; // 2845 : 240 - 0xf0
      12'hB1E: dout  = 8'b11110000; // 2846 : 240 - 0xf0
      12'hB1F: dout  = 8'b11110000; // 2847 : 240 - 0xf0
      12'hB20: dout  = 8'b00010000; // 2848 :  16 - 0x10 -- Background 0xb2
      12'hB21: dout  = 8'b00010000; // 2849 :  16 - 0x10
      12'hB22: dout  = 8'b00010000; // 2850 :  16 - 0x10
      12'hB23: dout  = 8'b00010000; // 2851 :  16 - 0x10
      12'hB24: dout  = 8'b00010000; // 2852 :  16 - 0x10
      12'hB25: dout  = 8'b00011111; // 2853 :  31 - 0x1f
      12'hB26: dout  = 8'b00011111; // 2854 :  31 - 0x1f
      12'hB27: dout  = 8'b00001111; // 2855 :  15 - 0xf
      12'hB28: dout  = 8'b00011111; // 2856 :  31 - 0x1f -- plane 1
      12'hB29: dout  = 8'b00011111; // 2857 :  31 - 0x1f
      12'hB2A: dout  = 8'b00011111; // 2858 :  31 - 0x1f
      12'hB2B: dout  = 8'b00011111; // 2859 :  31 - 0x1f
      12'hB2C: dout  = 8'b00011111; // 2860 :  31 - 0x1f
      12'hB2D: dout  = 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout  = 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout  = 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout  = 8'b00001000; // 2864 :   8 - 0x8 -- Background 0xb3
      12'hB31: dout  = 8'b00001000; // 2865 :   8 - 0x8
      12'hB32: dout  = 8'b00001000; // 2866 :   8 - 0x8
      12'hB33: dout  = 8'b00001000; // 2867 :   8 - 0x8
      12'hB34: dout  = 8'b00001000; // 2868 :   8 - 0x8
      12'hB35: dout  = 8'b11111000; // 2869 : 248 - 0xf8
      12'hB36: dout  = 8'b11111000; // 2870 : 248 - 0xf8
      12'hB37: dout  = 8'b11110000; // 2871 : 240 - 0xf0
      12'hB38: dout  = 8'b11110000; // 2872 : 240 - 0xf0 -- plane 1
      12'hB39: dout  = 8'b11110000; // 2873 : 240 - 0xf0
      12'hB3A: dout  = 8'b11110000; // 2874 : 240 - 0xf0
      12'hB3B: dout  = 8'b11110000; // 2875 : 240 - 0xf0
      12'hB3C: dout  = 8'b11110000; // 2876 : 240 - 0xf0
      12'hB3D: dout  = 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout  = 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Background 0xb4
      12'hB41: dout  = 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout  = 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout  = 8'b00111111; // 2883 :  63 - 0x3f
      12'hB44: dout  = 8'b01100000; // 2884 :  96 - 0x60
      12'hB45: dout  = 8'b01100000; // 2885 :  96 - 0x60
      12'hB46: dout  = 8'b01100000; // 2886 :  96 - 0x60
      12'hB47: dout  = 8'b01100000; // 2887 :  96 - 0x60
      12'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0 -- plane 1
      12'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout  = 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout  = 8'b00111111; // 2891 :  63 - 0x3f
      12'hB4C: dout  = 8'b01111111; // 2892 : 127 - 0x7f
      12'hB4D: dout  = 8'b01111111; // 2893 : 127 - 0x7f
      12'hB4E: dout  = 8'b01111111; // 2894 : 127 - 0x7f
      12'hB4F: dout  = 8'b01111111; // 2895 : 127 - 0x7f
      12'hB50: dout  = 8'b00000000; // 2896 :   0 - 0x0 -- Background 0xb5
      12'hB51: dout  = 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout  = 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout  = 8'b11111100; // 2899 : 252 - 0xfc
      12'hB54: dout  = 8'b00000110; // 2900 :   6 - 0x6
      12'hB55: dout  = 8'b00000110; // 2901 :   6 - 0x6
      12'hB56: dout  = 8'b00000110; // 2902 :   6 - 0x6
      12'hB57: dout  = 8'b00000110; // 2903 :   6 - 0x6
      12'hB58: dout  = 8'b00000000; // 2904 :   0 - 0x0 -- plane 1
      12'hB59: dout  = 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout  = 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout  = 8'b11111000; // 2907 : 248 - 0xf8
      12'hB5C: dout  = 8'b11111000; // 2908 : 248 - 0xf8
      12'hB5D: dout  = 8'b11111000; // 2909 : 248 - 0xf8
      12'hB5E: dout  = 8'b11111000; // 2910 : 248 - 0xf8
      12'hB5F: dout  = 8'b11111000; // 2911 : 248 - 0xf8
      12'hB60: dout  = 8'b01100000; // 2912 :  96 - 0x60 -- Background 0xb6
      12'hB61: dout  = 8'b01100000; // 2913 :  96 - 0x60
      12'hB62: dout  = 8'b01100000; // 2914 :  96 - 0x60
      12'hB63: dout  = 8'b01100000; // 2915 :  96 - 0x60
      12'hB64: dout  = 8'b01111111; // 2916 : 127 - 0x7f
      12'hB65: dout  = 8'b01111111; // 2917 : 127 - 0x7f
      12'hB66: dout  = 8'b00111111; // 2918 :  63 - 0x3f
      12'hB67: dout  = 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout  = 8'b01111111; // 2920 : 127 - 0x7f -- plane 1
      12'hB69: dout  = 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout  = 8'b01111111; // 2922 : 127 - 0x7f
      12'hB6B: dout  = 8'b01111111; // 2923 : 127 - 0x7f
      12'hB6C: dout  = 8'b01000000; // 2924 :  64 - 0x40
      12'hB6D: dout  = 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout  = 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout  = 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout  = 8'b00000110; // 2928 :   6 - 0x6 -- Background 0xb7
      12'hB71: dout  = 8'b00000110; // 2929 :   6 - 0x6
      12'hB72: dout  = 8'b00000110; // 2930 :   6 - 0x6
      12'hB73: dout  = 8'b00000110; // 2931 :   6 - 0x6
      12'hB74: dout  = 8'b11111110; // 2932 : 254 - 0xfe
      12'hB75: dout  = 8'b11111110; // 2933 : 254 - 0xfe
      12'hB76: dout  = 8'b11111100; // 2934 : 252 - 0xfc
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b11111000; // 2936 : 248 - 0xf8 -- plane 1
      12'hB79: dout  = 8'b11111000; // 2937 : 248 - 0xf8
      12'hB7A: dout  = 8'b11111000; // 2938 : 248 - 0xf8
      12'hB7B: dout  = 8'b11111000; // 2939 : 248 - 0xf8
      12'hB7C: dout  = 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout  = 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout  = 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout  = 8'b01100000; // 2944 :  96 - 0x60 -- Background 0xb8
      12'hB81: dout  = 8'b11110000; // 2945 : 240 - 0xf0
      12'hB82: dout  = 8'b11000011; // 2946 : 195 - 0xc3
      12'hB83: dout  = 8'b10000111; // 2947 : 135 - 0x87
      12'hB84: dout  = 8'b00000110; // 2948 :   6 - 0x6
      12'hB85: dout  = 8'b00000100; // 2949 :   4 - 0x4
      12'hB86: dout  = 8'b00000100; // 2950 :   4 - 0x4
      12'hB87: dout  = 8'b00000111; // 2951 :   7 - 0x7
      12'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout  = 8'b00000011; // 2954 :   3 - 0x3
      12'hB8B: dout  = 8'b00000111; // 2955 :   7 - 0x7
      12'hB8C: dout  = 8'b00000111; // 2956 :   7 - 0x7
      12'hB8D: dout  = 8'b00000111; // 2957 :   7 - 0x7
      12'hB8E: dout  = 8'b00000011; // 2958 :   3 - 0x3
      12'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout  = 8'b00000110; // 2960 :   6 - 0x6 -- Background 0xb9
      12'hB91: dout  = 8'b00001111; // 2961 :  15 - 0xf
      12'hB92: dout  = 8'b10000111; // 2962 : 135 - 0x87
      12'hB93: dout  = 8'b11000001; // 2963 : 193 - 0xc1
      12'hB94: dout  = 8'b00100011; // 2964 :  35 - 0x23
      12'hB95: dout  = 8'b00101110; // 2965 :  46 - 0x2e
      12'hB96: dout  = 8'b01100000; // 2966 :  96 - 0x60
      12'hB97: dout  = 8'b11100001; // 2967 : 225 - 0xe1
      12'hB98: dout  = 8'b00000000; // 2968 :   0 - 0x0 -- plane 1
      12'hB99: dout  = 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout  = 8'b11000001; // 2970 : 193 - 0xc1
      12'hB9B: dout  = 8'b11100010; // 2971 : 226 - 0xe2
      12'hB9C: dout  = 8'b11001100; // 2972 : 204 - 0xcc
      12'hB9D: dout  = 8'b11000000; // 2973 : 192 - 0xc0
      12'hB9E: dout  = 8'b10000000; // 2974 : 128 - 0x80
      12'hB9F: dout  = 8'b00000001; // 2975 :   1 - 0x1
      12'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Background 0xba
      12'hBA1: dout  = 8'b11001000; // 2977 : 200 - 0xc8
      12'hBA2: dout  = 8'b11111000; // 2978 : 248 - 0xf8
      12'hBA3: dout  = 8'b10110000; // 2979 : 176 - 0xb0
      12'hBA4: dout  = 8'b00010000; // 2980 :  16 - 0x10
      12'hBA5: dout  = 8'b00110000; // 2981 :  48 - 0x30
      12'hBA6: dout  = 8'b11001000; // 2982 : 200 - 0xc8
      12'hBA7: dout  = 8'b11111000; // 2983 : 248 - 0xf8
      12'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout  = 8'b11110000; // 2985 : 240 - 0xf0
      12'hBAA: dout  = 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout  = 8'b00100000; // 2987 :  32 - 0x20
      12'hBAC: dout  = 8'b00100000; // 2988 :  32 - 0x20
      12'hBAD: dout  = 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout  = 8'b11110000; // 2990 : 240 - 0xf0
      12'hBAF: dout  = 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout  = 8'b00000111; // 2992 :   7 - 0x7 -- Background 0xbb
      12'hBB1: dout  = 8'b00000011; // 2993 :   3 - 0x3
      12'hBB2: dout  = 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout  = 8'b01100000; // 2995 :  96 - 0x60
      12'hBB4: dout  = 8'b11110000; // 2996 : 240 - 0xf0
      12'hBB5: dout  = 8'b11010000; // 2997 : 208 - 0xd0
      12'hBB6: dout  = 8'b10010000; // 2998 : 144 - 0x90
      12'hBB7: dout  = 8'b01100000; // 2999 :  96 - 0x60
      12'hBB8: dout  = 8'b00000000; // 3000 :   0 - 0x0 -- plane 1
      12'hBB9: dout  = 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout  = 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout  = 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout  = 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout  = 8'b01100000; // 3005 :  96 - 0x60
      12'hBBE: dout  = 8'b01100000; // 3006 :  96 - 0x60
      12'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout  = 8'b11100001; // 3008 : 225 - 0xe1 -- Background 0xbc
      12'hBC1: dout  = 8'b11000011; // 3009 : 195 - 0xc3
      12'hBC2: dout  = 8'b00001110; // 3010 :  14 - 0xe
      12'hBC3: dout  = 8'b00000110; // 3011 :   6 - 0x6
      12'hBC4: dout  = 8'b00001111; // 3012 :  15 - 0xf
      12'hBC5: dout  = 8'b00001101; // 3013 :  13 - 0xd
      12'hBC6: dout  = 8'b00001001; // 3014 :   9 - 0x9
      12'hBC7: dout  = 8'b00000110; // 3015 :   6 - 0x6
      12'hBC8: dout  = 8'b00000010; // 3016 :   2 - 0x2 -- plane 1
      12'hBC9: dout  = 8'b00001100; // 3017 :  12 - 0xc
      12'hBCA: dout  = 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout  = 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout  = 8'b00000110; // 3021 :   6 - 0x6
      12'hBCE: dout  = 8'b00000110; // 3022 :   6 - 0x6
      12'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout  = 8'b11100000; // 3024 : 224 - 0xe0 -- Background 0xbd
      12'hBD1: dout  = 8'b01100000; // 3025 :  96 - 0x60
      12'hBD2: dout  = 8'b11100011; // 3026 : 227 - 0xe3
      12'hBD3: dout  = 8'b11100111; // 3027 : 231 - 0xe7
      12'hBD4: dout  = 8'b00000110; // 3028 :   6 - 0x6
      12'hBD5: dout  = 8'b00000100; // 3029 :   4 - 0x4
      12'hBD6: dout  = 8'b00000100; // 3030 :   4 - 0x4
      12'hBD7: dout  = 8'b00000111; // 3031 :   7 - 0x7
      12'hBD8: dout  = 8'b00000000; // 3032 :   0 - 0x0 -- plane 1
      12'hBD9: dout  = 8'b10000000; // 3033 : 128 - 0x80
      12'hBDA: dout  = 8'b00000011; // 3034 :   3 - 0x3
      12'hBDB: dout  = 8'b00000111; // 3035 :   7 - 0x7
      12'hBDC: dout  = 8'b00000111; // 3036 :   7 - 0x7
      12'hBDD: dout  = 8'b00000111; // 3037 :   7 - 0x7
      12'hBDE: dout  = 8'b00000011; // 3038 :   3 - 0x3
      12'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout  = 8'b00000111; // 3040 :   7 - 0x7 -- Background 0xbe
      12'hBE1: dout  = 8'b00000011; // 3041 :   3 - 0x3
      12'hBE2: dout  = 8'b10000111; // 3042 : 135 - 0x87
      12'hBE3: dout  = 8'b11000111; // 3043 : 199 - 0xc7
      12'hBE4: dout  = 8'b00100000; // 3044 :  32 - 0x20
      12'hBE5: dout  = 8'b00100000; // 3045 :  32 - 0x20
      12'hBE6: dout  = 8'b01100000; // 3046 :  96 - 0x60
      12'hBE7: dout  = 8'b11100000; // 3047 : 224 - 0xe0
      12'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout  = 8'b00000100; // 3049 :   4 - 0x4
      12'hBEA: dout  = 8'b11000000; // 3050 : 192 - 0xc0
      12'hBEB: dout  = 8'b11100000; // 3051 : 224 - 0xe0
      12'hBEC: dout  = 8'b11000000; // 3052 : 192 - 0xc0
      12'hBED: dout  = 8'b11000000; // 3053 : 192 - 0xc0
      12'hBEE: dout  = 8'b10000000; // 3054 : 128 - 0x80
      12'hBEF: dout  = 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout  = 8'b00000111; // 3056 :   7 - 0x7 -- Background 0xbf
      12'hBF1: dout  = 8'b00000011; // 3057 :   3 - 0x3
      12'hBF2: dout  = 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout  = 8'b00001100; // 3059 :  12 - 0xc
      12'hBF4: dout  = 8'b11101100; // 3060 : 236 - 0xec
      12'hBF5: dout  = 8'b01100100; // 3061 : 100 - 0x64
      12'hBF6: dout  = 8'b11101100; // 3062 : 236 - 0xec
      12'hBF7: dout  = 8'b11101101; // 3063 : 237 - 0xed
      12'hBF8: dout  = 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout  = 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout  = 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout  = 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout  = 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout  = 8'b10001000; // 3069 : 136 - 0x88
      12'hBFE: dout  = 8'b00001000; // 3070 :   8 - 0x8
      12'hBFF: dout  = 8'b00001011; // 3071 :  11 - 0xb
      12'hC00: dout  = 8'b11100000; // 3072 : 224 - 0xe0 -- Background 0xc0
      12'hC01: dout  = 8'b11000000; // 3073 : 192 - 0xc0
      12'hC02: dout  = 8'b00000000; // 3074 :   0 - 0x0
      12'hC03: dout  = 8'b00110000; // 3075 :  48 - 0x30
      12'hC04: dout  = 8'b00110111; // 3076 :  55 - 0x37
      12'hC05: dout  = 8'b00010011; // 3077 :  19 - 0x13
      12'hC06: dout  = 8'b00110111; // 3078 :  55 - 0x37
      12'hC07: dout  = 8'b01110111; // 3079 : 119 - 0x77
      12'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout  = 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout  = 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout  = 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout  = 8'b00100100; // 3085 :  36 - 0x24
      12'hC0E: dout  = 8'b00100000; // 3086 :  32 - 0x20
      12'hC0F: dout  = 8'b10100000; // 3087 : 160 - 0xa0
      12'hC10: dout  = 8'b00001111; // 3088 :  15 - 0xf -- Background 0xc1
      12'hC11: dout  = 8'b00001100; // 3089 :  12 - 0xc
      12'hC12: dout  = 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout  = 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout  = 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout  = 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout  = 8'b00000000; // 3094 :   0 - 0x0
      12'hC17: dout  = 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout  = 8'b00000000; // 3096 :   0 - 0x0 -- plane 1
      12'hC19: dout  = 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout  = 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout  = 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout  = 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout  = 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout  = 8'b11110000; // 3104 : 240 - 0xf0 -- Background 0xc2
      12'hC21: dout  = 8'b00110000; // 3105 :  48 - 0x30
      12'hC22: dout  = 8'b00000000; // 3106 :   0 - 0x0
      12'hC23: dout  = 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout  = 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout  = 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout  = 8'b00000000; // 3110 :   0 - 0x0
      12'hC27: dout  = 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout  = 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout  = 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout  = 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout  = 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout  = 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout  = 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Background 0xc3
      12'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout  = 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout  = 8'b00000100; // 3123 :   4 - 0x4
      12'hC34: dout  = 8'b00001101; // 3124 :  13 - 0xd
      12'hC35: dout  = 8'b00001111; // 3125 :  15 - 0xf
      12'hC36: dout  = 8'b00001100; // 3126 :  12 - 0xc
      12'hC37: dout  = 8'b00001100; // 3127 :  12 - 0xc
      12'hC38: dout  = 8'b00000000; // 3128 :   0 - 0x0 -- plane 1
      12'hC39: dout  = 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout  = 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout  = 8'b00001000; // 3131 :   8 - 0x8
      12'hC3C: dout  = 8'b00001011; // 3132 :  11 - 0xb
      12'hC3D: dout  = 8'b00001000; // 3133 :   8 - 0x8
      12'hC3E: dout  = 8'b00001000; // 3134 :   8 - 0x8
      12'hC3F: dout  = 8'b00001000; // 3135 :   8 - 0x8
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Background 0xc4
      12'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout  = 8'b00010000; // 3139 :  16 - 0x10
      12'hC44: dout  = 8'b01110000; // 3140 : 112 - 0x70
      12'hC45: dout  = 8'b11110000; // 3141 : 240 - 0xf0
      12'hC46: dout  = 8'b00110000; // 3142 :  48 - 0x30
      12'hC47: dout  = 8'b00110000; // 3143 :  48 - 0x30
      12'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout  = 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout  = 8'b00100000; // 3147 :  32 - 0x20
      12'hC4C: dout  = 8'b10100000; // 3148 : 160 - 0xa0
      12'hC4D: dout  = 8'b00100000; // 3149 :  32 - 0x20
      12'hC4E: dout  = 8'b00100000; // 3150 :  32 - 0x20
      12'hC4F: dout  = 8'b00100000; // 3151 :  32 - 0x20
      12'hC50: dout  = 8'b11100100; // 3152 : 228 - 0xe4 -- Background 0xc5
      12'hC51: dout  = 8'b00100100; // 3153 :  36 - 0x24
      12'hC52: dout  = 8'b11100100; // 3154 : 228 - 0xe4
      12'hC53: dout  = 8'b11101111; // 3155 : 239 - 0xef
      12'hC54: dout  = 8'b00000111; // 3156 :   7 - 0x7
      12'hC55: dout  = 8'b00000110; // 3157 :   6 - 0x6
      12'hC56: dout  = 8'b00000100; // 3158 :   4 - 0x4
      12'hC57: dout  = 8'b00000100; // 3159 :   4 - 0x4
      12'hC58: dout  = 8'b00001000; // 3160 :   8 - 0x8 -- plane 1
      12'hC59: dout  = 8'b11001000; // 3161 : 200 - 0xc8
      12'hC5A: dout  = 8'b00001000; // 3162 :   8 - 0x8
      12'hC5B: dout  = 8'b00000011; // 3163 :   3 - 0x3
      12'hC5C: dout  = 8'b00000111; // 3164 :   7 - 0x7
      12'hC5D: dout  = 8'b00000111; // 3165 :   7 - 0x7
      12'hC5E: dout  = 8'b00000111; // 3166 :   7 - 0x7
      12'hC5F: dout  = 8'b00000011; // 3167 :   3 - 0x3
      12'hC60: dout  = 8'b00010111; // 3168 :  23 - 0x17 -- Background 0xc6
      12'hC61: dout  = 8'b00010001; // 3169 :  17 - 0x11
      12'hC62: dout  = 8'b00010111; // 3170 :  23 - 0x17
      12'hC63: dout  = 8'b10110111; // 3171 : 183 - 0xb7
      12'hC64: dout  = 8'b11000000; // 3172 : 192 - 0xc0
      12'hC65: dout  = 8'b00100000; // 3173 :  32 - 0x20
      12'hC66: dout  = 8'b00100000; // 3174 :  32 - 0x20
      12'hC67: dout  = 8'b01100000; // 3175 :  96 - 0x60
      12'hC68: dout  = 8'b00100000; // 3176 :  32 - 0x20 -- plane 1
      12'hC69: dout  = 8'b00100110; // 3177 :  38 - 0x26
      12'hC6A: dout  = 8'b00100000; // 3178 :  32 - 0x20
      12'hC6B: dout  = 8'b11000000; // 3179 : 192 - 0xc0
      12'hC6C: dout  = 8'b11100000; // 3180 : 224 - 0xe0
      12'hC6D: dout  = 8'b11000000; // 3181 : 192 - 0xc0
      12'hC6E: dout  = 8'b11000000; // 3182 : 192 - 0xc0
      12'hC6F: dout  = 8'b10000000; // 3183 : 128 - 0x80
      12'hC70: dout  = 8'b00000111; // 3184 :   7 - 0x7 -- Background 0xc7
      12'hC71: dout  = 8'b00000111; // 3185 :   7 - 0x7
      12'hC72: dout  = 8'b00000011; // 3186 :   3 - 0x3
      12'hC73: dout  = 8'b00000000; // 3187 :   0 - 0x0
      12'hC74: dout  = 8'b11100000; // 3188 : 224 - 0xe0
      12'hC75: dout  = 8'b00100000; // 3189 :  32 - 0x20
      12'hC76: dout  = 8'b11100000; // 3190 : 224 - 0xe0
      12'hC77: dout  = 8'b11100000; // 3191 : 224 - 0xe0
      12'hC78: dout  = 8'b00000000; // 3192 :   0 - 0x0 -- plane 1
      12'hC79: dout  = 8'b00000000; // 3193 :   0 - 0x0
      12'hC7A: dout  = 8'b00000000; // 3194 :   0 - 0x0
      12'hC7B: dout  = 8'b00000000; // 3195 :   0 - 0x0
      12'hC7C: dout  = 8'b00000000; // 3196 :   0 - 0x0
      12'hC7D: dout  = 8'b11000000; // 3197 : 192 - 0xc0
      12'hC7E: dout  = 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout  = 8'b11100000; // 3200 : 224 - 0xe0 -- Background 0xc8
      12'hC81: dout  = 8'b11100000; // 3201 : 224 - 0xe0
      12'hC82: dout  = 8'b11000000; // 3202 : 192 - 0xc0
      12'hC83: dout  = 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout  = 8'b00000111; // 3204 :   7 - 0x7
      12'hC85: dout  = 8'b00000001; // 3205 :   1 - 0x1
      12'hC86: dout  = 8'b00000111; // 3206 :   7 - 0x7
      12'hC87: dout  = 8'b00000111; // 3207 :   7 - 0x7
      12'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout  = 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout  = 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout  = 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout  = 8'b00000110; // 3213 :   6 - 0x6
      12'hC8E: dout  = 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout  = 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout  = 8'b00000001; // 3216 :   1 - 0x1 -- Background 0xc9
      12'hC91: dout  = 8'b00010011; // 3217 :  19 - 0x13
      12'hC92: dout  = 8'b00011111; // 3218 :  31 - 0x1f
      12'hC93: dout  = 8'b00001101; // 3219 :  13 - 0xd
      12'hC94: dout  = 8'b00000100; // 3220 :   4 - 0x4
      12'hC95: dout  = 8'b00001100; // 3221 :  12 - 0xc
      12'hC96: dout  = 8'b00010011; // 3222 :  19 - 0x13
      12'hC97: dout  = 8'b00011111; // 3223 :  31 - 0x1f
      12'hC98: dout  = 8'b00000000; // 3224 :   0 - 0x0 -- plane 1
      12'hC99: dout  = 8'b00001111; // 3225 :  15 - 0xf
      12'hC9A: dout  = 8'b00000000; // 3226 :   0 - 0x0
      12'hC9B: dout  = 8'b00001000; // 3227 :   8 - 0x8
      12'hC9C: dout  = 8'b00001000; // 3228 :   8 - 0x8
      12'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout  = 8'b00001111; // 3230 :  15 - 0xf
      12'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout  = 8'b01100000; // 3232 :  96 - 0x60 -- Background 0xca
      12'hCA1: dout  = 8'b01110000; // 3233 : 112 - 0x70
      12'hCA2: dout  = 8'b10100011; // 3234 : 163 - 0xa3
      12'hCA3: dout  = 8'b10000111; // 3235 : 135 - 0x87
      12'hCA4: dout  = 8'b11000110; // 3236 : 198 - 0xc6
      12'hCA5: dout  = 8'b01110100; // 3237 : 116 - 0x74
      12'hCA6: dout  = 8'b00000100; // 3238 :   4 - 0x4
      12'hCA7: dout  = 8'b10000111; // 3239 : 135 - 0x87
      12'hCA8: dout  = 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout  = 8'b00000000; // 3241 :   0 - 0x0
      12'hCAA: dout  = 8'b10000011; // 3242 : 131 - 0x83
      12'hCAB: dout  = 8'b01000111; // 3243 :  71 - 0x47
      12'hCAC: dout  = 8'b00110111; // 3244 :  55 - 0x37
      12'hCAD: dout  = 8'b00000111; // 3245 :   7 - 0x7
      12'hCAE: dout  = 8'b00000011; // 3246 :   3 - 0x3
      12'hCAF: dout  = 8'b10000000; // 3247 : 128 - 0x80
      12'hCB0: dout  = 8'b00000110; // 3248 :   6 - 0x6 -- Background 0xcb
      12'hCB1: dout  = 8'b00001111; // 3249 :  15 - 0xf
      12'hCB2: dout  = 8'b10000011; // 3250 : 131 - 0x83
      12'hCB3: dout  = 8'b11000001; // 3251 : 193 - 0xc1
      12'hCB4: dout  = 8'b00100000; // 3252 :  32 - 0x20
      12'hCB5: dout  = 8'b00100000; // 3253 :  32 - 0x20
      12'hCB6: dout  = 8'b01100000; // 3254 :  96 - 0x60
      12'hCB7: dout  = 8'b11100000; // 3255 : 224 - 0xe0
      12'hCB8: dout  = 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout  = 8'b00000000; // 3257 :   0 - 0x0
      12'hCBA: dout  = 8'b11000000; // 3258 : 192 - 0xc0
      12'hCBB: dout  = 8'b11100000; // 3259 : 224 - 0xe0
      12'hCBC: dout  = 8'b11000000; // 3260 : 192 - 0xc0
      12'hCBD: dout  = 8'b11000000; // 3261 : 192 - 0xc0
      12'hCBE: dout  = 8'b10000000; // 3262 : 128 - 0x80
      12'hCBF: dout  = 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout  = 8'b10000111; // 3264 : 135 - 0x87 -- Background 0xcc
      12'hCC1: dout  = 8'b01000011; // 3265 :  67 - 0x43
      12'hCC2: dout  = 8'b00110000; // 3266 :  48 - 0x30
      12'hCC3: dout  = 8'b01100000; // 3267 :  96 - 0x60
      12'hCC4: dout  = 8'b11110000; // 3268 : 240 - 0xf0
      12'hCC5: dout  = 8'b11010000; // 3269 : 208 - 0xd0
      12'hCC6: dout  = 8'b10010000; // 3270 : 144 - 0x90
      12'hCC7: dout  = 8'b01100000; // 3271 :  96 - 0x60
      12'hCC8: dout  = 8'b01000000; // 3272 :  64 - 0x40 -- plane 1
      12'hCC9: dout  = 8'b00110000; // 3273 :  48 - 0x30
      12'hCCA: dout  = 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout  = 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout  = 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout  = 8'b01100000; // 3277 :  96 - 0x60
      12'hCCE: dout  = 8'b01100000; // 3278 :  96 - 0x60
      12'hCCF: dout  = 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout  = 8'b11100000; // 3280 : 224 - 0xe0 -- Background 0xcd
      12'hCD1: dout  = 8'b11000000; // 3281 : 192 - 0xc0
      12'hCD2: dout  = 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout  = 8'b00000110; // 3283 :   6 - 0x6
      12'hCD4: dout  = 8'b00001111; // 3284 :  15 - 0xf
      12'hCD5: dout  = 8'b00001101; // 3285 :  13 - 0xd
      12'hCD6: dout  = 8'b00001001; // 3286 :   9 - 0x9
      12'hCD7: dout  = 8'b00000110; // 3287 :   6 - 0x6
      12'hCD8: dout  = 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout  = 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout  = 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout  = 8'b00000000; // 3291 :   0 - 0x0
      12'hCDC: dout  = 8'b00000000; // 3292 :   0 - 0x0
      12'hCDD: dout  = 8'b00000110; // 3293 :   6 - 0x6
      12'hCDE: dout  = 8'b00000110; // 3294 :   6 - 0x6
      12'hCDF: dout  = 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout  = 8'b11111100; // 3296 : 252 - 0xfc -- Background 0xce
      12'hCE1: dout  = 8'b11000000; // 3297 : 192 - 0xc0
      12'hCE2: dout  = 8'b11010001; // 3298 : 209 - 0xd1
      12'hCE3: dout  = 8'b11000010; // 3299 : 194 - 0xc2
      12'hCE4: dout  = 8'b10011110; // 3300 : 158 - 0x9e
      12'hCE5: dout  = 8'b10111111; // 3301 : 191 - 0xbf
      12'hCE6: dout  = 8'b10110000; // 3302 : 176 - 0xb0
      12'hCE7: dout  = 8'b10110011; // 3303 : 179 - 0xb3
      12'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout  = 8'b00000001; // 3305 :   1 - 0x1
      12'hCEA: dout  = 8'b00011011; // 3306 :  27 - 0x1b
      12'hCEB: dout  = 8'b00010011; // 3307 :  19 - 0x13
      12'hCEC: dout  = 8'b00011111; // 3308 :  31 - 0x1f
      12'hCED: dout  = 8'b00111111; // 3309 :  63 - 0x3f
      12'hCEE: dout  = 8'b00111111; // 3310 :  63 - 0x3f
      12'hCEF: dout  = 8'b00111111; // 3311 :  63 - 0x3f
      12'hCF0: dout  = 8'b00000111; // 3312 :   7 - 0x7 -- Background 0xcf
      12'hCF1: dout  = 8'b11110011; // 3313 : 243 - 0xf3
      12'hCF2: dout  = 8'b00001011; // 3314 :  11 - 0xb
      12'hCF3: dout  = 8'b01111011; // 3315 : 123 - 0x7b
      12'hCF4: dout  = 8'b01111011; // 3316 : 123 - 0x7b
      12'hCF5: dout  = 8'b11111001; // 3317 : 249 - 0xf9
      12'hCF6: dout  = 8'b00001101; // 3318 :  13 - 0xd
      12'hCF7: dout  = 8'b11101101; // 3319 : 237 - 0xed
      12'hCF8: dout  = 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout  = 8'b11111000; // 3321 : 248 - 0xf8
      12'hCFA: dout  = 8'b00001000; // 3322 :   8 - 0x8
      12'hCFB: dout  = 8'b00001000; // 3323 :   8 - 0x8
      12'hCFC: dout  = 8'b00001000; // 3324 :   8 - 0x8
      12'hCFD: dout  = 8'b11111000; // 3325 : 248 - 0xf8
      12'hCFE: dout  = 8'b11110000; // 3326 : 240 - 0xf0
      12'hCFF: dout  = 8'b11010000; // 3327 : 208 - 0xd0
      12'hD00: dout  = 8'b11111111; // 3328 : 255 - 0xff -- Background 0xd0
      12'hD01: dout  = 8'b11111111; // 3329 : 255 - 0xff
      12'hD02: dout  = 8'b11111111; // 3330 : 255 - 0xff
      12'hD03: dout  = 8'b11111111; // 3331 : 255 - 0xff
      12'hD04: dout  = 8'b11101110; // 3332 : 238 - 0xee
      12'hD05: dout  = 8'b11101110; // 3333 : 238 - 0xee
      12'hD06: dout  = 8'b11101110; // 3334 : 238 - 0xee
      12'hD07: dout  = 8'b11101110; // 3335 : 238 - 0xee
      12'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout  = 8'b01111100; // 3338 : 124 - 0x7c
      12'hD0B: dout  = 8'b11111110; // 3339 : 254 - 0xfe
      12'hD0C: dout  = 8'b11101110; // 3340 : 238 - 0xee
      12'hD0D: dout  = 8'b11101110; // 3341 : 238 - 0xee
      12'hD0E: dout  = 8'b11101110; // 3342 : 238 - 0xee
      12'hD0F: dout  = 8'b11101110; // 3343 : 238 - 0xee
      12'hD10: dout  = 8'b11111111; // 3344 : 255 - 0xff -- Background 0xd1
      12'hD11: dout  = 8'b11111111; // 3345 : 255 - 0xff
      12'hD12: dout  = 8'b11111111; // 3346 : 255 - 0xff
      12'hD13: dout  = 8'b11111011; // 3347 : 251 - 0xfb
      12'hD14: dout  = 8'b11111011; // 3348 : 251 - 0xfb
      12'hD15: dout  = 8'b11111011; // 3349 : 251 - 0xfb
      12'hD16: dout  = 8'b11111011; // 3350 : 251 - 0xfb
      12'hD17: dout  = 8'b11111011; // 3351 : 251 - 0xfb
      12'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout  = 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout  = 8'b00111000; // 3354 :  56 - 0x38
      12'hD1B: dout  = 8'b01111000; // 3355 : 120 - 0x78
      12'hD1C: dout  = 8'b01111000; // 3356 : 120 - 0x78
      12'hD1D: dout  = 8'b00111000; // 3357 :  56 - 0x38
      12'hD1E: dout  = 8'b00111000; // 3358 :  56 - 0x38
      12'hD1F: dout  = 8'b00111000; // 3359 :  56 - 0x38
      12'hD20: dout  = 8'b11111111; // 3360 : 255 - 0xff -- Background 0xd2
      12'hD21: dout  = 8'b11111111; // 3361 : 255 - 0xff
      12'hD22: dout  = 8'b11111111; // 3362 : 255 - 0xff
      12'hD23: dout  = 8'b11111111; // 3363 : 255 - 0xff
      12'hD24: dout  = 8'b11101110; // 3364 : 238 - 0xee
      12'hD25: dout  = 8'b10001110; // 3365 : 142 - 0x8e
      12'hD26: dout  = 8'b11111110; // 3366 : 254 - 0xfe
      12'hD27: dout  = 8'b11111110; // 3367 : 254 - 0xfe
      12'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout  = 8'b01111100; // 3370 : 124 - 0x7c
      12'hD2B: dout  = 8'b11111110; // 3371 : 254 - 0xfe
      12'hD2C: dout  = 8'b11101110; // 3372 : 238 - 0xee
      12'hD2D: dout  = 8'b00001110; // 3373 :  14 - 0xe
      12'hD2E: dout  = 8'b00001110; // 3374 :  14 - 0xe
      12'hD2F: dout  = 8'b01111110; // 3375 : 126 - 0x7e
      12'hD30: dout  = 8'b11111111; // 3376 : 255 - 0xff -- Background 0xd3
      12'hD31: dout  = 8'b11111111; // 3377 : 255 - 0xff
      12'hD32: dout  = 8'b11111111; // 3378 : 255 - 0xff
      12'hD33: dout  = 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout  = 8'b11101110; // 3380 : 238 - 0xee
      12'hD35: dout  = 8'b10001110; // 3381 : 142 - 0x8e
      12'hD36: dout  = 8'b11111100; // 3382 : 252 - 0xfc
      12'hD37: dout  = 8'b11111101; // 3383 : 253 - 0xfd
      12'hD38: dout  = 8'b00000000; // 3384 :   0 - 0x0 -- plane 1
      12'hD39: dout  = 8'b00000000; // 3385 :   0 - 0x0
      12'hD3A: dout  = 8'b01111100; // 3386 : 124 - 0x7c
      12'hD3B: dout  = 8'b11111110; // 3387 : 254 - 0xfe
      12'hD3C: dout  = 8'b11101110; // 3388 : 238 - 0xee
      12'hD3D: dout  = 8'b00001110; // 3389 :  14 - 0xe
      12'hD3E: dout  = 8'b00111100; // 3390 :  60 - 0x3c
      12'hD3F: dout  = 8'b00111100; // 3391 :  60 - 0x3c
      12'hD40: dout  = 8'b11111111; // 3392 : 255 - 0xff -- Background 0xd4
      12'hD41: dout  = 8'b11111111; // 3393 : 255 - 0xff
      12'hD42: dout  = 8'b11111111; // 3394 : 255 - 0xff
      12'hD43: dout  = 8'b11111110; // 3395 : 254 - 0xfe
      12'hD44: dout  = 8'b11101110; // 3396 : 238 - 0xee
      12'hD45: dout  = 8'b11101110; // 3397 : 238 - 0xee
      12'hD46: dout  = 8'b11101110; // 3398 : 238 - 0xee
      12'hD47: dout  = 8'b11101110; // 3399 : 238 - 0xee
      12'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout  = 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout  = 8'b00111110; // 3402 :  62 - 0x3e
      12'hD4B: dout  = 8'b01111110; // 3403 : 126 - 0x7e
      12'hD4C: dout  = 8'b11101110; // 3404 : 238 - 0xee
      12'hD4D: dout  = 8'b11101110; // 3405 : 238 - 0xee
      12'hD4E: dout  = 8'b11101110; // 3406 : 238 - 0xee
      12'hD4F: dout  = 8'b11101110; // 3407 : 238 - 0xee
      12'hD50: dout  = 8'b11111111; // 3408 : 255 - 0xff -- Background 0xd5
      12'hD51: dout  = 8'b11111111; // 3409 : 255 - 0xff
      12'hD52: dout  = 8'b11111111; // 3410 : 255 - 0xff
      12'hD53: dout  = 8'b11111101; // 3411 : 253 - 0xfd
      12'hD54: dout  = 8'b11100001; // 3412 : 225 - 0xe1
      12'hD55: dout  = 8'b11101111; // 3413 : 239 - 0xef
      12'hD56: dout  = 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout  = 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout  = 8'b11111100; // 3418 : 252 - 0xfc
      12'hD5B: dout  = 8'b11111100; // 3419 : 252 - 0xfc
      12'hD5C: dout  = 8'b11100000; // 3420 : 224 - 0xe0
      12'hD5D: dout  = 8'b11100000; // 3421 : 224 - 0xe0
      12'hD5E: dout  = 8'b11111100; // 3422 : 252 - 0xfc
      12'hD5F: dout  = 8'b11111110; // 3423 : 254 - 0xfe
      12'hD60: dout  = 8'b11111111; // 3424 : 255 - 0xff -- Background 0xd6
      12'hD61: dout  = 8'b11111111; // 3425 : 255 - 0xff
      12'hD62: dout  = 8'b11111111; // 3426 : 255 - 0xff
      12'hD63: dout  = 8'b11111101; // 3427 : 253 - 0xfd
      12'hD64: dout  = 8'b11100001; // 3428 : 225 - 0xe1
      12'hD65: dout  = 8'b11101111; // 3429 : 239 - 0xef
      12'hD66: dout  = 8'b11111111; // 3430 : 255 - 0xff
      12'hD67: dout  = 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout  = 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout  = 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout  = 8'b01111100; // 3434 : 124 - 0x7c
      12'hD6B: dout  = 8'b11111100; // 3435 : 252 - 0xfc
      12'hD6C: dout  = 8'b11100000; // 3436 : 224 - 0xe0
      12'hD6D: dout  = 8'b11100000; // 3437 : 224 - 0xe0
      12'hD6E: dout  = 8'b11111100; // 3438 : 252 - 0xfc
      12'hD6F: dout  = 8'b11111110; // 3439 : 254 - 0xfe
      12'hD70: dout  = 8'b11111111; // 3440 : 255 - 0xff -- Background 0xd7
      12'hD71: dout  = 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout  = 8'b11111111; // 3442 : 255 - 0xff
      12'hD73: dout  = 8'b11111110; // 3443 : 254 - 0xfe
      12'hD74: dout  = 8'b11101110; // 3444 : 238 - 0xee
      12'hD75: dout  = 8'b10001110; // 3445 : 142 - 0x8e
      12'hD76: dout  = 8'b11111110; // 3446 : 254 - 0xfe
      12'hD77: dout  = 8'b11111100; // 3447 : 252 - 0xfc
      12'hD78: dout  = 8'b00000000; // 3448 :   0 - 0x0 -- plane 1
      12'hD79: dout  = 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout  = 8'b11111110; // 3450 : 254 - 0xfe
      12'hD7B: dout  = 8'b11111110; // 3451 : 254 - 0xfe
      12'hD7C: dout  = 8'b11101110; // 3452 : 238 - 0xee
      12'hD7D: dout  = 8'b00001110; // 3453 :  14 - 0xe
      12'hD7E: dout  = 8'b00001110; // 3454 :  14 - 0xe
      12'hD7F: dout  = 8'b00011100; // 3455 :  28 - 0x1c
      12'hD80: dout  = 8'b11111111; // 3456 : 255 - 0xff -- Background 0xd8
      12'hD81: dout  = 8'b11111111; // 3457 : 255 - 0xff
      12'hD82: dout  = 8'b11111111; // 3458 : 255 - 0xff
      12'hD83: dout  = 8'b11111111; // 3459 : 255 - 0xff
      12'hD84: dout  = 8'b11101110; // 3460 : 238 - 0xee
      12'hD85: dout  = 8'b11101110; // 3461 : 238 - 0xee
      12'hD86: dout  = 8'b11111100; // 3462 : 252 - 0xfc
      12'hD87: dout  = 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout  = 8'b00000000; // 3464 :   0 - 0x0 -- plane 1
      12'hD89: dout  = 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout  = 8'b01111100; // 3466 : 124 - 0x7c
      12'hD8B: dout  = 8'b11111110; // 3467 : 254 - 0xfe
      12'hD8C: dout  = 8'b11101110; // 3468 : 238 - 0xee
      12'hD8D: dout  = 8'b11101110; // 3469 : 238 - 0xee
      12'hD8E: dout  = 8'b01111100; // 3470 : 124 - 0x7c
      12'hD8F: dout  = 8'b11111110; // 3471 : 254 - 0xfe
      12'hD90: dout  = 8'b11111111; // 3472 : 255 - 0xff -- Background 0xd9
      12'hD91: dout  = 8'b11111111; // 3473 : 255 - 0xff
      12'hD92: dout  = 8'b11111111; // 3474 : 255 - 0xff
      12'hD93: dout  = 8'b11111111; // 3475 : 255 - 0xff
      12'hD94: dout  = 8'b11101110; // 3476 : 238 - 0xee
      12'hD95: dout  = 8'b11101110; // 3477 : 238 - 0xee
      12'hD96: dout  = 8'b11101110; // 3478 : 238 - 0xee
      12'hD97: dout  = 8'b11101110; // 3479 : 238 - 0xee
      12'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout  = 8'b00000000; // 3481 :   0 - 0x0
      12'hD9A: dout  = 8'b01111100; // 3482 : 124 - 0x7c
      12'hD9B: dout  = 8'b11111110; // 3483 : 254 - 0xfe
      12'hD9C: dout  = 8'b11101110; // 3484 : 238 - 0xee
      12'hD9D: dout  = 8'b11101110; // 3485 : 238 - 0xee
      12'hD9E: dout  = 8'b11101110; // 3486 : 238 - 0xee
      12'hD9F: dout  = 8'b11101110; // 3487 : 238 - 0xee
      12'hDA0: dout  = 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xda
      12'hDA1: dout  = 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout  = 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout  = 8'b10000000; // 3491 : 128 - 0x80
      12'hDA4: dout  = 8'b00000000; // 3492 :   0 - 0x0
      12'hDA5: dout  = 8'b00000000; // 3493 :   0 - 0x0
      12'hDA6: dout  = 8'b00000100; // 3494 :   4 - 0x4
      12'hDA7: dout  = 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout  = 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout  = 8'b00100000; // 3497 :  32 - 0x20
      12'hDAA: dout  = 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout  = 8'b00000010; // 3499 :   2 - 0x2
      12'hDAC: dout  = 8'b00000000; // 3500 :   0 - 0x0
      12'hDAD: dout  = 8'b00100000; // 3501 :  32 - 0x20
      12'hDAE: dout  = 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout  = 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xdb
      12'hDB1: dout  = 8'b00000100; // 3505 :   4 - 0x4
      12'hDB2: dout  = 8'b00000000; // 3506 :   0 - 0x0
      12'hDB3: dout  = 8'b00010001; // 3507 :  17 - 0x11
      12'hDB4: dout  = 8'b00000000; // 3508 :   0 - 0x0
      12'hDB5: dout  = 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout  = 8'b00000000; // 3510 :   0 - 0x0
      12'hDB7: dout  = 8'b00100000; // 3511 :  32 - 0x20
      12'hDB8: dout  = 8'b00100000; // 3512 :  32 - 0x20 -- plane 1
      12'hDB9: dout  = 8'b00000000; // 3513 :   0 - 0x0
      12'hDBA: dout  = 8'b00000000; // 3514 :   0 - 0x0
      12'hDBB: dout  = 8'b00000000; // 3515 :   0 - 0x0
      12'hDBC: dout  = 8'b10000000; // 3516 : 128 - 0x80
      12'hDBD: dout  = 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout  = 8'b00000100; // 3518 :   4 - 0x4
      12'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xdc
      12'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout  = 8'b00000000; // 3522 :   0 - 0x0
      12'hDC3: dout  = 8'b00100000; // 3523 :  32 - 0x20
      12'hDC4: dout  = 8'b00000000; // 3524 :   0 - 0x0
      12'hDC5: dout  = 8'b00000000; // 3525 :   0 - 0x0
      12'hDC6: dout  = 8'b00000000; // 3526 :   0 - 0x0
      12'hDC7: dout  = 8'b00000100; // 3527 :   4 - 0x4
      12'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0 -- plane 1
      12'hDC9: dout  = 8'b00001000; // 3529 :   8 - 0x8
      12'hDCA: dout  = 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout  = 8'b00000000; // 3531 :   0 - 0x0
      12'hDCC: dout  = 8'b00000010; // 3532 :   2 - 0x2
      12'hDCD: dout  = 8'b00000000; // 3533 :   0 - 0x0
      12'hDCE: dout  = 8'b01000000; // 3534 :  64 - 0x40
      12'hDCF: dout  = 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout  = 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xdd
      12'hDD1: dout  = 8'b00000000; // 3537 :   0 - 0x0
      12'hDD2: dout  = 8'b00010001; // 3538 :  17 - 0x11
      12'hDD3: dout  = 8'b00000000; // 3539 :   0 - 0x0
      12'hDD4: dout  = 8'b00000000; // 3540 :   0 - 0x0
      12'hDD5: dout  = 8'b10000000; // 3541 : 128 - 0x80
      12'hDD6: dout  = 8'b00000000; // 3542 :   0 - 0x0
      12'hDD7: dout  = 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout  = 8'b00000000; // 3544 :   0 - 0x0 -- plane 1
      12'hDD9: dout  = 8'b01000000; // 3545 :  64 - 0x40
      12'hDDA: dout  = 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout  = 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout  = 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout  = 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout  = 8'b00000010; // 3550 :   2 - 0x2
      12'hDDF: dout  = 8'b00100000; // 3551 :  32 - 0x20
      12'hDE0: dout  = 8'b10110011; // 3552 : 179 - 0xb3 -- Background 0xde
      12'hDE1: dout  = 8'b10110011; // 3553 : 179 - 0xb3
      12'hDE2: dout  = 8'b10110011; // 3554 : 179 - 0xb3
      12'hDE3: dout  = 8'b10110011; // 3555 : 179 - 0xb3
      12'hDE4: dout  = 8'b10110000; // 3556 : 176 - 0xb0
      12'hDE5: dout  = 8'b10101111; // 3557 : 175 - 0xaf
      12'hDE6: dout  = 8'b10011111; // 3558 : 159 - 0x9f
      12'hDE7: dout  = 8'b11000000; // 3559 : 192 - 0xc0
      12'hDE8: dout  = 8'b00111110; // 3560 :  62 - 0x3e -- plane 1
      12'hDE9: dout  = 8'b00111111; // 3561 :  63 - 0x3f
      12'hDEA: dout  = 8'b00111110; // 3562 :  62 - 0x3e
      12'hDEB: dout  = 8'b00111100; // 3563 :  60 - 0x3c
      12'hDEC: dout  = 8'b00111111; // 3564 :  63 - 0x3f
      12'hDED: dout  = 8'b00110000; // 3565 :  48 - 0x30
      12'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout  = 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout  = 8'b11101101; // 3568 : 237 - 0xed -- Background 0xdf
      12'hDF1: dout  = 8'b11001101; // 3569 : 205 - 0xcd
      12'hDF2: dout  = 8'b11001101; // 3570 : 205 - 0xcd
      12'hDF3: dout  = 8'b00001101; // 3571 :  13 - 0xd
      12'hDF4: dout  = 8'b00001101; // 3572 :  13 - 0xd
      12'hDF5: dout  = 8'b11111101; // 3573 : 253 - 0xfd
      12'hDF6: dout  = 8'b11111101; // 3574 : 253 - 0xfd
      12'hDF7: dout  = 8'b00000011; // 3575 :   3 - 0x3
      12'hDF8: dout  = 8'b00010000; // 3576 :  16 - 0x10 -- plane 1
      12'hDF9: dout  = 8'b10110000; // 3577 : 176 - 0xb0
      12'hDFA: dout  = 8'b00110000; // 3578 :  48 - 0x30
      12'hDFB: dout  = 8'b11110000; // 3579 : 240 - 0xf0
      12'hDFC: dout  = 8'b11110000; // 3580 : 240 - 0xf0
      12'hDFD: dout  = 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout  = 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout  = 8'b11101110; // 3584 : 238 - 0xee -- Background 0xe0
      12'hE01: dout  = 8'b11101110; // 3585 : 238 - 0xee
      12'hE02: dout  = 8'b11101110; // 3586 : 238 - 0xee
      12'hE03: dout  = 8'b11101110; // 3587 : 238 - 0xee
      12'hE04: dout  = 8'b11111110; // 3588 : 254 - 0xfe
      12'hE05: dout  = 8'b11111100; // 3589 : 252 - 0xfc
      12'hE06: dout  = 8'b11000001; // 3590 : 193 - 0xc1
      12'hE07: dout  = 8'b11111111; // 3591 : 255 - 0xff
      12'hE08: dout  = 8'b11101110; // 3592 : 238 - 0xee -- plane 1
      12'hE09: dout  = 8'b11101110; // 3593 : 238 - 0xee
      12'hE0A: dout  = 8'b11101110; // 3594 : 238 - 0xee
      12'hE0B: dout  = 8'b11101110; // 3595 : 238 - 0xee
      12'hE0C: dout  = 8'b11111110; // 3596 : 254 - 0xfe
      12'hE0D: dout  = 8'b01111100; // 3597 : 124 - 0x7c
      12'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout  = 8'b11111011; // 3600 : 251 - 0xfb -- Background 0xe1
      12'hE11: dout  = 8'b11111011; // 3601 : 251 - 0xfb
      12'hE12: dout  = 8'b11111011; // 3602 : 251 - 0xfb
      12'hE13: dout  = 8'b11111011; // 3603 : 251 - 0xfb
      12'hE14: dout  = 8'b11111111; // 3604 : 255 - 0xff
      12'hE15: dout  = 8'b11111101; // 3605 : 253 - 0xfd
      12'hE16: dout  = 8'b11000001; // 3606 : 193 - 0xc1
      12'hE17: dout  = 8'b11111111; // 3607 : 255 - 0xff
      12'hE18: dout  = 8'b00111000; // 3608 :  56 - 0x38 -- plane 1
      12'hE19: dout  = 8'b00111000; // 3609 :  56 - 0x38
      12'hE1A: dout  = 8'b00111000; // 3610 :  56 - 0x38
      12'hE1B: dout  = 8'b00111000; // 3611 :  56 - 0x38
      12'hE1C: dout  = 8'b01111100; // 3612 : 124 - 0x7c
      12'hE1D: dout  = 8'b01111100; // 3613 : 124 - 0x7c
      12'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout  = 8'b11111100; // 3616 : 252 - 0xfc -- Background 0xe2
      12'hE21: dout  = 8'b11100001; // 3617 : 225 - 0xe1
      12'hE22: dout  = 8'b11101111; // 3618 : 239 - 0xef
      12'hE23: dout  = 8'b11101111; // 3619 : 239 - 0xef
      12'hE24: dout  = 8'b11111111; // 3620 : 255 - 0xff
      12'hE25: dout  = 8'b11111110; // 3621 : 254 - 0xfe
      12'hE26: dout  = 8'b10000000; // 3622 : 128 - 0x80
      12'hE27: dout  = 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout  = 8'b11111100; // 3624 : 252 - 0xfc -- plane 1
      12'hE29: dout  = 8'b11100000; // 3625 : 224 - 0xe0
      12'hE2A: dout  = 8'b11100000; // 3626 : 224 - 0xe0
      12'hE2B: dout  = 8'b11100000; // 3627 : 224 - 0xe0
      12'hE2C: dout  = 8'b11111110; // 3628 : 254 - 0xfe
      12'hE2D: dout  = 8'b11111110; // 3629 : 254 - 0xfe
      12'hE2E: dout  = 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout  = 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout  = 8'b11101110; // 3632 : 238 - 0xee -- Background 0xe3
      12'hE31: dout  = 8'b11111110; // 3633 : 254 - 0xfe
      12'hE32: dout  = 8'b11111110; // 3634 : 254 - 0xfe
      12'hE33: dout  = 8'b11111110; // 3635 : 254 - 0xfe
      12'hE34: dout  = 8'b11111110; // 3636 : 254 - 0xfe
      12'hE35: dout  = 8'b11111100; // 3637 : 252 - 0xfc
      12'hE36: dout  = 8'b11000001; // 3638 : 193 - 0xc1
      12'hE37: dout  = 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout  = 8'b00001110; // 3640 :  14 - 0xe -- plane 1
      12'hE39: dout  = 8'b00001110; // 3641 :  14 - 0xe
      12'hE3A: dout  = 8'b00001110; // 3642 :  14 - 0xe
      12'hE3B: dout  = 8'b11101110; // 3643 : 238 - 0xee
      12'hE3C: dout  = 8'b11111110; // 3644 : 254 - 0xfe
      12'hE3D: dout  = 8'b01111100; // 3645 : 124 - 0x7c
      12'hE3E: dout  = 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout  = 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout  = 8'b11101110; // 3648 : 238 - 0xee -- Background 0xe4
      12'hE41: dout  = 8'b11101110; // 3649 : 238 - 0xee
      12'hE42: dout  = 8'b11111110; // 3650 : 254 - 0xfe
      12'hE43: dout  = 8'b11111110; // 3651 : 254 - 0xfe
      12'hE44: dout  = 8'b10001110; // 3652 : 142 - 0x8e
      12'hE45: dout  = 8'b11111110; // 3653 : 254 - 0xfe
      12'hE46: dout  = 8'b11111000; // 3654 : 248 - 0xf8
      12'hE47: dout  = 8'b11111111; // 3655 : 255 - 0xff
      12'hE48: dout  = 8'b11101110; // 3656 : 238 - 0xee -- plane 1
      12'hE49: dout  = 8'b11101110; // 3657 : 238 - 0xee
      12'hE4A: dout  = 8'b11111110; // 3658 : 254 - 0xfe
      12'hE4B: dout  = 8'b11111110; // 3659 : 254 - 0xfe
      12'hE4C: dout  = 8'b00001110; // 3660 :  14 - 0xe
      12'hE4D: dout  = 8'b00001110; // 3661 :  14 - 0xe
      12'hE4E: dout  = 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout  = 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout  = 8'b10001110; // 3664 : 142 - 0x8e -- Background 0xe5
      12'hE51: dout  = 8'b11111110; // 3665 : 254 - 0xfe
      12'hE52: dout  = 8'b11111110; // 3666 : 254 - 0xfe
      12'hE53: dout  = 8'b11111110; // 3667 : 254 - 0xfe
      12'hE54: dout  = 8'b11111110; // 3668 : 254 - 0xfe
      12'hE55: dout  = 8'b11111100; // 3669 : 252 - 0xfc
      12'hE56: dout  = 8'b11000001; // 3670 : 193 - 0xc1
      12'hE57: dout  = 8'b11111111; // 3671 : 255 - 0xff
      12'hE58: dout  = 8'b00001110; // 3672 :  14 - 0xe -- plane 1
      12'hE59: dout  = 8'b00001110; // 3673 :  14 - 0xe
      12'hE5A: dout  = 8'b00001110; // 3674 :  14 - 0xe
      12'hE5B: dout  = 8'b11101110; // 3675 : 238 - 0xee
      12'hE5C: dout  = 8'b11111110; // 3676 : 254 - 0xfe
      12'hE5D: dout  = 8'b01111100; // 3677 : 124 - 0x7c
      12'hE5E: dout  = 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout  = 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout  = 8'b11101110; // 3680 : 238 - 0xee -- Background 0xe6
      12'hE61: dout  = 8'b11101110; // 3681 : 238 - 0xee
      12'hE62: dout  = 8'b11101110; // 3682 : 238 - 0xee
      12'hE63: dout  = 8'b11101110; // 3683 : 238 - 0xee
      12'hE64: dout  = 8'b11111110; // 3684 : 254 - 0xfe
      12'hE65: dout  = 8'b11111100; // 3685 : 252 - 0xfc
      12'hE66: dout  = 8'b11000001; // 3686 : 193 - 0xc1
      12'hE67: dout  = 8'b11111111; // 3687 : 255 - 0xff
      12'hE68: dout  = 8'b11101110; // 3688 : 238 - 0xee -- plane 1
      12'hE69: dout  = 8'b11101110; // 3689 : 238 - 0xee
      12'hE6A: dout  = 8'b11101110; // 3690 : 238 - 0xee
      12'hE6B: dout  = 8'b11101110; // 3691 : 238 - 0xee
      12'hE6C: dout  = 8'b11111110; // 3692 : 254 - 0xfe
      12'hE6D: dout  = 8'b01111100; // 3693 : 124 - 0x7c
      12'hE6E: dout  = 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout  = 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout  = 8'b11111101; // 3696 : 253 - 0xfd -- Background 0xe7
      12'hE71: dout  = 8'b11111101; // 3697 : 253 - 0xfd
      12'hE72: dout  = 8'b11111001; // 3698 : 249 - 0xf9
      12'hE73: dout  = 8'b11111011; // 3699 : 251 - 0xfb
      12'hE74: dout  = 8'b11111011; // 3700 : 251 - 0xfb
      12'hE75: dout  = 8'b11111011; // 3701 : 251 - 0xfb
      12'hE76: dout  = 8'b11100011; // 3702 : 227 - 0xe3
      12'hE77: dout  = 8'b11111111; // 3703 : 255 - 0xff
      12'hE78: dout  = 8'b00011100; // 3704 :  28 - 0x1c -- plane 1
      12'hE79: dout  = 8'b00011100; // 3705 :  28 - 0x1c
      12'hE7A: dout  = 8'b00111000; // 3706 :  56 - 0x38
      12'hE7B: dout  = 8'b00111000; // 3707 :  56 - 0x38
      12'hE7C: dout  = 8'b00111000; // 3708 :  56 - 0x38
      12'hE7D: dout  = 8'b00111000; // 3709 :  56 - 0x38
      12'hE7E: dout  = 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout  = 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout  = 8'b11101110; // 3712 : 238 - 0xee -- Background 0xe8
      12'hE81: dout  = 8'b11101110; // 3713 : 238 - 0xee
      12'hE82: dout  = 8'b11101110; // 3714 : 238 - 0xee
      12'hE83: dout  = 8'b11101110; // 3715 : 238 - 0xee
      12'hE84: dout  = 8'b11111110; // 3716 : 254 - 0xfe
      12'hE85: dout  = 8'b11111100; // 3717 : 252 - 0xfc
      12'hE86: dout  = 8'b11000001; // 3718 : 193 - 0xc1
      12'hE87: dout  = 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout  = 8'b11101110; // 3720 : 238 - 0xee -- plane 1
      12'hE89: dout  = 8'b11101110; // 3721 : 238 - 0xee
      12'hE8A: dout  = 8'b11101110; // 3722 : 238 - 0xee
      12'hE8B: dout  = 8'b11101110; // 3723 : 238 - 0xee
      12'hE8C: dout  = 8'b11111110; // 3724 : 254 - 0xfe
      12'hE8D: dout  = 8'b01111100; // 3725 : 124 - 0x7c
      12'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout  = 8'b11111110; // 3728 : 254 - 0xfe -- Background 0xe9
      12'hE91: dout  = 8'b11111110; // 3729 : 254 - 0xfe
      12'hE92: dout  = 8'b11001110; // 3730 : 206 - 0xce
      12'hE93: dout  = 8'b11111110; // 3731 : 254 - 0xfe
      12'hE94: dout  = 8'b11111110; // 3732 : 254 - 0xfe
      12'hE95: dout  = 8'b11111100; // 3733 : 252 - 0xfc
      12'hE96: dout  = 8'b11000001; // 3734 : 193 - 0xc1
      12'hE97: dout  = 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout  = 8'b11111110; // 3736 : 254 - 0xfe -- plane 1
      12'hE99: dout  = 8'b01111110; // 3737 : 126 - 0x7e
      12'hE9A: dout  = 8'b00001110; // 3738 :  14 - 0xe
      12'hE9B: dout  = 8'b00001110; // 3739 :  14 - 0xe
      12'hE9C: dout  = 8'b01111110; // 3740 : 126 - 0x7e
      12'hE9D: dout  = 8'b01111100; // 3741 : 124 - 0x7c
      12'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      12'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout  = 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xea
      12'hEA1: dout  = 8'b01110000; // 3745 : 112 - 0x70
      12'hEA2: dout  = 8'b00111000; // 3746 :  56 - 0x38
      12'hEA3: dout  = 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout  = 8'b00000010; // 3748 :   2 - 0x2
      12'hEA5: dout  = 8'b00000111; // 3749 :   7 - 0x7
      12'hEA6: dout  = 8'b00000011; // 3750 :   3 - 0x3
      12'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout  = 8'b00000000; // 3752 :   0 - 0x0 -- plane 1
      12'hEA9: dout  = 8'b01110000; // 3753 : 112 - 0x70
      12'hEAA: dout  = 8'b00111000; // 3754 :  56 - 0x38
      12'hEAB: dout  = 8'b00000000; // 3755 :   0 - 0x0
      12'hEAC: dout  = 8'b00000010; // 3756 :   2 - 0x2
      12'hEAD: dout  = 8'b00000111; // 3757 :   7 - 0x7
      12'hEAE: dout  = 8'b00000011; // 3758 :   3 - 0x3
      12'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout  = 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xeb
      12'hEB1: dout  = 8'b00001100; // 3761 :  12 - 0xc
      12'hEB2: dout  = 8'b00000110; // 3762 :   6 - 0x6
      12'hEB3: dout  = 8'b00000110; // 3763 :   6 - 0x6
      12'hEB4: dout  = 8'b01100000; // 3764 :  96 - 0x60
      12'hEB5: dout  = 8'b01110000; // 3765 : 112 - 0x70
      12'hEB6: dout  = 8'b00110000; // 3766 :  48 - 0x30
      12'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout  = 8'b00000000; // 3768 :   0 - 0x0 -- plane 1
      12'hEB9: dout  = 8'b00001100; // 3769 :  12 - 0xc
      12'hEBA: dout  = 8'b00000110; // 3770 :   6 - 0x6
      12'hEBB: dout  = 8'b00000110; // 3771 :   6 - 0x6
      12'hEBC: dout  = 8'b01100000; // 3772 :  96 - 0x60
      12'hEBD: dout  = 8'b01110000; // 3773 : 112 - 0x70
      12'hEBE: dout  = 8'b00110000; // 3774 :  48 - 0x30
      12'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xec
      12'hEC1: dout  = 8'b11000000; // 3777 : 192 - 0xc0
      12'hEC2: dout  = 8'b11100000; // 3778 : 224 - 0xe0
      12'hEC3: dout  = 8'b01100000; // 3779 :  96 - 0x60
      12'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout  = 8'b00001100; // 3781 :  12 - 0xc
      12'hEC6: dout  = 8'b00001110; // 3782 :  14 - 0xe
      12'hEC7: dout  = 8'b00000110; // 3783 :   6 - 0x6
      12'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout  = 8'b11000000; // 3785 : 192 - 0xc0
      12'hECA: dout  = 8'b11100000; // 3786 : 224 - 0xe0
      12'hECB: dout  = 8'b01100000; // 3787 :  96 - 0x60
      12'hECC: dout  = 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout  = 8'b00001100; // 3789 :  12 - 0xc
      12'hECE: dout  = 8'b00001110; // 3790 :  14 - 0xe
      12'hECF: dout  = 8'b00000110; // 3791 :   6 - 0x6
      12'hED0: dout  = 8'b01100000; // 3792 :  96 - 0x60 -- Background 0xed
      12'hED1: dout  = 8'b01110000; // 3793 : 112 - 0x70
      12'hED2: dout  = 8'b00110000; // 3794 :  48 - 0x30
      12'hED3: dout  = 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout  = 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout  = 8'b00001100; // 3797 :  12 - 0xc
      12'hED6: dout  = 8'b00001110; // 3798 :  14 - 0xe
      12'hED7: dout  = 8'b00000110; // 3799 :   6 - 0x6
      12'hED8: dout  = 8'b01100000; // 3800 :  96 - 0x60 -- plane 1
      12'hED9: dout  = 8'b01110000; // 3801 : 112 - 0x70
      12'hEDA: dout  = 8'b00110000; // 3802 :  48 - 0x30
      12'hEDB: dout  = 8'b00000000; // 3803 :   0 - 0x0
      12'hEDC: dout  = 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout  = 8'b00001100; // 3805 :  12 - 0xc
      12'hEDE: dout  = 8'b00001110; // 3806 :  14 - 0xe
      12'hEDF: dout  = 8'b00000110; // 3807 :   6 - 0x6
      12'hEE0: dout  = 8'b11111111; // 3808 : 255 - 0xff -- Background 0xee
      12'hEE1: dout  = 8'b11111111; // 3809 : 255 - 0xff
      12'hEE2: dout  = 8'b10111101; // 3810 : 189 - 0xbd
      12'hEE3: dout  = 8'b11111111; // 3811 : 255 - 0xff
      12'hEE4: dout  = 8'b11111111; // 3812 : 255 - 0xff
      12'hEE5: dout  = 8'b11111011; // 3813 : 251 - 0xfb
      12'hEE6: dout  = 8'b11111111; // 3814 : 255 - 0xff
      12'hEE7: dout  = 8'b11111111; // 3815 : 255 - 0xff
      12'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0 -- plane 1
      12'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout  = 8'b01000010; // 3818 :  66 - 0x42
      12'hEEB: dout  = 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout  = 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout  = 8'b00000100; // 3821 :   4 - 0x4
      12'hEEE: dout  = 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout  = 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout  = 8'b11111111; // 3824 : 255 - 0xff -- Background 0xef
      12'hEF1: dout  = 8'b11111111; // 3825 : 255 - 0xff
      12'hEF2: dout  = 8'b11111011; // 3826 : 251 - 0xfb
      12'hEF3: dout  = 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout  = 8'b11011111; // 3828 : 223 - 0xdf
      12'hEF5: dout  = 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout  = 8'b11111111; // 3830 : 255 - 0xff
      12'hEF7: dout  = 8'b11111111; // 3831 : 255 - 0xff
      12'hEF8: dout  = 8'b00000000; // 3832 :   0 - 0x0 -- plane 1
      12'hEF9: dout  = 8'b00000000; // 3833 :   0 - 0x0
      12'hEFA: dout  = 8'b00000100; // 3834 :   4 - 0x4
      12'hEFB: dout  = 8'b00000000; // 3835 :   0 - 0x0
      12'hEFC: dout  = 8'b00100000; // 3836 :  32 - 0x20
      12'hEFD: dout  = 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout  = 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout  = 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xf0
      12'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout  = 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout  = 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b00000000; // 3856 :   0 - 0x0 -- Background 0xf1
      12'hF11: dout  = 8'b10000000; // 3857 : 128 - 0x80
      12'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout  = 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b10000000; // 3864 : 128 - 0x80 -- plane 1
      12'hF19: dout  = 8'b10000000; // 3865 : 128 - 0x80
      12'hF1A: dout  = 8'b10000000; // 3866 : 128 - 0x80
      12'hF1B: dout  = 8'b10000000; // 3867 : 128 - 0x80
      12'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout  = 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xf2
      12'hF21: dout  = 8'b11000000; // 3873 : 192 - 0xc0
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout  = 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout  = 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout  = 8'b11000000; // 3880 : 192 - 0xc0 -- plane 1
      12'hF29: dout  = 8'b11000000; // 3881 : 192 - 0xc0
      12'hF2A: dout  = 8'b11000000; // 3882 : 192 - 0xc0
      12'hF2B: dout  = 8'b11000000; // 3883 : 192 - 0xc0
      12'hF2C: dout  = 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout  = 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout  = 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout  = 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout  = 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xf3
      12'hF31: dout  = 8'b11100000; // 3889 : 224 - 0xe0
      12'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout  = 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout  = 8'b11100000; // 3896 : 224 - 0xe0 -- plane 1
      12'hF39: dout  = 8'b11100000; // 3897 : 224 - 0xe0
      12'hF3A: dout  = 8'b11100000; // 3898 : 224 - 0xe0
      12'hF3B: dout  = 8'b11100000; // 3899 : 224 - 0xe0
      12'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout  = 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout  = 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xf4
      12'hF41: dout  = 8'b11110000; // 3905 : 240 - 0xf0
      12'hF42: dout  = 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout  = 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout  = 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout  = 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout  = 8'b11110000; // 3912 : 240 - 0xf0 -- plane 1
      12'hF49: dout  = 8'b11110000; // 3913 : 240 - 0xf0
      12'hF4A: dout  = 8'b11110000; // 3914 : 240 - 0xf0
      12'hF4B: dout  = 8'b11110000; // 3915 : 240 - 0xf0
      12'hF4C: dout  = 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout  = 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xf5
      12'hF51: dout  = 8'b11111000; // 3921 : 248 - 0xf8
      12'hF52: dout  = 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout  = 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout  = 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout  = 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout  = 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout  = 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout  = 8'b11111000; // 3928 : 248 - 0xf8 -- plane 1
      12'hF59: dout  = 8'b11111000; // 3929 : 248 - 0xf8
      12'hF5A: dout  = 8'b11111000; // 3930 : 248 - 0xf8
      12'hF5B: dout  = 8'b11111000; // 3931 : 248 - 0xf8
      12'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xf6
      12'hF61: dout  = 8'b11111100; // 3937 : 252 - 0xfc
      12'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout  = 8'b11111100; // 3944 : 252 - 0xfc -- plane 1
      12'hF69: dout  = 8'b11111100; // 3945 : 252 - 0xfc
      12'hF6A: dout  = 8'b11111100; // 3946 : 252 - 0xfc
      12'hF6B: dout  = 8'b11111100; // 3947 : 252 - 0xfc
      12'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xf7
      12'hF71: dout  = 8'b11111110; // 3953 : 254 - 0xfe
      12'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout  = 8'b11111110; // 3960 : 254 - 0xfe -- plane 1
      12'hF79: dout  = 8'b11111110; // 3961 : 254 - 0xfe
      12'hF7A: dout  = 8'b11111110; // 3962 : 254 - 0xfe
      12'hF7B: dout  = 8'b11111110; // 3963 : 254 - 0xfe
      12'hF7C: dout  = 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout  = 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout  = 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf8
      12'hF81: dout  = 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout  = 8'b11111111; // 3976 : 255 - 0xff -- plane 1
      12'hF89: dout  = 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout  = 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout  = 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout  = 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout  = 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout  = 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout  = 8'b11111111; // 3984 : 255 - 0xff -- Background 0xf9
      12'hF91: dout  = 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout  = 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout  = 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout  = 8'b10000000; // 3988 : 128 - 0x80
      12'hF95: dout  = 8'b10000000; // 3989 : 128 - 0x80
      12'hF96: dout  = 8'b11000000; // 3990 : 192 - 0xc0
      12'hF97: dout  = 8'b11000000; // 3991 : 192 - 0xc0
      12'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0 -- plane 1
      12'hF99: dout  = 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout  = 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout  = 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout  = 8'b01111111; // 3996 : 127 - 0x7f
      12'hF9D: dout  = 8'b01000000; // 3997 :  64 - 0x40
      12'hF9E: dout  = 8'b01000000; // 3998 :  64 - 0x40
      12'hF9F: dout  = 8'b01000000; // 3999 :  64 - 0x40
      12'hFA0: dout  = 8'b11111111; // 4000 : 255 - 0xff -- Background 0xfa
      12'hFA1: dout  = 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout  = 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout  = 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout  = 8'b00000000; // 4008 :   0 - 0x0 -- plane 1
      12'hFA9: dout  = 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout  = 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout  = 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout  = 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout  = 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout  = 8'b11111111; // 4016 : 255 - 0xff -- Background 0xfb
      12'hFB1: dout  = 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout  = 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout  = 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout  = 8'b00000001; // 4020 :   1 - 0x1
      12'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout  = 8'b00000010; // 4022 :   2 - 0x2
      12'hFB7: dout  = 8'b00000010; // 4023 :   2 - 0x2
      12'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout  = 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout  = 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout  = 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout  = 8'b11111110; // 4028 : 254 - 0xfe
      12'hFBD: dout  = 8'b00000010; // 4029 :   2 - 0x2
      12'hFBE: dout  = 8'b00000010; // 4030 :   2 - 0x2
      12'hFBF: dout  = 8'b00000010; // 4031 :   2 - 0x2
      12'hFC0: dout  = 8'b11000000; // 4032 : 192 - 0xc0 -- Background 0xfc
      12'hFC1: dout  = 8'b11000000; // 4033 : 192 - 0xc0
      12'hFC2: dout  = 8'b10000000; // 4034 : 128 - 0x80
      12'hFC3: dout  = 8'b10000000; // 4035 : 128 - 0x80
      12'hFC4: dout  = 8'b11000000; // 4036 : 192 - 0xc0
      12'hFC5: dout  = 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout  = 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout  = 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout  = 8'b01000000; // 4040 :  64 - 0x40 -- plane 1
      12'hFC9: dout  = 8'b01000000; // 4041 :  64 - 0x40
      12'hFCA: dout  = 8'b01000000; // 4042 :  64 - 0x40
      12'hFCB: dout  = 8'b01111111; // 4043 : 127 - 0x7f
      12'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Background 0xfd
      12'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout  = 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout  = 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout  = 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout  = 8'b00000000; // 4056 :   0 - 0x0 -- plane 1
      12'hFD9: dout  = 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout  = 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout  = 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout  = 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout  = 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout  = 8'b00000010; // 4064 :   2 - 0x2 -- Background 0xfe
      12'hFE1: dout  = 8'b00000010; // 4065 :   2 - 0x2
      12'hFE2: dout  = 8'b00000000; // 4066 :   0 - 0x0
      12'hFE3: dout  = 8'b00000000; // 4067 :   0 - 0x0
      12'hFE4: dout  = 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout  = 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout  = 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout  = 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout  = 8'b00000010; // 4072 :   2 - 0x2 -- plane 1
      12'hFE9: dout  = 8'b00000010; // 4073 :   2 - 0x2
      12'hFEA: dout  = 8'b00000010; // 4074 :   2 - 0x2
      12'hFEB: dout  = 8'b11111110; // 4075 : 254 - 0xfe
      12'hFEC: dout  = 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout  = 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout  = 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout  = 8'b11111111; // 4080 : 255 - 0xff -- Background 0xff
      12'hFF1: dout  = 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout  = 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout  = 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout  = 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout  = 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout  = 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout  = 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout  = 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout  = 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout  = 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout  = 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout  = 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
