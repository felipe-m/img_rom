--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables

---  Original memory dump file name: smario_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_SMARIO_color1 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_SMARIO_color1;

architecture BEHAVIORAL of ROM_PTABLE_SMARIO_color1 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant nametable_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00000000", --    0 -  0x0  :    0 - 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00011111", --    4 -  0x4  :   31 - 0x1f
    "00111111", --    5 -  0x5  :   63 - 0x3f
    "00111111", --    6 -  0x6  :   63 - 0x3f
    "01111111", --    7 -  0x7  :  127 - 0x7f
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00100000", --    9 -  0x9  :   32 - 0x20
    "01100000", --   10 -  0xa  :   96 - 0x60
    "00000000", --   11 -  0xb  :    0 - 0x0
    "11110000", --   12 -  0xc  :  240 - 0xf0
    "11111100", --   13 -  0xd  :  252 - 0xfc
    "11111110", --   14 -  0xe  :  254 - 0xfe
    "11111110", --   15 -  0xf  :  254 - 0xfe
    "01111111", --   16 - 0x10  :  127 - 0x7f
    "01111111", --   17 - 0x11  :  127 - 0x7f
    "00011111", --   18 - 0x12  :   31 - 0x1f
    "00000111", --   19 - 0x13  :    7 - 0x7
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00011110", --   21 - 0x15  :   30 - 0x1e
    "00111111", --   22 - 0x16  :   63 - 0x3f
    "01111111", --   23 - 0x17  :  127 - 0x7f
    "11111100", --   24 - 0x18  :  252 - 0xfc
    "11111100", --   25 - 0x19  :  252 - 0xfc
    "11111000", --   26 - 0x1a  :  248 - 0xf8
    "11000000", --   27 - 0x1b  :  192 - 0xc0
    "11000010", --   28 - 0x1c  :  194 - 0xc2
    "01100111", --   29 - 0x1d  :  103 - 0x67
    "00101111", --   30 - 0x1e  :   47 - 0x2f
    "00110111", --   31 - 0x1f  :   55 - 0x37
    "01111111", --   32 - 0x20  :  127 - 0x7f
    "01111110", --   33 - 0x21  :  126 - 0x7e
    "11111100", --   34 - 0x22  :  252 - 0xfc
    "11110000", --   35 - 0x23  :  240 - 0xf0
    "11111000", --   36 - 0x24  :  248 - 0xf8
    "11111000", --   37 - 0x25  :  248 - 0xf8
    "11110000", --   38 - 0x26  :  240 - 0xf0
    "01110000", --   39 - 0x27  :  112 - 0x70
    "00110111", --   40 - 0x28  :   55 - 0x37
    "00110110", --   41 - 0x29  :   54 - 0x36
    "01011100", --   42 - 0x2a  :   92 - 0x5c
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000001", --   45 - 0x2d  :    1 - 0x1
    "00000011", --   46 - 0x2e  :    3 - 0x3
    "00011111", --   47 - 0x2f  :   31 - 0x1f
    "00001000", --   48 - 0x30  :    8 - 0x8
    "00100100", --   49 - 0x31  :   36 - 0x24
    "11100011", --   50 - 0x32  :  227 - 0xe3
    "11110000", --   51 - 0x33  :  240 - 0xf0
    "11111000", --   52 - 0x34  :  248 - 0xf8
    "01110000", --   53 - 0x35  :  112 - 0x70
    "01110000", --   54 - 0x36  :  112 - 0x70
    "00111000", --   55 - 0x37  :   56 - 0x38
    "00011111", --   56 - 0x38  :   31 - 0x1f
    "00011111", --   57 - 0x39  :   31 - 0x1f
    "00011111", --   58 - 0x3a  :   31 - 0x1f
    "00011111", --   59 - 0x3b  :   31 - 0x1f
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00001111", --   70 - 0x46  :   15 - 0xf
    "00011111", --   71 - 0x47  :   31 - 0x1f
    "00000000", --   72 - 0x48  :    0 - 0x0
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00010000", --   75 - 0x4b  :   16 - 0x10
    "00110000", --   76 - 0x4c  :   48 - 0x30
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "11111000", --   78 - 0x4e  :  248 - 0xf8
    "11111110", --   79 - 0x4f  :  254 - 0xfe
    "00011111", --   80 - 0x50  :   31 - 0x1f
    "00111111", --   81 - 0x51  :   63 - 0x3f
    "00111111", --   82 - 0x52  :   63 - 0x3f
    "00011111", --   83 - 0x53  :   31 - 0x1f
    "00000111", --   84 - 0x54  :    7 - 0x7
    "00001000", --   85 - 0x55  :    8 - 0x8
    "00010111", --   86 - 0x56  :   23 - 0x17
    "00010111", --   87 - 0x57  :   23 - 0x17
    "11111111", --   88 - 0x58  :  255 - 0xff
    "11111111", --   89 - 0x59  :  255 - 0xff
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111110", --   91 - 0x5b  :  254 - 0xfe
    "11111100", --   92 - 0x5c  :  252 - 0xfc
    "11100000", --   93 - 0x5d  :  224 - 0xe0
    "01000000", --   94 - 0x5e  :   64 - 0x40
    "10100000", --   95 - 0x5f  :  160 - 0xa0
    "00110111", --   96 - 0x60  :   55 - 0x37
    "00100111", --   97 - 0x61  :   39 - 0x27
    "00100011", --   98 - 0x62  :   35 - 0x23
    "00000011", --   99 - 0x63  :    3 - 0x3
    "00000001", --  100 - 0x64  :    1 - 0x1
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11001100", --  104 - 0x68  :  204 - 0xcc
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111111", --  106 - 0x6a  :  255 - 0xff
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111111", --  108 - 0x6c  :  255 - 0xff
    "01110000", --  109 - 0x6d  :  112 - 0x70
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00001000", --  111 - 0x6f  :    8 - 0x8
    "11110000", --  112 - 0x70  :  240 - 0xf0
    "11110000", --  113 - 0x71  :  240 - 0xf0
    "11110000", --  114 - 0x72  :  240 - 0xf0
    "11110000", --  115 - 0x73  :  240 - 0xf0
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "10000000", --  118 - 0x76  :  128 - 0x80
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00010000", --  120 - 0x78  :   16 - 0x10
    "01100000", --  121 - 0x79  :   96 - 0x60
    "10000000", --  122 - 0x7a  :  128 - 0x80
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "01111000", --  124 - 0x7c  :  120 - 0x78
    "01111000", --  125 - 0x7d  :  120 - 0x78
    "01111110", --  126 - 0x7e  :  126 - 0x7e
    "01111110", --  127 - 0x7f  :  126 - 0x7e
    "00000000", --  128 - 0x80  :    0 - 0x0
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00011111", --  133 - 0x85  :   31 - 0x1f
    "00111111", --  134 - 0x86  :   63 - 0x3f
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00100000", --  138 - 0x8a  :   32 - 0x20
    "01100000", --  139 - 0x8b  :   96 - 0x60
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "11110000", --  141 - 0x8d  :  240 - 0xf0
    "11111100", --  142 - 0x8e  :  252 - 0xfc
    "11111110", --  143 - 0x8f  :  254 - 0xfe
    "01111111", --  144 - 0x90  :  127 - 0x7f
    "01111111", --  145 - 0x91  :  127 - 0x7f
    "00111111", --  146 - 0x92  :   63 - 0x3f
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00010110", --  149 - 0x95  :   22 - 0x16
    "00101111", --  150 - 0x96  :   47 - 0x2f
    "00101111", --  151 - 0x97  :   47 - 0x2f
    "11111110", --  152 - 0x98  :  254 - 0xfe
    "11111100", --  153 - 0x99  :  252 - 0xfc
    "11111100", --  154 - 0x9a  :  252 - 0xfc
    "11111000", --  155 - 0x9b  :  248 - 0xf8
    "11000000", --  156 - 0x9c  :  192 - 0xc0
    "01100000", --  157 - 0x9d  :   96 - 0x60
    "00100000", --  158 - 0x9e  :   32 - 0x20
    "00110000", --  159 - 0x9f  :   48 - 0x30
    "00101111", --  160 - 0xa0  :   47 - 0x2f
    "00101111", --  161 - 0xa1  :   47 - 0x2f
    "00101111", --  162 - 0xa2  :   47 - 0x2f
    "00001111", --  163 - 0xa3  :   15 - 0xf
    "00000111", --  164 - 0xa4  :    7 - 0x7
    "00000011", --  165 - 0xa5  :    3 - 0x3
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00010000", --  168 - 0xa8  :   16 - 0x10
    "11110000", --  169 - 0xa9  :  240 - 0xf0
    "11110000", --  170 - 0xaa  :  240 - 0xf0
    "11110000", --  171 - 0xab  :  240 - 0xf0
    "11110000", --  172 - 0xac  :  240 - 0xf0
    "11100000", --  173 - 0xad  :  224 - 0xe0
    "11000000", --  174 - 0xae  :  192 - 0xc0
    "11100000", --  175 - 0xaf  :  224 - 0xe0
    "00000001", --  176 - 0xb0  :    1 - 0x1
    "00000011", --  177 - 0xb1  :    3 - 0x3
    "00000001", --  178 - 0xb2  :    1 - 0x1
    "00000100", --  179 - 0xb3  :    4 - 0x4
    "00000111", --  180 - 0xb4  :    7 - 0x7
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00001111", --  182 - 0xb6  :   15 - 0xf
    "00000011", --  183 - 0xb7  :    3 - 0x3
    "11111000", --  184 - 0xb8  :  248 - 0xf8
    "11110000", --  185 - 0xb9  :  240 - 0xf0
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "01110000", --  187 - 0xbb  :  112 - 0x70
    "10110000", --  188 - 0xbc  :  176 - 0xb0
    "10000000", --  189 - 0xbd  :  128 - 0x80
    "11100000", --  190 - 0xbe  :  224 - 0xe0
    "11100000", --  191 - 0xbf  :  224 - 0xe0
    "00000000", --  192 - 0xc0  :    0 - 0x0
    "00110000", --  193 - 0xc1  :   48 - 0x30
    "01110000", --  194 - 0xc2  :  112 - 0x70
    "01111111", --  195 - 0xc3  :  127 - 0x7f
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11110111", --  198 - 0xc6  :  247 - 0xf7
    "11110011", --  199 - 0xc7  :  243 - 0xf3
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00011000", --  201 - 0xc9  :   24 - 0x18
    "00010000", --  202 - 0xca  :   16 - 0x10
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "11111000", --  204 - 0xcc  :  248 - 0xf8
    "11111000", --  205 - 0xcd  :  248 - 0xf8
    "11111110", --  206 - 0xce  :  254 - 0xfe
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "11100111", --  208 - 0xd0  :  231 - 0xe7
    "00001111", --  209 - 0xd1  :   15 - 0xf
    "00001111", --  210 - 0xd2  :   15 - 0xf
    "00011111", --  211 - 0xd3  :   31 - 0x1f
    "00011111", --  212 - 0xd4  :   31 - 0x1f
    "00011111", --  213 - 0xd5  :   31 - 0x1f
    "00001111", --  214 - 0xd6  :   15 - 0xf
    "00000111", --  215 - 0xd7  :    7 - 0x7
    "11111111", --  216 - 0xd8  :  255 - 0xff
    "11111110", --  217 - 0xd9  :  254 - 0xfe
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "11000110", --  219 - 0xdb  :  198 - 0xc6
    "10001110", --  220 - 0xdc  :  142 - 0x8e
    "11101110", --  221 - 0xdd  :  238 - 0xee
    "11111111", --  222 - 0xde  :  255 - 0xff
    "11111111", --  223 - 0xdf  :  255 - 0xff
    "00000011", --  224 - 0xe0  :    3 - 0x3
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00001110", --  227 - 0xe3  :   14 - 0xe
    "00000111", --  228 - 0xe4  :    7 - 0x7
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00111111", --  230 - 0xe6  :   63 - 0x3f
    "00111111", --  231 - 0xe7  :   63 - 0x3f
    "11111111", --  232 - 0xe8  :  255 - 0xff
    "01111111", --  233 - 0xe9  :  127 - 0x7f
    "00111111", --  234 - 0xea  :   63 - 0x3f
    "00001110", --  235 - 0xeb  :   14 - 0xe
    "11000000", --  236 - 0xec  :  192 - 0xc0
    "11000000", --  237 - 0xed  :  192 - 0xc0
    "11100000", --  238 - 0xee  :  224 - 0xe0
    "11100000", --  239 - 0xef  :  224 - 0xe0
    "00000000", --  240 - 0xf0  :    0 - 0x0
    "10000000", --  241 - 0xf1  :  128 - 0x80
    "11001000", --  242 - 0xf2  :  200 - 0xc8
    "11111110", --  243 - 0xf3  :  254 - 0xfe
    "01111111", --  244 - 0xf4  :  127 - 0x7f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00011110", --  246 - 0xf6  :   30 - 0x1e
    "00001110", --  247 - 0xf7  :   14 - 0xe
    "11100000", --  248 - 0xf8  :  224 - 0xe0
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00011111", --  262 - 0x106  :   31 - 0x1f
    "00111111", --  263 - 0x107  :   63 - 0x3f
    "00001110", --  264 - 0x108  :   14 - 0xe
    "00011111", --  265 - 0x109  :   31 - 0x1f
    "00011111", --  266 - 0x10a  :   31 - 0x1f
    "00011111", --  267 - 0x10b  :   31 - 0x1f
    "00011111", --  268 - 0x10c  :   31 - 0x1f
    "00000011", --  269 - 0x10d  :    3 - 0x3
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "00111111", --  272 - 0x110  :   63 - 0x3f
    "00111111", --  273 - 0x111  :   63 - 0x3f
    "01111111", --  274 - 0x112  :  127 - 0x7f
    "01111111", --  275 - 0x113  :  127 - 0x7f
    "00011111", --  276 - 0x114  :   31 - 0x1f
    "00000000", --  277 - 0x115  :    0 - 0x0
    "01111110", --  278 - 0x116  :  126 - 0x7e
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111111", --  280 - 0x118  :  255 - 0xff
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11111110", --  282 - 0x11a  :  254 - 0xfe
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111110", --  284 - 0x11c  :  254 - 0xfe
    "11011110", --  285 - 0x11d  :  222 - 0xde
    "01011100", --  286 - 0x11e  :   92 - 0x5c
    "01101100", --  287 - 0x11f  :  108 - 0x6c
    "11111111", --  288 - 0x120  :  255 - 0xff
    "11111111", --  289 - 0x121  :  255 - 0xff
    "11111110", --  290 - 0x122  :  254 - 0xfe
    "11111100", --  291 - 0x123  :  252 - 0xfc
    "11111000", --  292 - 0x124  :  248 - 0xf8
    "10110000", --  293 - 0x125  :  176 - 0xb0
    "01100000", --  294 - 0x126  :   96 - 0x60
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00101000", --  296 - 0x128  :   40 - 0x28
    "00110000", --  297 - 0x129  :   48 - 0x30
    "00011000", --  298 - 0x12a  :   24 - 0x18
    "01000000", --  299 - 0x12b  :   64 - 0x40
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000001", --  301 - 0x12d  :    1 - 0x1
    "00000011", --  302 - 0x12e  :    3 - 0x3
    "00001111", --  303 - 0x12f  :   15 - 0xf
    "00010000", --  304 - 0x130  :   16 - 0x10
    "11101100", --  305 - 0x131  :  236 - 0xec
    "11100011", --  306 - 0x132  :  227 - 0xe3
    "11100000", --  307 - 0x133  :  224 - 0xe0
    "11100000", --  308 - 0x134  :  224 - 0xe0
    "11100000", --  309 - 0x135  :  224 - 0xe0
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "10000000", --  311 - 0x137  :  128 - 0x80
    "00001111", --  312 - 0x138  :   15 - 0xf
    "00001111", --  313 - 0x139  :   15 - 0xf
    "00001111", --  314 - 0x13a  :   15 - 0xf
    "00001111", --  315 - 0x13b  :   15 - 0xf
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00011111", --  320 - 0x140  :   31 - 0x1f
    "00111111", --  321 - 0x141  :   63 - 0x3f
    "00111111", --  322 - 0x142  :   63 - 0x3f
    "00011111", --  323 - 0x143  :   31 - 0x1f
    "00000111", --  324 - 0x144  :    7 - 0x7
    "00001001", --  325 - 0x145  :    9 - 0x9
    "00010011", --  326 - 0x146  :   19 - 0x13
    "00010111", --  327 - 0x147  :   23 - 0x17
    "11111111", --  328 - 0x148  :  255 - 0xff
    "11111111", --  329 - 0x149  :  255 - 0xff
    "11111110", --  330 - 0x14a  :  254 - 0xfe
    "11111111", --  331 - 0x14b  :  255 - 0xff
    "11111110", --  332 - 0x14c  :  254 - 0xfe
    "11111100", --  333 - 0x14d  :  252 - 0xfc
    "11111000", --  334 - 0x14e  :  248 - 0xf8
    "11100000", --  335 - 0x14f  :  224 - 0xe0
    "00010111", --  336 - 0x150  :   23 - 0x17
    "00010111", --  337 - 0x151  :   23 - 0x17
    "00000011", --  338 - 0x152  :    3 - 0x3
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "11010000", --  344 - 0x158  :  208 - 0xd0
    "10010000", --  345 - 0x159  :  144 - 0x90
    "00011000", --  346 - 0x15a  :   24 - 0x18
    "00001000", --  347 - 0x15b  :    8 - 0x8
    "01000000", --  348 - 0x15c  :   64 - 0x40
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00110000", --  352 - 0x160  :   48 - 0x30
    "11110000", --  353 - 0x161  :  240 - 0xf0
    "11110000", --  354 - 0x162  :  240 - 0xf0
    "11110001", --  355 - 0x163  :  241 - 0xf1
    "11110110", --  356 - 0x164  :  246 - 0xf6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "10000100", --  358 - 0x166  :  132 - 0x84
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00011111", --  368 - 0x170  :   31 - 0x1f
    "00011111", --  369 - 0x171  :   31 - 0x1f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111110", --  371 - 0x173  :   62 - 0x3e
    "01111100", --  372 - 0x174  :  124 - 0x7c
    "01111000", --  373 - 0x175  :  120 - 0x78
    "11110000", --  374 - 0x176  :  240 - 0xf0
    "11100000", --  375 - 0x177  :  224 - 0xe0
    "10110000", --  376 - 0x178  :  176 - 0xb0
    "10010000", --  377 - 0x179  :  144 - 0x90
    "00011000", --  378 - 0x17a  :   24 - 0x18
    "00001000", --  379 - 0x17b  :    8 - 0x8
    "01000000", --  380 - 0x17c  :   64 - 0x40
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "11000000", --  384 - 0x180  :  192 - 0xc0
    "11100000", --  385 - 0x181  :  224 - 0xe0
    "11111100", --  386 - 0x182  :  252 - 0xfc
    "11111110", --  387 - 0x183  :  254 - 0xfe
    "11111111", --  388 - 0x184  :  255 - 0xff
    "01111111", --  389 - 0x185  :  127 - 0x7f
    "00000011", --  390 - 0x186  :    3 - 0x3
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00010000", --  394 - 0x18a  :   16 - 0x10
    "00111000", --  395 - 0x18b  :   56 - 0x38
    "00111110", --  396 - 0x18c  :   62 - 0x3e
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00111000", --  398 - 0x18e  :   56 - 0x38
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000000", --  400 - 0x190  :    0 - 0x0
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000111", --  403 - 0x193  :    7 - 0x7
    "00001111", --  404 - 0x194  :   15 - 0xf
    "00001111", --  405 - 0x195  :   15 - 0xf
    "00001111", --  406 - 0x196  :   15 - 0xf
    "00000011", --  407 - 0x197  :    3 - 0x3
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "11110000", --  411 - 0x19b  :  240 - 0xf0
    "11111100", --  412 - 0x19c  :  252 - 0xfc
    "11111110", --  413 - 0x19d  :  254 - 0xfe
    "11111100", --  414 - 0x19e  :  252 - 0xfc
    "11111000", --  415 - 0x19f  :  248 - 0xf8
    "00000111", --  416 - 0x1a0  :    7 - 0x7
    "00001111", --  417 - 0x1a1  :   15 - 0xf
    "00011011", --  418 - 0x1a2  :   27 - 0x1b
    "00011000", --  419 - 0x1a3  :   24 - 0x18
    "00010000", --  420 - 0x1a4  :   16 - 0x10
    "00110000", --  421 - 0x1a5  :   48 - 0x30
    "00100001", --  422 - 0x1a6  :   33 - 0x21
    "00000001", --  423 - 0x1a7  :    1 - 0x1
    "10101000", --  424 - 0x1a8  :  168 - 0xa8
    "11111100", --  425 - 0x1a9  :  252 - 0xfc
    "11111000", --  426 - 0x1aa  :  248 - 0xf8
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "11000000", --  430 - 0x1ae  :  192 - 0xc0
    "11100000", --  431 - 0x1af  :  224 - 0xe0
    "00000000", --  432 - 0x1b0  :    0 - 0x0
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00001111", --  434 - 0x1b2  :   15 - 0xf
    "00011111", --  435 - 0x1b3  :   31 - 0x1f
    "00011111", --  436 - 0x1b4  :   31 - 0x1f
    "00011111", --  437 - 0x1b5  :   31 - 0x1f
    "00000111", --  438 - 0x1b6  :    7 - 0x7
    "00111100", --  439 - 0x1b7  :   60 - 0x3c
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "11100000", --  442 - 0x1ba  :  224 - 0xe0
    "11111000", --  443 - 0x1bb  :  248 - 0xf8
    "11111100", --  444 - 0x1bc  :  252 - 0xfc
    "11111000", --  445 - 0x1bd  :  248 - 0xf8
    "11110000", --  446 - 0x1be  :  240 - 0xf0
    "11000000", --  447 - 0x1bf  :  192 - 0xc0
    "11111100", --  448 - 0x1c0  :  252 - 0xfc
    "11101101", --  449 - 0x1c1  :  237 - 0xed
    "11000000", --  450 - 0x1c2  :  192 - 0xc0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "01100000", --  453 - 0x1c5  :   96 - 0x60
    "01110000", --  454 - 0x1c6  :  112 - 0x70
    "00111000", --  455 - 0x1c7  :   56 - 0x38
    "01111110", --  456 - 0x1c8  :  126 - 0x7e
    "00011110", --  457 - 0x1c9  :   30 - 0x1e
    "00000100", --  458 - 0x1ca  :    4 - 0x4
    "00001100", --  459 - 0x1cb  :   12 - 0xc
    "00001100", --  460 - 0x1cc  :   12 - 0xc
    "00001100", --  461 - 0x1cd  :   12 - 0xc
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00001111", --  466 - 0x1d2  :   15 - 0xf
    "00011111", --  467 - 0x1d3  :   31 - 0x1f
    "00011111", --  468 - 0x1d4  :   31 - 0x1f
    "00011111", --  469 - 0x1d5  :   31 - 0x1f
    "00000111", --  470 - 0x1d6  :    7 - 0x7
    "00001101", --  471 - 0x1d7  :   13 - 0xd
    "00011110", --  472 - 0x1d8  :   30 - 0x1e
    "00011100", --  473 - 0x1d9  :   28 - 0x1c
    "00011110", --  474 - 0x1da  :   30 - 0x1e
    "00001111", --  475 - 0x1db  :   15 - 0xf
    "00000111", --  476 - 0x1dc  :    7 - 0x7
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000111", --  478 - 0x1de  :    7 - 0x7
    "00000111", --  479 - 0x1df  :    7 - 0x7
    "01100000", --  480 - 0x1e0  :   96 - 0x60
    "10010000", --  481 - 0x1e1  :  144 - 0x90
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "10000000", --  483 - 0x1e3  :  128 - 0x80
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "11100000", --  485 - 0x1e5  :  224 - 0xe0
    "11110000", --  486 - 0x1e6  :  240 - 0xf0
    "10000000", --  487 - 0x1e7  :  128 - 0x80
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "00010000", --  489 - 0x1e9  :   16 - 0x10
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "01111111", --  491 - 0x1eb  :  127 - 0x7f
    "01111111", --  492 - 0x1ec  :  127 - 0x7f
    "00111111", --  493 - 0x1ed  :   63 - 0x3f
    "00000011", --  494 - 0x1ee  :    3 - 0x3
    "00001111", --  495 - 0x1ef  :   15 - 0xf
    "00000000", --  496 - 0x1f0  :    0 - 0x0
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "11100000", --  498 - 0x1f2  :  224 - 0xe0
    "11111000", --  499 - 0x1f3  :  248 - 0xf8
    "11111100", --  500 - 0x1f4  :  252 - 0xfc
    "11111000", --  501 - 0x1f5  :  248 - 0xf8
    "10110000", --  502 - 0x1f6  :  176 - 0xb0
    "00111000", --  503 - 0x1f7  :   56 - 0x38
    "00011111", --  504 - 0x1f8  :   31 - 0x1f
    "00000111", --  505 - 0x1f9  :    7 - 0x7
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00001110", --  507 - 0x1fb  :   14 - 0xe
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "01010011", --  509 - 0x1fd  :   83 - 0x53
    "01111100", --  510 - 0x1fe  :  124 - 0x7c
    "00111100", --  511 - 0x1ff  :   60 - 0x3c
    "11111000", --  512 - 0x200  :  248 - 0xf8
    "11111000", --  513 - 0x201  :  248 - 0xf8
    "11110000", --  514 - 0x202  :  240 - 0xf0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "10000000", --  517 - 0x205  :  128 - 0x80
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000111", --  520 - 0x208  :    7 - 0x7
    "00000111", --  521 - 0x209  :    7 - 0x7
    "00000011", --  522 - 0x20a  :    3 - 0x3
    "11110111", --  523 - 0x20b  :  247 - 0xf7
    "11111111", --  524 - 0x20c  :  255 - 0xff
    "11111111", --  525 - 0x20d  :  255 - 0xff
    "11111110", --  526 - 0x20e  :  254 - 0xfe
    "11111100", --  527 - 0x20f  :  252 - 0xfc
    "00111110", --  528 - 0x210  :   62 - 0x3e
    "01111111", --  529 - 0x211  :  127 - 0x7f
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11100010", --  531 - 0x213  :  226 - 0xe2
    "01010000", --  532 - 0x214  :   80 - 0x50
    "00111000", --  533 - 0x215  :   56 - 0x38
    "01110000", --  534 - 0x216  :  112 - 0x70
    "01000000", --  535 - 0x217  :   64 - 0x40
    "11101000", --  536 - 0x218  :  232 - 0xe8
    "01110001", --  537 - 0x219  :  113 - 0x71
    "00000001", --  538 - 0x21a  :    1 - 0x1
    "01001011", --  539 - 0x21b  :   75 - 0x4b
    "00000011", --  540 - 0x21c  :    3 - 0x3
    "00000011", --  541 - 0x21d  :    3 - 0x3
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000101", --  544 - 0x220  :    5 - 0x5
    "00000011", --  545 - 0x221  :    3 - 0x3
    "00000001", --  546 - 0x222  :    1 - 0x1
    "00110000", --  547 - 0x223  :   48 - 0x30
    "00110000", --  548 - 0x224  :   48 - 0x30
    "00110000", --  549 - 0x225  :   48 - 0x30
    "00100110", --  550 - 0x226  :   38 - 0x26
    "00000100", --  551 - 0x227  :    4 - 0x4
    "11111110", --  552 - 0x228  :  254 - 0xfe
    "11111100", --  553 - 0x229  :  252 - 0xfc
    "11100000", --  554 - 0x22a  :  224 - 0xe0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000101", --  560 - 0x230  :    5 - 0x5
    "00000011", --  561 - 0x231  :    3 - 0x3
    "00000001", --  562 - 0x232  :    1 - 0x1
    "00010000", --  563 - 0x233  :   16 - 0x10
    "00110000", --  564 - 0x234  :   48 - 0x30
    "00001100", --  565 - 0x235  :   12 - 0xc
    "00011100", --  566 - 0x236  :   28 - 0x1c
    "00011000", --  567 - 0x237  :   24 - 0x18
    "11000000", --  568 - 0x238  :  192 - 0xc0
    "11100000", --  569 - 0x239  :  224 - 0xe0
    "11110000", --  570 - 0x23a  :  240 - 0xf0
    "01111000", --  571 - 0x23b  :  120 - 0x78
    "00011000", --  572 - 0x23c  :   24 - 0x18
    "00001000", --  573 - 0x23d  :    8 - 0x8
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000111", --  576 - 0x240  :    7 - 0x7
    "00001111", --  577 - 0x241  :   15 - 0xf
    "00111110", --  578 - 0x242  :   62 - 0x3e
    "01111100", --  579 - 0x243  :  124 - 0x7c
    "00110000", --  580 - 0x244  :   48 - 0x30
    "00001100", --  581 - 0x245  :   12 - 0xc
    "00011100", --  582 - 0x246  :   28 - 0x1c
    "00011000", --  583 - 0x247  :   24 - 0x18
    "01100000", --  584 - 0x248  :   96 - 0x60
    "01100000", --  585 - 0x249  :   96 - 0x60
    "01100000", --  586 - 0x24a  :   96 - 0x60
    "10000000", --  587 - 0x24b  :  128 - 0x80
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "01110011", --  592 - 0x250  :  115 - 0x73
    "11110011", --  593 - 0x251  :  243 - 0xf3
    "11110000", --  594 - 0x252  :  240 - 0xf0
    "11110100", --  595 - 0x253  :  244 - 0xf4
    "11110000", --  596 - 0x254  :  240 - 0xf0
    "11110000", --  597 - 0x255  :  240 - 0xf0
    "01110000", --  598 - 0x256  :  112 - 0x70
    "01100000", --  599 - 0x257  :   96 - 0x60
    "00000000", --  600 - 0x258  :    0 - 0x0
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00111100", --  604 - 0x25c  :   60 - 0x3c
    "00111100", --  605 - 0x25d  :   60 - 0x3c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "01111111", --  608 - 0x260  :  127 - 0x7f
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "00011111", --  610 - 0x262  :   31 - 0x1f
    "00000111", --  611 - 0x263  :    7 - 0x7
    "00001011", --  612 - 0x264  :   11 - 0xb
    "00011011", --  613 - 0x265  :   27 - 0x1b
    "00111011", --  614 - 0x266  :   59 - 0x3b
    "01111011", --  615 - 0x267  :  123 - 0x7b
    "11111100", --  616 - 0x268  :  252 - 0xfc
    "11111100", --  617 - 0x269  :  252 - 0xfc
    "11111000", --  618 - 0x26a  :  248 - 0xf8
    "11100000", --  619 - 0x26b  :  224 - 0xe0
    "11010000", --  620 - 0x26c  :  208 - 0xd0
    "11011000", --  621 - 0x26d  :  216 - 0xd8
    "11011100", --  622 - 0x26e  :  220 - 0xdc
    "11011110", --  623 - 0x26f  :  222 - 0xde
    "11000100", --  624 - 0x270  :  196 - 0xc4
    "11100000", --  625 - 0x271  :  224 - 0xe0
    "11100000", --  626 - 0x272  :  224 - 0xe0
    "01000000", --  627 - 0x273  :   64 - 0x40
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00111100", --  629 - 0x275  :   60 - 0x3c
    "00111100", --  630 - 0x276  :   60 - 0x3c
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "00011101", --  632 - 0x278  :   29 - 0x1d
    "00111100", --  633 - 0x279  :   60 - 0x3c
    "00111010", --  634 - 0x27a  :   58 - 0x3a
    "00111000", --  635 - 0x27b  :   56 - 0x38
    "00110000", --  636 - 0x27c  :   48 - 0x30
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00011100", --  638 - 0x27e  :   28 - 0x1c
    "00111100", --  639 - 0x27f  :   60 - 0x3c
    "00100010", --  640 - 0x280  :   34 - 0x22
    "01010101", --  641 - 0x281  :   85 - 0x55
    "01010101", --  642 - 0x282  :   85 - 0x55
    "01010101", --  643 - 0x283  :   85 - 0x55
    "01010101", --  644 - 0x284  :   85 - 0x55
    "01010101", --  645 - 0x285  :   85 - 0x55
    "01110111", --  646 - 0x286  :  119 - 0x77
    "00100010", --  647 - 0x287  :   34 - 0x22
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0
    "00000000", --  657 - 0x291  :    0 - 0x0
    "11001111", --  658 - 0x292  :  207 - 0xcf
    "00000111", --  659 - 0x293  :    7 - 0x7
    "01111111", --  660 - 0x294  :  127 - 0x7f
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00111100", --  666 - 0x29a  :   60 - 0x3c
    "11111100", --  667 - 0x29b  :  252 - 0xfc
    "11111110", --  668 - 0x29c  :  254 - 0xfe
    "11100000", --  669 - 0x29d  :  224 - 0xe0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "01000000", --  672 - 0x2a0  :   64 - 0x40
    "11100000", --  673 - 0x2a1  :  224 - 0xe0
    "01000000", --  674 - 0x2a2  :   64 - 0x40
    "00111111", --  675 - 0x2a3  :   63 - 0x3f
    "00111110", --  676 - 0x2a4  :   62 - 0x3e
    "00111110", --  677 - 0x2a5  :   62 - 0x3e
    "00110000", --  678 - 0x2a6  :   48 - 0x30
    "00111000", --  679 - 0x2a7  :   56 - 0x38
    "00000000", --  680 - 0x2a8  :    0 - 0x0
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "11111000", --  683 - 0x2ab  :  248 - 0xf8
    "11111000", --  684 - 0x2ac  :  248 - 0xf8
    "11111000", --  685 - 0x2ad  :  248 - 0xf8
    "00011000", --  686 - 0x2ae  :   24 - 0x18
    "00111000", --  687 - 0x2af  :   56 - 0x38
    "00111100", --  688 - 0x2b0  :   60 - 0x3c
    "00111001", --  689 - 0x2b1  :   57 - 0x39
    "00111011", --  690 - 0x2b2  :   59 - 0x3b
    "00111111", --  691 - 0x2b3  :   63 - 0x3f
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "01111000", --  696 - 0x2b8  :  120 - 0x78
    "00111000", --  697 - 0x2b9  :   56 - 0x38
    "10111000", --  698 - 0x2ba  :  184 - 0xb8
    "11111000", --  699 - 0x2bb  :  248 - 0xf8
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00111111", --  704 - 0x2c0  :   63 - 0x3f
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "00001111", --  706 - 0x2c2  :   15 - 0xf
    "01110111", --  707 - 0x2c3  :  119 - 0x77
    "01110111", --  708 - 0x2c4  :  119 - 0x77
    "11110111", --  709 - 0x2c5  :  247 - 0xf7
    "11110111", --  710 - 0x2c6  :  247 - 0xf7
    "11110111", --  711 - 0x2c7  :  247 - 0xf7
    "11111111", --  712 - 0x2c8  :  255 - 0xff
    "11111110", --  713 - 0x2c9  :  254 - 0xfe
    "11111110", --  714 - 0x2ca  :  254 - 0xfe
    "11111110", --  715 - 0x2cb  :  254 - 0xfe
    "11111010", --  716 - 0x2cc  :  250 - 0xfa
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11110011", --  718 - 0x2ce  :  243 - 0xf3
    "11100111", --  719 - 0x2cf  :  231 - 0xe7
    "11110000", --  720 - 0x2d0  :  240 - 0xf0
    "11111000", --  721 - 0x2d1  :  248 - 0xf8
    "11111100", --  722 - 0x2d2  :  252 - 0xfc
    "01111100", --  723 - 0x2d3  :  124 - 0x7c
    "01111000", --  724 - 0x2d4  :  120 - 0x78
    "00111000", --  725 - 0x2d5  :   56 - 0x38
    "00111100", --  726 - 0x2d6  :   60 - 0x3c
    "11111100", --  727 - 0x2d7  :  252 - 0xfc
    "11111111", --  728 - 0x2d8  :  255 - 0xff
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "11000011", --  730 - 0x2da  :  195 - 0xc3
    "10000001", --  731 - 0x2db  :  129 - 0x81
    "10000001", --  732 - 0x2dc  :  129 - 0x81
    "11000011", --  733 - 0x2dd  :  195 - 0xc3
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00001011", --  745 - 0x2e9  :   11 - 0xb
    "00011111", --  746 - 0x2ea  :   31 - 0x1f
    "00011111", --  747 - 0x2eb  :   31 - 0x1f
    "00011110", --  748 - 0x2ec  :   30 - 0x1e
    "00111110", --  749 - 0x2ed  :   62 - 0x3e
    "00001100", --  750 - 0x2ee  :   12 - 0xc
    "00000100", --  751 - 0x2ef  :    4 - 0x4
    "00000000", --  752 - 0x2f0  :    0 - 0x0
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000011", --  760 - 0x2f8  :    3 - 0x3
    "00001111", --  761 - 0x2f9  :   15 - 0xf
    "00001111", --  762 - 0x2fa  :   15 - 0xf
    "00001111", --  763 - 0x2fb  :   15 - 0xf
    "00001111", --  764 - 0x2fc  :   15 - 0xf
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0
    "00011000", --  769 - 0x301  :   24 - 0x18
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "01111110", --  771 - 0x303  :  126 - 0x7e
    "01110110", --  772 - 0x304  :  118 - 0x76
    "11111011", --  773 - 0x305  :  251 - 0xfb
    "11111011", --  774 - 0x306  :  251 - 0xfb
    "11111011", --  775 - 0x307  :  251 - 0xfb
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00010000", --  777 - 0x309  :   16 - 0x10
    "00010000", --  778 - 0x30a  :   16 - 0x10
    "00100000", --  779 - 0x30b  :   32 - 0x20
    "00100000", --  780 - 0x30c  :   32 - 0x20
    "00100000", --  781 - 0x30d  :   32 - 0x20
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "00100000", --  783 - 0x30f  :   32 - 0x20
    "00000000", --  784 - 0x310  :    0 - 0x0
    "00001000", --  785 - 0x311  :    8 - 0x8
    "00001000", --  786 - 0x312  :    8 - 0x8
    "00001000", --  787 - 0x313  :    8 - 0x8
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00001000", --  789 - 0x315  :    8 - 0x8
    "00001000", --  790 - 0x316  :    8 - 0x8
    "00001000", --  791 - 0x317  :    8 - 0x8
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00010000", --  793 - 0x319  :   16 - 0x10
    "00010000", --  794 - 0x31a  :   16 - 0x10
    "00111000", --  795 - 0x31b  :   56 - 0x38
    "00111000", --  796 - 0x31c  :   56 - 0x38
    "00111000", --  797 - 0x31d  :   56 - 0x38
    "00111000", --  798 - 0x31e  :   56 - 0x38
    "00111000", --  799 - 0x31f  :   56 - 0x38
    "00000000", --  800 - 0x320  :    0 - 0x0
    "00011000", --  801 - 0x321  :   24 - 0x18
    "00111100", --  802 - 0x322  :   60 - 0x3c
    "00001110", --  803 - 0x323  :   14 - 0xe
    "00001110", --  804 - 0x324  :   14 - 0xe
    "00000100", --  805 - 0x325  :    4 - 0x4
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000100", --  810 - 0x32a  :    4 - 0x4
    "00000110", --  811 - 0x32b  :    6 - 0x6
    "00011110", --  812 - 0x32c  :   30 - 0x1e
    "00111100", --  813 - 0x32d  :   60 - 0x3c
    "00011000", --  814 - 0x32e  :   24 - 0x18
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000001", --  818 - 0x332  :    1 - 0x1
    "00001010", --  819 - 0x333  :   10 - 0xa
    "00010111", --  820 - 0x334  :   23 - 0x17
    "00001111", --  821 - 0x335  :   15 - 0xf
    "00101111", --  822 - 0x336  :   47 - 0x2f
    "00011111", --  823 - 0x337  :   31 - 0x1f
    "00000000", --  824 - 0x338  :    0 - 0x0
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000101", --  828 - 0x33c  :    5 - 0x5
    "00000111", --  829 - 0x33d  :    7 - 0x7
    "00001111", --  830 - 0x33e  :   15 - 0xf
    "00000111", --  831 - 0x33f  :    7 - 0x7
    "00000000", --  832 - 0x340  :    0 - 0x0
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000001", --  838 - 0x346  :    1 - 0x1
    "00000011", --  839 - 0x347  :    3 - 0x3
    "00000000", --  840 - 0x348  :    0 - 0x0
    "01100000", --  841 - 0x349  :   96 - 0x60
    "11110000", --  842 - 0x34a  :  240 - 0xf0
    "11111000", --  843 - 0x34b  :  248 - 0xf8
    "01111100", --  844 - 0x34c  :  124 - 0x7c
    "00111110", --  845 - 0x34d  :   62 - 0x3e
    "01111110", --  846 - 0x34e  :  126 - 0x7e
    "01111111", --  847 - 0x34f  :  127 - 0x7f
    "00111111", --  848 - 0x350  :   63 - 0x3f
    "01011111", --  849 - 0x351  :   95 - 0x5f
    "01111111", --  850 - 0x352  :  127 - 0x7f
    "00111110", --  851 - 0x353  :   62 - 0x3e
    "00001110", --  852 - 0x354  :   14 - 0xe
    "00001010", --  853 - 0x355  :   10 - 0xa
    "01010001", --  854 - 0x356  :   81 - 0x51
    "00100000", --  855 - 0x357  :   32 - 0x20
    "00000000", --  856 - 0x358  :    0 - 0x0
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00001110", --  862 - 0x35e  :   14 - 0xe
    "00011111", --  863 - 0x35f  :   31 - 0x1f
    "00111111", --  864 - 0x360  :   63 - 0x3f
    "01111111", --  865 - 0x361  :  127 - 0x7f
    "01111111", --  866 - 0x362  :  127 - 0x7f
    "11111110", --  867 - 0x363  :  254 - 0xfe
    "11101100", --  868 - 0x364  :  236 - 0xec
    "11001010", --  869 - 0x365  :  202 - 0xca
    "01010001", --  870 - 0x366  :   81 - 0x51
    "00100000", --  871 - 0x367  :   32 - 0x20
    "00000000", --  872 - 0x368  :    0 - 0x0
    "01000000", --  873 - 0x369  :   64 - 0x40
    "01100011", --  874 - 0x36a  :   99 - 0x63
    "01110111", --  875 - 0x36b  :  119 - 0x77
    "01111100", --  876 - 0x36c  :  124 - 0x7c
    "00111000", --  877 - 0x36d  :   56 - 0x38
    "11111000", --  878 - 0x36e  :  248 - 0xf8
    "11100100", --  879 - 0x36f  :  228 - 0xe4
    "00000000", --  880 - 0x370  :    0 - 0x0
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000011", --  882 - 0x372  :    3 - 0x3
    "00000111", --  883 - 0x373  :    7 - 0x7
    "00001100", --  884 - 0x374  :   12 - 0xc
    "00011000", --  885 - 0x375  :   24 - 0x18
    "11111000", --  886 - 0x376  :  248 - 0xf8
    "11100100", --  887 - 0x377  :  228 - 0xe4
    "00000011", --  888 - 0x378  :    3 - 0x3
    "01000100", --  889 - 0x379  :   68 - 0x44
    "00101000", --  890 - 0x37a  :   40 - 0x28
    "00010000", --  891 - 0x37b  :   16 - 0x10
    "00001000", --  892 - 0x37c  :    8 - 0x8
    "00000100", --  893 - 0x37d  :    4 - 0x4
    "00000011", --  894 - 0x37e  :    3 - 0x3
    "00000100", --  895 - 0x37f  :    4 - 0x4
    "00000011", --  896 - 0x380  :    3 - 0x3
    "00000111", --  897 - 0x381  :    7 - 0x7
    "00001111", --  898 - 0x382  :   15 - 0xf
    "00011111", --  899 - 0x383  :   31 - 0x1f
    "00100111", --  900 - 0x384  :   39 - 0x27
    "01111011", --  901 - 0x385  :  123 - 0x7b
    "01111000", --  902 - 0x386  :  120 - 0x78
    "11111011", --  903 - 0x387  :  251 - 0xfb
    "11000000", --  904 - 0x388  :  192 - 0xc0
    "11100000", --  905 - 0x389  :  224 - 0xe0
    "11110000", --  906 - 0x38a  :  240 - 0xf0
    "11111000", --  907 - 0x38b  :  248 - 0xf8
    "11100100", --  908 - 0x38c  :  228 - 0xe4
    "11011110", --  909 - 0x38d  :  222 - 0xde
    "00011110", --  910 - 0x38e  :   30 - 0x1e
    "11011111", --  911 - 0x38f  :  223 - 0xdf
    "11111111", --  912 - 0x390  :  255 - 0xff
    "11111111", --  913 - 0x391  :  255 - 0xff
    "01111111", --  914 - 0x392  :  127 - 0x7f
    "00001111", --  915 - 0x393  :   15 - 0xf
    "00001111", --  916 - 0x394  :   15 - 0xf
    "00000111", --  917 - 0x395  :    7 - 0x7
    "00000011", --  918 - 0x396  :    3 - 0x3
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111110", --  922 - 0x39a  :  254 - 0xfe
    "11110000", --  923 - 0x39b  :  240 - 0xf0
    "11110000", --  924 - 0x39c  :  240 - 0xf0
    "11000000", --  925 - 0x39d  :  192 - 0xc0
    "10000000", --  926 - 0x39e  :  128 - 0x80
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00011000", --  930 - 0x3a2  :   24 - 0x18
    "00100100", --  931 - 0x3a3  :   36 - 0x24
    "00100100", --  932 - 0x3a4  :   36 - 0x24
    "00011000", --  933 - 0x3a5  :   24 - 0x18
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00111100", --  936 - 0x3a8  :   60 - 0x3c
    "01111110", --  937 - 0x3a9  :  126 - 0x7e
    "11111111", --  938 - 0x3aa  :  255 - 0xff
    "11111111", --  939 - 0x3ab  :  255 - 0xff
    "11111111", --  940 - 0x3ac  :  255 - 0xff
    "11111111", --  941 - 0x3ad  :  255 - 0xff
    "01111110", --  942 - 0x3ae  :  126 - 0x7e
    "00111100", --  943 - 0x3af  :   60 - 0x3c
    "00000011", --  944 - 0x3b0  :    3 - 0x3
    "00000111", --  945 - 0x3b1  :    7 - 0x7
    "00001111", --  946 - 0x3b2  :   15 - 0xf
    "00011111", --  947 - 0x3b3  :   31 - 0x1f
    "00111111", --  948 - 0x3b4  :   63 - 0x3f
    "01100011", --  949 - 0x3b5  :   99 - 0x63
    "01000001", --  950 - 0x3b6  :   65 - 0x41
    "11000001", --  951 - 0x3b7  :  193 - 0xc1
    "11000000", --  952 - 0x3b8  :  192 - 0xc0
    "10000000", --  953 - 0x3b9  :  128 - 0x80
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "10001100", --  956 - 0x3bc  :  140 - 0x8c
    "11111110", --  957 - 0x3bd  :  254 - 0xfe
    "11111110", --  958 - 0x3be  :  254 - 0xfe
    "11110011", --  959 - 0x3bf  :  243 - 0xf3
    "11000001", --  960 - 0x3c0  :  193 - 0xc1
    "11100011", --  961 - 0x3c1  :  227 - 0xe3
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "01000111", --  963 - 0x3c3  :   71 - 0x47
    "00001111", --  964 - 0x3c4  :   15 - 0xf
    "00001111", --  965 - 0x3c5  :   15 - 0xf
    "00001111", --  966 - 0x3c6  :   15 - 0xf
    "00000111", --  967 - 0x3c7  :    7 - 0x7
    "11110001", --  968 - 0x3c8  :  241 - 0xf1
    "11111001", --  969 - 0x3c9  :  249 - 0xf9
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "11100010", --  971 - 0x3cb  :  226 - 0xe2
    "11110000", --  972 - 0x3cc  :  240 - 0xf0
    "11110000", --  973 - 0x3cd  :  240 - 0xf0
    "11110000", --  974 - 0x3ce  :  240 - 0xf0
    "11100000", --  975 - 0x3cf  :  224 - 0xe0
    "00010110", --  976 - 0x3d0  :   22 - 0x16
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000101", --  980 - 0x3d4  :    5 - 0x5
    "00001101", --  981 - 0x3d5  :   13 - 0xd
    "00111111", --  982 - 0x3d6  :   63 - 0x3f
    "00011111", --  983 - 0x3d7  :   31 - 0x1f
    "10000000", --  984 - 0x3d8  :  128 - 0x80
    "10000000", --  985 - 0x3d9  :  128 - 0x80
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "10100000", --  989 - 0x3dd  :  160 - 0xa0
    "10100000", --  990 - 0x3de  :  160 - 0xa0
    "11100000", --  991 - 0x3df  :  224 - 0xe0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000100", --  993 - 0x3e1  :    4 - 0x4
    "01001110", --  994 - 0x3e2  :   78 - 0x4e
    "10001100", --  995 - 0x3e3  :  140 - 0x8c
    "00001100", --  996 - 0x3e4  :   12 - 0xc
    "01111111", --  997 - 0x3e5  :  127 - 0x7f
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000001", -- 1006 - 0x3ee  :    1 - 0x1
    "00000001", -- 1007 - 0x3ef  :    1 - 0x1
    "11111111", -- 1008 - 0x3f0  :  255 - 0xff
    "01111111", -- 1009 - 0x3f1  :  127 - 0x7f
    "00111111", -- 1010 - 0x3f2  :   63 - 0x3f
    "00011111", -- 1011 - 0x3f3  :   31 - 0x1f
    "00001111", -- 1012 - 0x3f4  :   15 - 0xf
    "00000111", -- 1013 - 0x3f5  :    7 - 0x7
    "00000011", -- 1014 - 0x3f6  :    3 - 0x3
    "00000001", -- 1015 - 0x3f7  :    1 - 0x1
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff
    "10000011", -- 1017 - 0x3f9  :  131 - 0x83
    "00101001", -- 1018 - 0x3fa  :   41 - 0x29
    "01101101", -- 1019 - 0x3fb  :  109 - 0x6d
    "01000101", -- 1020 - 0x3fc  :   69 - 0x45
    "00010001", -- 1021 - 0x3fd  :   17 - 0x11
    "00000001", -- 1022 - 0x3fe  :    1 - 0x1
    "11000111", -- 1023 - 0x3ff  :  199 - 0xc7
    "00001000", -- 1024 - 0x400  :    8 - 0x8
    "00001000", -- 1025 - 0x401  :    8 - 0x8
    "00000010", -- 1026 - 0x402  :    2 - 0x2
    "00011111", -- 1027 - 0x403  :   31 - 0x1f
    "00100010", -- 1028 - 0x404  :   34 - 0x22
    "00000010", -- 1029 - 0x405  :    2 - 0x2
    "00000010", -- 1030 - 0x406  :    2 - 0x2
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00001000", -- 1032 - 0x408  :    8 - 0x8
    "00001000", -- 1033 - 0x409  :    8 - 0x8
    "00001000", -- 1034 - 0x40a  :    8 - 0x8
    "00001000", -- 1035 - 0x40b  :    8 - 0x8
    "00001000", -- 1036 - 0x40c  :    8 - 0x8
    "00001000", -- 1037 - 0x40d  :    8 - 0x8
    "00001000", -- 1038 - 0x40e  :    8 - 0x8
    "00001000", -- 1039 - 0x40f  :    8 - 0x8
    "00010000", -- 1040 - 0x410  :   16 - 0x10
    "00011110", -- 1041 - 0x411  :   30 - 0x1e
    "00010000", -- 1042 - 0x412  :   16 - 0x10
    "01010000", -- 1043 - 0x413  :   80 - 0x50
    "00010000", -- 1044 - 0x414  :   16 - 0x10
    "00001000", -- 1045 - 0x415  :    8 - 0x8
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "11111110", -- 1051 - 0x41b  :  254 - 0xfe
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00011100", -- 1056 - 0x420  :   28 - 0x1c
    "00101010", -- 1057 - 0x421  :   42 - 0x2a
    "01110111", -- 1058 - 0x422  :  119 - 0x77
    "11101110", -- 1059 - 0x423  :  238 - 0xee
    "11011101", -- 1060 - 0x424  :  221 - 0xdd
    "10101010", -- 1061 - 0x425  :  170 - 0xaa
    "01110100", -- 1062 - 0x426  :  116 - 0x74
    "00101000", -- 1063 - 0x427  :   40 - 0x28
    "11111111", -- 1064 - 0x428  :  255 - 0xff
    "11111110", -- 1065 - 0x429  :  254 - 0xfe
    "11111110", -- 1066 - 0x42a  :  254 - 0xfe
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "11101111", -- 1068 - 0x42c  :  239 - 0xef
    "11101111", -- 1069 - 0x42d  :  239 - 0xef
    "11101111", -- 1070 - 0x42e  :  239 - 0xef
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "11111110", -- 1072 - 0x430  :  254 - 0xfe
    "11111110", -- 1073 - 0x431  :  254 - 0xfe
    "11111110", -- 1074 - 0x432  :  254 - 0xfe
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "11101111", -- 1076 - 0x434  :  239 - 0xef
    "11101111", -- 1077 - 0x435  :  239 - 0xef
    "11101111", -- 1078 - 0x436  :  239 - 0xef
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "01111111", -- 1081 - 0x439  :  127 - 0x7f
    "01011111", -- 1082 - 0x43a  :   95 - 0x5f
    "01111111", -- 1083 - 0x43b  :  127 - 0x7f
    "01111111", -- 1084 - 0x43c  :  127 - 0x7f
    "01111111", -- 1085 - 0x43d  :  127 - 0x7f
    "01111111", -- 1086 - 0x43e  :  127 - 0x7f
    "01111111", -- 1087 - 0x43f  :  127 - 0x7f
    "10111000", -- 1088 - 0x440  :  184 - 0xb8
    "10011110", -- 1089 - 0x441  :  158 - 0x9e
    "10000000", -- 1090 - 0x442  :  128 - 0x80
    "11000000", -- 1091 - 0x443  :  192 - 0xc0
    "11100000", -- 1092 - 0x444  :  224 - 0xe0
    "11110000", -- 1093 - 0x445  :  240 - 0xf0
    "11111000", -- 1094 - 0x446  :  248 - 0xf8
    "01111100", -- 1095 - 0x447  :  124 - 0x7c
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00100011", -- 1097 - 0x449  :   35 - 0x23
    "01010111", -- 1098 - 0x44a  :   87 - 0x57
    "01001111", -- 1099 - 0x44b  :   79 - 0x4f
    "01010111", -- 1100 - 0x44c  :   87 - 0x57
    "00100111", -- 1101 - 0x44d  :   39 - 0x27
    "11000011", -- 1102 - 0x44e  :  195 - 0xc3
    "00100001", -- 1103 - 0x44f  :   33 - 0x21
    "00000000", -- 1104 - 0x450  :    0 - 0x0
    "00110000", -- 1105 - 0x451  :   48 - 0x30
    "01110000", -- 1106 - 0x452  :  112 - 0x70
    "01110000", -- 1107 - 0x453  :  112 - 0x70
    "11110000", -- 1108 - 0x454  :  240 - 0xf0
    "11100000", -- 1109 - 0x455  :  224 - 0xe0
    "11000000", -- 1110 - 0x456  :  192 - 0xc0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00010011", -- 1112 - 0x458  :   19 - 0x13
    "00001111", -- 1113 - 0x459  :   15 - 0xf
    "00011110", -- 1114 - 0x45a  :   30 - 0x1e
    "11110000", -- 1115 - 0x45b  :  240 - 0xf0
    "11111100", -- 1116 - 0x45c  :  252 - 0xfc
    "11111000", -- 1117 - 0x45d  :  248 - 0xf8
    "11110000", -- 1118 - 0x45e  :  240 - 0xf0
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "10111110", -- 1120 - 0x460  :  190 - 0xbe
    "10010000", -- 1121 - 0x461  :  144 - 0x90
    "10000000", -- 1122 - 0x462  :  128 - 0x80
    "11000000", -- 1123 - 0x463  :  192 - 0xc0
    "11000000", -- 1124 - 0x464  :  192 - 0xc0
    "10000000", -- 1125 - 0x465  :  128 - 0x80
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000001", -- 1128 - 0x468  :    1 - 0x1
    "00000001", -- 1129 - 0x469  :    1 - 0x1
    "00000011", -- 1130 - 0x46a  :    3 - 0x3
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000111", -- 1132 - 0x46c  :    7 - 0x7
    "01111111", -- 1133 - 0x46d  :  127 - 0x7f
    "01111101", -- 1134 - 0x46e  :  125 - 0x7d
    "00111101", -- 1135 - 0x46f  :   61 - 0x3d
    "00000110", -- 1136 - 0x470  :    6 - 0x6
    "00000100", -- 1137 - 0x471  :    4 - 0x4
    "00110000", -- 1138 - 0x472  :   48 - 0x30
    "00100011", -- 1139 - 0x473  :   35 - 0x23
    "00000110", -- 1140 - 0x474  :    6 - 0x6
    "01100100", -- 1141 - 0x475  :  100 - 0x64
    "01100000", -- 1142 - 0x476  :   96 - 0x60
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "01100000", -- 1145 - 0x479  :   96 - 0x60
    "01100000", -- 1146 - 0x47a  :   96 - 0x60
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00100000", -- 1148 - 0x47c  :   32 - 0x20
    "00110000", -- 1149 - 0x47d  :   48 - 0x30
    "00000100", -- 1150 - 0x47e  :    4 - 0x4
    "00000110", -- 1151 - 0x47f  :    6 - 0x6
    "00000000", -- 1152 - 0x480  :    0 - 0x0
    "00000001", -- 1153 - 0x481  :    1 - 0x1
    "00000001", -- 1154 - 0x482  :    1 - 0x1
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "11111110", -- 1160 - 0x488  :  254 - 0xfe
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "01000000", -- 1163 - 0x48b  :   64 - 0x40
    "00000001", -- 1164 - 0x48c  :    1 - 0x1
    "00000011", -- 1165 - 0x48d  :    3 - 0x3
    "00000011", -- 1166 - 0x48e  :    3 - 0x3
    "00000011", -- 1167 - 0x48f  :    3 - 0x3
    "00000001", -- 1168 - 0x490  :    1 - 0x1
    "00000001", -- 1169 - 0x491  :    1 - 0x1
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "11100000", -- 1176 - 0x498  :  224 - 0xe0
    "11111110", -- 1177 - 0x499  :  254 - 0xfe
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "01111111", -- 1179 - 0x49b  :  127 - 0x7f
    "00000011", -- 1180 - 0x49c  :    3 - 0x3
    "00000010", -- 1181 - 0x49d  :    2 - 0x2
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000001", -- 1184 - 0x4a0  :    1 - 0x1
    "00001101", -- 1185 - 0x4a1  :   13 - 0xd
    "00001000", -- 1186 - 0x4a2  :    8 - 0x8
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00110110", -- 1188 - 0x4a4  :   54 - 0x36
    "00101100", -- 1189 - 0x4a5  :   44 - 0x2c
    "00001000", -- 1190 - 0x4a6  :    8 - 0x8
    "01100000", -- 1191 - 0x4a7  :   96 - 0x60
    "01100000", -- 1192 - 0x4a8  :   96 - 0x60
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00100000", -- 1194 - 0x4aa  :   32 - 0x20
    "00110000", -- 1195 - 0x4ab  :   48 - 0x30
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00001000", -- 1197 - 0x4ad  :    8 - 0x8
    "00001101", -- 1198 - 0x4ae  :   13 - 0xd
    "00000001", -- 1199 - 0x4af  :    1 - 0x1
    "00000001", -- 1200 - 0x4b0  :    1 - 0x1
    "00000001", -- 1201 - 0x4b1  :    1 - 0x1
    "00000011", -- 1202 - 0x4b2  :    3 - 0x3
    "01000011", -- 1203 - 0x4b3  :   67 - 0x43
    "01100111", -- 1204 - 0x4b4  :  103 - 0x67
    "01110111", -- 1205 - 0x4b5  :  119 - 0x77
    "01111011", -- 1206 - 0x4b6  :  123 - 0x7b
    "01111000", -- 1207 - 0x4b7  :  120 - 0x78
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "10000000", -- 1210 - 0x4ba  :  128 - 0x80
    "10000100", -- 1211 - 0x4bb  :  132 - 0x84
    "11001100", -- 1212 - 0x4bc  :  204 - 0xcc
    "11011100", -- 1213 - 0x4bd  :  220 - 0xdc
    "10111100", -- 1214 - 0x4be  :  188 - 0xbc
    "00111100", -- 1215 - 0x4bf  :   60 - 0x3c
    "00110011", -- 1216 - 0x4c0  :   51 - 0x33
    "00000111", -- 1217 - 0x4c1  :    7 - 0x7
    "00000111", -- 1218 - 0x4c2  :    7 - 0x7
    "11100011", -- 1219 - 0x4c3  :  227 - 0xe3
    "00111000", -- 1220 - 0x4c4  :   56 - 0x38
    "00111111", -- 1221 - 0x4c5  :   63 - 0x3f
    "00011100", -- 1222 - 0x4c6  :   28 - 0x1c
    "00001100", -- 1223 - 0x4c7  :   12 - 0xc
    "10011000", -- 1224 - 0x4c8  :  152 - 0x98
    "11000111", -- 1225 - 0x4c9  :  199 - 0xc7
    "11001000", -- 1226 - 0x4ca  :  200 - 0xc8
    "10010010", -- 1227 - 0x4cb  :  146 - 0x92
    "00110000", -- 1228 - 0x4cc  :   48 - 0x30
    "11111000", -- 1229 - 0x4cd  :  248 - 0xf8
    "01110000", -- 1230 - 0x4ce  :  112 - 0x70
    "01100000", -- 1231 - 0x4cf  :   96 - 0x60
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0
    "00000001", -- 1233 - 0x4d1  :    1 - 0x1
    "00000001", -- 1234 - 0x4d2  :    1 - 0x1
    "00000011", -- 1235 - 0x4d3  :    3 - 0x3
    "01000011", -- 1236 - 0x4d4  :   67 - 0x43
    "01100111", -- 1237 - 0x4d5  :  103 - 0x67
    "01110111", -- 1238 - 0x4d6  :  119 - 0x77
    "01111011", -- 1239 - 0x4d7  :  123 - 0x7b
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "10000000", -- 1243 - 0x4db  :  128 - 0x80
    "10000100", -- 1244 - 0x4dc  :  132 - 0x84
    "11001100", -- 1245 - 0x4dd  :  204 - 0xcc
    "11011100", -- 1246 - 0x4de  :  220 - 0xdc
    "10111100", -- 1247 - 0x4df  :  188 - 0xbc
    "01111000", -- 1248 - 0x4e0  :  120 - 0x78
    "00110011", -- 1249 - 0x4e1  :   51 - 0x33
    "00000111", -- 1250 - 0x4e2  :    7 - 0x7
    "00000111", -- 1251 - 0x4e3  :    7 - 0x7
    "11100011", -- 1252 - 0x4e4  :  227 - 0xe3
    "00111000", -- 1253 - 0x4e5  :   56 - 0x38
    "01111111", -- 1254 - 0x4e6  :  127 - 0x7f
    "11110000", -- 1255 - 0x4e7  :  240 - 0xf0
    "00111100", -- 1256 - 0x4e8  :   60 - 0x3c
    "10011000", -- 1257 - 0x4e9  :  152 - 0x98
    "11000111", -- 1258 - 0x4ea  :  199 - 0xc7
    "11001000", -- 1259 - 0x4eb  :  200 - 0xc8
    "10010010", -- 1260 - 0x4ec  :  146 - 0x92
    "00110000", -- 1261 - 0x4ed  :   48 - 0x30
    "11111000", -- 1262 - 0x4ee  :  248 - 0xf8
    "00111100", -- 1263 - 0x4ef  :   60 - 0x3c
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0
    "00010000", -- 1265 - 0x4f1  :   16 - 0x10
    "01111111", -- 1266 - 0x4f2  :  127 - 0x7f
    "01111111", -- 1267 - 0x4f3  :  127 - 0x7f
    "01111111", -- 1268 - 0x4f4  :  127 - 0x7f
    "00011111", -- 1269 - 0x4f5  :   31 - 0x1f
    "00001111", -- 1270 - 0x4f6  :   15 - 0xf
    "00001111", -- 1271 - 0x4f7  :   15 - 0xf
    "00000011", -- 1272 - 0x4f8  :    3 - 0x3
    "00110011", -- 1273 - 0x4f9  :   51 - 0x33
    "00111001", -- 1274 - 0x4fa  :   57 - 0x39
    "00111010", -- 1275 - 0x4fb  :   58 - 0x3a
    "00111000", -- 1276 - 0x4fc  :   56 - 0x38
    "00011000", -- 1277 - 0x4fd  :   24 - 0x18
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00010000", -- 1280 - 0x500  :   16 - 0x10
    "00111000", -- 1281 - 0x501  :   56 - 0x38
    "00111100", -- 1282 - 0x502  :   60 - 0x3c
    "01110100", -- 1283 - 0x503  :  116 - 0x74
    "01110110", -- 1284 - 0x504  :  118 - 0x76
    "01110110", -- 1285 - 0x505  :  118 - 0x76
    "01111110", -- 1286 - 0x506  :  126 - 0x7e
    "01111101", -- 1287 - 0x507  :  125 - 0x7d
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00010001", -- 1290 - 0x50a  :   17 - 0x11
    "00001010", -- 1291 - 0x50b  :   10 - 0xa
    "00110100", -- 1292 - 0x50c  :   52 - 0x34
    "00101010", -- 1293 - 0x50d  :   42 - 0x2a
    "01010001", -- 1294 - 0x50e  :   81 - 0x51
    "00100000", -- 1295 - 0x50f  :   32 - 0x20
    "01111111", -- 1296 - 0x510  :  127 - 0x7f
    "01100111", -- 1297 - 0x511  :  103 - 0x67
    "01100011", -- 1298 - 0x512  :   99 - 0x63
    "01110000", -- 1299 - 0x513  :  112 - 0x70
    "00111000", -- 1300 - 0x514  :   56 - 0x38
    "00111110", -- 1301 - 0x515  :   62 - 0x3e
    "01111100", -- 1302 - 0x516  :  124 - 0x7c
    "10111000", -- 1303 - 0x517  :  184 - 0xb8
    "01010001", -- 1304 - 0x518  :   81 - 0x51
    "00001010", -- 1305 - 0x519  :   10 - 0xa
    "00000100", -- 1306 - 0x51a  :    4 - 0x4
    "11101010", -- 1307 - 0x51b  :  234 - 0xea
    "01111001", -- 1308 - 0x51c  :  121 - 0x79
    "01111111", -- 1309 - 0x51d  :  127 - 0x7f
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "00111001", -- 1311 - 0x51f  :   57 - 0x39
    "01011000", -- 1312 - 0x520  :   88 - 0x58
    "00111000", -- 1313 - 0x521  :   56 - 0x38
    "00010000", -- 1314 - 0x522  :   16 - 0x10
    "00110000", -- 1315 - 0x523  :   48 - 0x30
    "11110000", -- 1316 - 0x524  :  240 - 0xf0
    "11110000", -- 1317 - 0x525  :  240 - 0xf0
    "11100000", -- 1318 - 0x526  :  224 - 0xe0
    "11000000", -- 1319 - 0x527  :  192 - 0xc0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00001000", -- 1321 - 0x529  :    8 - 0x8
    "00011100", -- 1322 - 0x52a  :   28 - 0x1c
    "00111100", -- 1323 - 0x52b  :   60 - 0x3c
    "01111010", -- 1324 - 0x52c  :  122 - 0x7a
    "01111010", -- 1325 - 0x52d  :  122 - 0x7a
    "01111010", -- 1326 - 0x52e  :  122 - 0x7a
    "01111110", -- 1327 - 0x52f  :  126 - 0x7e
    "00000000", -- 1328 - 0x530  :    0 - 0x0
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00010001", -- 1331 - 0x533  :   17 - 0x11
    "00001010", -- 1332 - 0x534  :   10 - 0xa
    "00110100", -- 1333 - 0x535  :   52 - 0x34
    "00101010", -- 1334 - 0x536  :   42 - 0x2a
    "01010001", -- 1335 - 0x537  :   81 - 0x51
    "01111111", -- 1336 - 0x538  :  127 - 0x7f
    "01111101", -- 1337 - 0x539  :  125 - 0x7d
    "00111111", -- 1338 - 0x53a  :   63 - 0x3f
    "00110111", -- 1339 - 0x53b  :   55 - 0x37
    "00110011", -- 1340 - 0x53c  :   51 - 0x33
    "00111011", -- 1341 - 0x53d  :   59 - 0x3b
    "00111010", -- 1342 - 0x53e  :   58 - 0x3a
    "01111000", -- 1343 - 0x53f  :  120 - 0x78
    "00100000", -- 1344 - 0x540  :   32 - 0x20
    "01010001", -- 1345 - 0x541  :   81 - 0x51
    "00001010", -- 1346 - 0x542  :   10 - 0xa
    "00000100", -- 1347 - 0x543  :    4 - 0x4
    "11101010", -- 1348 - 0x544  :  234 - 0xea
    "00111001", -- 1349 - 0x545  :   57 - 0x39
    "01111111", -- 1350 - 0x546  :  127 - 0x7f
    "11110000", -- 1351 - 0x547  :  240 - 0xf0
    "10111100", -- 1352 - 0x548  :  188 - 0xbc
    "01011000", -- 1353 - 0x549  :   88 - 0x58
    "00111000", -- 1354 - 0x54a  :   56 - 0x38
    "00010000", -- 1355 - 0x54b  :   16 - 0x10
    "00110000", -- 1356 - 0x54c  :   48 - 0x30
    "11111000", -- 1357 - 0x54d  :  248 - 0xf8
    "11111100", -- 1358 - 0x54e  :  252 - 0xfc
    "00111110", -- 1359 - 0x54f  :   62 - 0x3e
    "00000000", -- 1360 - 0x550  :    0 - 0x0
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000110", -- 1363 - 0x553  :    6 - 0x6
    "00001110", -- 1364 - 0x554  :   14 - 0xe
    "00001100", -- 1365 - 0x555  :   12 - 0xc
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00001111", -- 1374 - 0x55e  :   15 - 0xf
    "00011000", -- 1375 - 0x55f  :   24 - 0x18
    "00000000", -- 1376 - 0x560  :    0 - 0x0
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "11111000", -- 1380 - 0x564  :  248 - 0xf8
    "00111110", -- 1381 - 0x565  :   62 - 0x3e
    "00111011", -- 1382 - 0x566  :   59 - 0x3b
    "00011000", -- 1383 - 0x567  :   24 - 0x18
    "00010000", -- 1384 - 0x568  :   16 - 0x10
    "00010100", -- 1385 - 0x569  :   20 - 0x14
    "00010000", -- 1386 - 0x56a  :   16 - 0x10
    "00010000", -- 1387 - 0x56b  :   16 - 0x10
    "00111000", -- 1388 - 0x56c  :   56 - 0x38
    "01111000", -- 1389 - 0x56d  :  120 - 0x78
    "11111000", -- 1390 - 0x56e  :  248 - 0xf8
    "00110000", -- 1391 - 0x56f  :   48 - 0x30
    "00000000", -- 1392 - 0x570  :    0 - 0x0
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000110", -- 1396 - 0x574  :    6 - 0x6
    "00001110", -- 1397 - 0x575  :   14 - 0xe
    "00001100", -- 1398 - 0x576  :   12 - 0xc
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00001111", -- 1407 - 0x57f  :   15 - 0xf
    "00000000", -- 1408 - 0x580  :    0 - 0x0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "11111000", -- 1413 - 0x585  :  248 - 0xf8
    "01111110", -- 1414 - 0x586  :  126 - 0x7e
    "11110011", -- 1415 - 0x587  :  243 - 0xf3
    "00011000", -- 1416 - 0x588  :   24 - 0x18
    "00010000", -- 1417 - 0x589  :   16 - 0x10
    "00010100", -- 1418 - 0x58a  :   20 - 0x14
    "00010000", -- 1419 - 0x58b  :   16 - 0x10
    "00010000", -- 1420 - 0x58c  :   16 - 0x10
    "00111000", -- 1421 - 0x58d  :   56 - 0x38
    "01111100", -- 1422 - 0x58e  :  124 - 0x7c
    "11011110", -- 1423 - 0x58f  :  222 - 0xde
    "00000000", -- 1424 - 0x590  :    0 - 0x0
    "00001101", -- 1425 - 0x591  :   13 - 0xd
    "00011110", -- 1426 - 0x592  :   30 - 0x1e
    "00011110", -- 1427 - 0x593  :   30 - 0x1e
    "00011110", -- 1428 - 0x594  :   30 - 0x1e
    "00011111", -- 1429 - 0x595  :   31 - 0x1f
    "00001111", -- 1430 - 0x596  :   15 - 0xf
    "00000111", -- 1431 - 0x597  :    7 - 0x7
    "01111000", -- 1432 - 0x598  :  120 - 0x78
    "11110000", -- 1433 - 0x599  :  240 - 0xf0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00011010", -- 1435 - 0x59b  :   26 - 0x1a
    "00111111", -- 1436 - 0x59c  :   63 - 0x3f
    "00110101", -- 1437 - 0x59d  :   53 - 0x35
    "00110101", -- 1438 - 0x59e  :   53 - 0x35
    "00111111", -- 1439 - 0x59f  :   63 - 0x3f
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "10000000", -- 1442 - 0x5a2  :  128 - 0x80
    "11100000", -- 1443 - 0x5a3  :  224 - 0xe0
    "11100000", -- 1444 - 0x5a4  :  224 - 0xe0
    "01110000", -- 1445 - 0x5a5  :  112 - 0x70
    "01110011", -- 1446 - 0x5a6  :  115 - 0x73
    "00100001", -- 1447 - 0x5a7  :   33 - 0x21
    "00011010", -- 1448 - 0x5a8  :   26 - 0x1a
    "00000111", -- 1449 - 0x5a9  :    7 - 0x7
    "00001100", -- 1450 - 0x5aa  :   12 - 0xc
    "00011000", -- 1451 - 0x5ab  :   24 - 0x18
    "01111000", -- 1452 - 0x5ac  :  120 - 0x78
    "11111110", -- 1453 - 0x5ad  :  254 - 0xfe
    "11111100", -- 1454 - 0x5ae  :  252 - 0xfc
    "11110000", -- 1455 - 0x5af  :  240 - 0xf0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0
    "00000001", -- 1457 - 0x5b1  :    1 - 0x1
    "00000010", -- 1458 - 0x5b2  :    2 - 0x2
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00111000", -- 1460 - 0x5b4  :   56 - 0x38
    "01111100", -- 1461 - 0x5b5  :  124 - 0x7c
    "01111110", -- 1462 - 0x5b6  :  126 - 0x7e
    "00111111", -- 1463 - 0x5b7  :   63 - 0x3f
    "00111111", -- 1464 - 0x5b8  :   63 - 0x3f
    "01000000", -- 1465 - 0x5b9  :   64 - 0x40
    "01100000", -- 1466 - 0x5ba  :   96 - 0x60
    "01100000", -- 1467 - 0x5bb  :   96 - 0x60
    "00100000", -- 1468 - 0x5bc  :   32 - 0x20
    "00110000", -- 1469 - 0x5bd  :   48 - 0x30
    "00010011", -- 1470 - 0x5be  :   19 - 0x13
    "00000001", -- 1471 - 0x5bf  :    1 - 0x1
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0
    "11100000", -- 1473 - 0x5c1  :  224 - 0xe0
    "00110000", -- 1474 - 0x5c2  :   48 - 0x30
    "11010000", -- 1475 - 0x5c3  :  208 - 0xd0
    "11010000", -- 1476 - 0x5c4  :  208 - 0xd0
    "11010000", -- 1477 - 0x5c5  :  208 - 0xd0
    "11010000", -- 1478 - 0x5c6  :  208 - 0xd0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000111", -- 1480 - 0x5c8  :    7 - 0x7
    "00001111", -- 1481 - 0x5c9  :   15 - 0xf
    "00000010", -- 1482 - 0x5ca  :    2 - 0x2
    "00011101", -- 1483 - 0x5cb  :   29 - 0x1d
    "00011111", -- 1484 - 0x5cc  :   31 - 0x1f
    "00011010", -- 1485 - 0x5cd  :   26 - 0x1a
    "00011010", -- 1486 - 0x5ce  :   26 - 0x1a
    "00000010", -- 1487 - 0x5cf  :    2 - 0x2
    "00111000", -- 1488 - 0x5d0  :   56 - 0x38
    "01111100", -- 1489 - 0x5d1  :  124 - 0x7c
    "11111100", -- 1490 - 0x5d2  :  252 - 0xfc
    "11111100", -- 1491 - 0x5d3  :  252 - 0xfc
    "11111100", -- 1492 - 0x5d4  :  252 - 0xfc
    "11111110", -- 1493 - 0x5d5  :  254 - 0xfe
    "10111110", -- 1494 - 0x5d6  :  190 - 0xbe
    "10111110", -- 1495 - 0x5d7  :  190 - 0xbe
    "00011100", -- 1496 - 0x5d8  :   28 - 0x1c
    "00111110", -- 1497 - 0x5d9  :   62 - 0x3e
    "00111111", -- 1498 - 0x5da  :   63 - 0x3f
    "00111111", -- 1499 - 0x5db  :   63 - 0x3f
    "00111111", -- 1500 - 0x5dc  :   63 - 0x3f
    "01111111", -- 1501 - 0x5dd  :  127 - 0x7f
    "01111101", -- 1502 - 0x5de  :  125 - 0x7d
    "01111101", -- 1503 - 0x5df  :  125 - 0x7d
    "01111101", -- 1504 - 0x5e0  :  125 - 0x7d
    "01111111", -- 1505 - 0x5e1  :  127 - 0x7f
    "01011111", -- 1506 - 0x5e2  :   95 - 0x5f
    "00111011", -- 1507 - 0x5e3  :   59 - 0x3b
    "00111100", -- 1508 - 0x5e4  :   60 - 0x3c
    "00111111", -- 1509 - 0x5e5  :   63 - 0x3f
    "00011110", -- 1510 - 0x5e6  :   30 - 0x1e
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00011100", -- 1512 - 0x5e8  :   28 - 0x1c
    "00111110", -- 1513 - 0x5e9  :   62 - 0x3e
    "00111111", -- 1514 - 0x5ea  :   63 - 0x3f
    "00011111", -- 1515 - 0x5eb  :   31 - 0x1f
    "00111111", -- 1516 - 0x5ec  :   63 - 0x3f
    "01111111", -- 1517 - 0x5ed  :  127 - 0x7f
    "01111101", -- 1518 - 0x5ee  :  125 - 0x7d
    "01111101", -- 1519 - 0x5ef  :  125 - 0x7d
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "01100000", -- 1523 - 0x5f3  :   96 - 0x60
    "01100010", -- 1524 - 0x5f4  :   98 - 0x62
    "01100101", -- 1525 - 0x5f5  :  101 - 0x65
    "00111111", -- 1526 - 0x5f6  :   63 - 0x3f
    "00011111", -- 1527 - 0x5f7  :   31 - 0x1f
    "01110000", -- 1528 - 0x5f8  :  112 - 0x70
    "00111100", -- 1529 - 0x5f9  :   60 - 0x3c
    "00111100", -- 1530 - 0x5fa  :   60 - 0x3c
    "00011000", -- 1531 - 0x5fb  :   24 - 0x18
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000010", -- 1534 - 0x5fe  :    2 - 0x2
    "00000111", -- 1535 - 0x5ff  :    7 - 0x7
    "11001111", -- 1536 - 0x600  :  207 - 0xcf
    "01111010", -- 1537 - 0x601  :  122 - 0x7a
    "01011010", -- 1538 - 0x602  :   90 - 0x5a
    "00010000", -- 1539 - 0x603  :   16 - 0x10
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "11000000", -- 1542 - 0x606  :  192 - 0xc0
    "10000000", -- 1543 - 0x607  :  128 - 0x80
    "10000101", -- 1544 - 0x608  :  133 - 0x85
    "10000100", -- 1545 - 0x609  :  132 - 0x84
    "10000110", -- 1546 - 0x60a  :  134 - 0x86
    "11000110", -- 1547 - 0x60b  :  198 - 0xc6
    "11100111", -- 1548 - 0x60c  :  231 - 0xe7
    "01110011", -- 1549 - 0x60d  :  115 - 0x73
    "01110011", -- 1550 - 0x60e  :  115 - 0x73
    "11100001", -- 1551 - 0x60f  :  225 - 0xe1
    "10000000", -- 1552 - 0x610  :  128 - 0x80
    "01001110", -- 1553 - 0x611  :   78 - 0x4e
    "01110111", -- 1554 - 0x612  :  119 - 0x77
    "11110011", -- 1555 - 0x613  :  243 - 0xf3
    "11111011", -- 1556 - 0x614  :  251 - 0xfb
    "11111001", -- 1557 - 0x615  :  249 - 0xf9
    "11111010", -- 1558 - 0x616  :  250 - 0xfa
    "01111000", -- 1559 - 0x617  :  120 - 0x78
    "00010001", -- 1560 - 0x618  :   17 - 0x11
    "00111001", -- 1561 - 0x619  :   57 - 0x39
    "01111101", -- 1562 - 0x61a  :  125 - 0x7d
    "00111001", -- 1563 - 0x61b  :   57 - 0x39
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "11100000", -- 1566 - 0x61e  :  224 - 0xe0
    "11100111", -- 1567 - 0x61f  :  231 - 0xe7
    "00000000", -- 1568 - 0x620  :    0 - 0x0
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000111", -- 1570 - 0x622  :    7 - 0x7
    "00000111", -- 1571 - 0x623  :    7 - 0x7
    "00010110", -- 1572 - 0x624  :   22 - 0x16
    "00010000", -- 1573 - 0x625  :   16 - 0x10
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00111000", -- 1575 - 0x627  :   56 - 0x38
    "11001111", -- 1576 - 0x628  :  207 - 0xcf
    "00011111", -- 1577 - 0x629  :   31 - 0x1f
    "00010111", -- 1578 - 0x62a  :   23 - 0x17
    "00010000", -- 1579 - 0x62b  :   16 - 0x10
    "00110011", -- 1580 - 0x62c  :   51 - 0x33
    "00110000", -- 1581 - 0x62d  :   48 - 0x30
    "00110000", -- 1582 - 0x62e  :   48 - 0x30
    "00100000", -- 1583 - 0x62f  :   32 - 0x20
    "00111000", -- 1584 - 0x630  :   56 - 0x38
    "00110000", -- 1585 - 0x631  :   48 - 0x30
    "01000000", -- 1586 - 0x632  :   64 - 0x40
    "11000111", -- 1587 - 0x633  :  199 - 0xc7
    "00000111", -- 1588 - 0x634  :    7 - 0x7
    "01100110", -- 1589 - 0x635  :  102 - 0x66
    "11100000", -- 1590 - 0x636  :  224 - 0xe0
    "01101100", -- 1591 - 0x637  :  108 - 0x6c
    "01100000", -- 1592 - 0x638  :   96 - 0x60
    "11000000", -- 1593 - 0x639  :  192 - 0xc0
    "10000000", -- 1594 - 0x63a  :  128 - 0x80
    "00000100", -- 1595 - 0x63b  :    4 - 0x4
    "10011110", -- 1596 - 0x63c  :  158 - 0x9e
    "11111111", -- 1597 - 0x63d  :  255 - 0xff
    "11110000", -- 1598 - 0x63e  :  240 - 0xf0
    "11111000", -- 1599 - 0x63f  :  248 - 0xf8
    "00100100", -- 1600 - 0x640  :   36 - 0x24
    "00000001", -- 1601 - 0x641  :    1 - 0x1
    "00000111", -- 1602 - 0x642  :    7 - 0x7
    "11111110", -- 1603 - 0x643  :  254 - 0xfe
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "01111111", -- 1605 - 0x645  :  127 - 0x7f
    "00111111", -- 1606 - 0x646  :   63 - 0x3f
    "01111111", -- 1607 - 0x647  :  127 - 0x7f
    "11001111", -- 1608 - 0x648  :  207 - 0xcf
    "01111010", -- 1609 - 0x649  :  122 - 0x7a
    "00001010", -- 1610 - 0x64a  :   10 - 0xa
    "11111110", -- 1611 - 0x64b  :  254 - 0xfe
    "11111100", -- 1612 - 0x64c  :  252 - 0xfc
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "10000101", -- 1616 - 0x650  :  133 - 0x85
    "10000110", -- 1617 - 0x651  :  134 - 0x86
    "10000011", -- 1618 - 0x652  :  131 - 0x83
    "11000011", -- 1619 - 0x653  :  195 - 0xc3
    "11100001", -- 1620 - 0x654  :  225 - 0xe1
    "01110000", -- 1621 - 0x655  :  112 - 0x70
    "01110000", -- 1622 - 0x656  :  112 - 0x70
    "11100000", -- 1623 - 0x657  :  224 - 0xe0
    "01100000", -- 1624 - 0x658  :   96 - 0x60
    "11000000", -- 1625 - 0x659  :  192 - 0xc0
    "10000000", -- 1626 - 0x65a  :  128 - 0x80
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "10011000", -- 1628 - 0x65c  :  152 - 0x98
    "11111100", -- 1629 - 0x65d  :  252 - 0xfc
    "11111110", -- 1630 - 0x65e  :  254 - 0xfe
    "11111111", -- 1631 - 0x65f  :  255 - 0xff
    "00100100", -- 1632 - 0x660  :   36 - 0x24
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000111", -- 1634 - 0x662  :    7 - 0x7
    "11111110", -- 1635 - 0x663  :  254 - 0xfe
    "11111111", -- 1636 - 0x664  :  255 - 0xff
    "01111111", -- 1637 - 0x665  :  127 - 0x7f
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "00000011", -- 1639 - 0x667  :    3 - 0x3
    "00000011", -- 1640 - 0x668  :    3 - 0x3
    "00001111", -- 1641 - 0x669  :   15 - 0xf
    "00100011", -- 1642 - 0x66a  :   35 - 0x23
    "01100010", -- 1643 - 0x66b  :   98 - 0x62
    "01100100", -- 1644 - 0x66c  :  100 - 0x64
    "00111100", -- 1645 - 0x66d  :   60 - 0x3c
    "00011100", -- 1646 - 0x66e  :   28 - 0x1c
    "00011110", -- 1647 - 0x66f  :   30 - 0x1e
    "00011111", -- 1648 - 0x670  :   31 - 0x1f
    "00111101", -- 1649 - 0x671  :   61 - 0x3d
    "01101101", -- 1650 - 0x672  :  109 - 0x6d
    "01001111", -- 1651 - 0x673  :   79 - 0x4f
    "11101110", -- 1652 - 0x674  :  238 - 0xee
    "11110011", -- 1653 - 0x675  :  243 - 0xf3
    "00100000", -- 1654 - 0x676  :   32 - 0x20
    "00000011", -- 1655 - 0x677  :    3 - 0x3
    "00000111", -- 1656 - 0x678  :    7 - 0x7
    "00000111", -- 1657 - 0x679  :    7 - 0x7
    "00011111", -- 1658 - 0x67a  :   31 - 0x1f
    "00111111", -- 1659 - 0x67b  :   63 - 0x3f
    "00001111", -- 1660 - 0x67c  :   15 - 0xf
    "01000111", -- 1661 - 0x67d  :   71 - 0x47
    "00000011", -- 1662 - 0x67e  :    3 - 0x3
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000011", -- 1666 - 0x682  :    3 - 0x3
    "00000111", -- 1667 - 0x683  :    7 - 0x7
    "00001111", -- 1668 - 0x684  :   15 - 0xf
    "00001111", -- 1669 - 0x685  :   15 - 0xf
    "00011111", -- 1670 - 0x686  :   31 - 0x1f
    "00011111", -- 1671 - 0x687  :   31 - 0x1f
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00100011", -- 1673 - 0x689  :   35 - 0x23
    "01010111", -- 1674 - 0x68a  :   87 - 0x57
    "01001111", -- 1675 - 0x68b  :   79 - 0x4f
    "01010111", -- 1676 - 0x68c  :   87 - 0x57
    "00101111", -- 1677 - 0x68d  :   47 - 0x2f
    "11011111", -- 1678 - 0x68e  :  223 - 0xdf
    "00100001", -- 1679 - 0x68f  :   33 - 0x21
    "00000000", -- 1680 - 0x690  :    0 - 0x0
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "10000000", -- 1684 - 0x694  :  128 - 0x80
    "10000000", -- 1685 - 0x695  :  128 - 0x80
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00100011", -- 1688 - 0x698  :   35 - 0x23
    "00001111", -- 1689 - 0x699  :   15 - 0xf
    "00011110", -- 1690 - 0x69a  :   30 - 0x1e
    "11110000", -- 1691 - 0x69b  :  240 - 0xf0
    "00011100", -- 1692 - 0x69c  :   28 - 0x1c
    "00111111", -- 1693 - 0x69d  :   63 - 0x3f
    "00011111", -- 1694 - 0x69e  :   31 - 0x1f
    "00011110", -- 1695 - 0x69f  :   30 - 0x1e
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0
    "10000000", -- 1697 - 0x6a1  :  128 - 0x80
    "00011000", -- 1698 - 0x6a2  :   24 - 0x18
    "00110000", -- 1699 - 0x6a3  :   48 - 0x30
    "00110100", -- 1700 - 0x6a4  :   52 - 0x34
    "11111110", -- 1701 - 0x6a5  :  254 - 0xfe
    "11111110", -- 1702 - 0x6a6  :  254 - 0xfe
    "11111110", -- 1703 - 0x6a7  :  254 - 0xfe
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000001", -- 1706 - 0x6aa  :    1 - 0x1
    "00000100", -- 1707 - 0x6ab  :    4 - 0x4
    "00000110", -- 1708 - 0x6ac  :    6 - 0x6
    "00000110", -- 1709 - 0x6ad  :    6 - 0x6
    "00000111", -- 1710 - 0x6ae  :    7 - 0x7
    "00000111", -- 1711 - 0x6af  :    7 - 0x7
    "00001111", -- 1712 - 0x6b0  :   15 - 0xf
    "00111111", -- 1713 - 0x6b1  :   63 - 0x3f
    "01111111", -- 1714 - 0x6b2  :  127 - 0x7f
    "11111000", -- 1715 - 0x6b3  :  248 - 0xf8
    "11111000", -- 1716 - 0x6b4  :  248 - 0xf8
    "01111111", -- 1717 - 0x6b5  :  127 - 0x7f
    "00111111", -- 1718 - 0x6b6  :   63 - 0x3f
    "00001111", -- 1719 - 0x6b7  :   15 - 0xf
    "00011111", -- 1720 - 0x6b8  :   31 - 0x1f
    "00011111", -- 1721 - 0x6b9  :   31 - 0x1f
    "00011111", -- 1722 - 0x6ba  :   31 - 0x1f
    "00001011", -- 1723 - 0x6bb  :   11 - 0xb
    "00000001", -- 1724 - 0x6bc  :    1 - 0x1
    "00000001", -- 1725 - 0x6bd  :    1 - 0x1
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000011", -- 1728 - 0x6c0  :    3 - 0x3
    "00011111", -- 1729 - 0x6c1  :   31 - 0x1f
    "00111111", -- 1730 - 0x6c2  :   63 - 0x3f
    "00111111", -- 1731 - 0x6c3  :   63 - 0x3f
    "01111000", -- 1732 - 0x6c4  :  120 - 0x78
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000011", -- 1734 - 0x6c6  :    3 - 0x3
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00100011", -- 1744 - 0x6d0  :   35 - 0x23
    "00100111", -- 1745 - 0x6d1  :   39 - 0x27
    "00011111", -- 1746 - 0x6d2  :   31 - 0x1f
    "00000111", -- 1747 - 0x6d3  :    7 - 0x7
    "00001111", -- 1748 - 0x6d4  :   15 - 0xf
    "00011111", -- 1749 - 0x6d5  :   31 - 0x1f
    "01111111", -- 1750 - 0x6d6  :  127 - 0x7f
    "00111111", -- 1751 - 0x6d7  :   63 - 0x3f
    "11100000", -- 1752 - 0x6d8  :  224 - 0xe0
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "10000000", -- 1754 - 0x6da  :  128 - 0x80
    "01000000", -- 1755 - 0x6db  :   64 - 0x40
    "11100000", -- 1756 - 0x6dc  :  224 - 0xe0
    "11100000", -- 1757 - 0x6dd  :  224 - 0xe0
    "11100000", -- 1758 - 0x6de  :  224 - 0xe0
    "11000000", -- 1759 - 0x6df  :  192 - 0xc0
    "00000011", -- 1760 - 0x6e0  :    3 - 0x3
    "00000111", -- 1761 - 0x6e1  :    7 - 0x7
    "00001111", -- 1762 - 0x6e2  :   15 - 0xf
    "00011111", -- 1763 - 0x6e3  :   31 - 0x1f
    "00111111", -- 1764 - 0x6e4  :   63 - 0x3f
    "01111111", -- 1765 - 0x6e5  :  127 - 0x7f
    "11111111", -- 1766 - 0x6e6  :  255 - 0xff
    "00011111", -- 1767 - 0x6e7  :   31 - 0x1f
    "00011111", -- 1768 - 0x6e8  :   31 - 0x1f
    "00010000", -- 1769 - 0x6e9  :   16 - 0x10
    "00001100", -- 1770 - 0x6ea  :   12 - 0xc
    "00010010", -- 1771 - 0x6eb  :   18 - 0x12
    "00010010", -- 1772 - 0x6ec  :   18 - 0x12
    "00101100", -- 1773 - 0x6ed  :   44 - 0x2c
    "00111111", -- 1774 - 0x6ee  :   63 - 0x3f
    "00111111", -- 1775 - 0x6ef  :   63 - 0x3f
    "00110111", -- 1776 - 0x6f0  :   55 - 0x37
    "00110110", -- 1777 - 0x6f1  :   54 - 0x36
    "00110110", -- 1778 - 0x6f2  :   54 - 0x36
    "00110110", -- 1779 - 0x6f3  :   54 - 0x36
    "00010110", -- 1780 - 0x6f4  :   22 - 0x16
    "00010110", -- 1781 - 0x6f5  :   22 - 0x16
    "00010010", -- 1782 - 0x6f6  :   18 - 0x12
    "00000010", -- 1783 - 0x6f7  :    2 - 0x2
    "00010000", -- 1784 - 0x6f8  :   16 - 0x10
    "01111110", -- 1785 - 0x6f9  :  126 - 0x7e
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11110110", -- 1788 - 0x6fc  :  246 - 0xf6
    "01110110", -- 1789 - 0x6fd  :  118 - 0x76
    "00111010", -- 1790 - 0x6fe  :   58 - 0x3a
    "00011010", -- 1791 - 0x6ff  :   26 - 0x1a
    "00000000", -- 1792 - 0x700  :    0 - 0x0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00111000", -- 1794 - 0x702  :   56 - 0x38
    "00000100", -- 1795 - 0x703  :    4 - 0x4
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00111000", -- 1803 - 0x70b  :   56 - 0x38
    "01000000", -- 1804 - 0x70c  :   64 - 0x40
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "11111100", -- 1808 - 0x710  :  252 - 0xfc
    "10100000", -- 1809 - 0x711  :  160 - 0xa0
    "10000000", -- 1810 - 0x712  :  128 - 0x80
    "10000000", -- 1811 - 0x713  :  128 - 0x80
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000111", -- 1816 - 0x718  :    7 - 0x7
    "00100111", -- 1817 - 0x719  :   39 - 0x27
    "01010111", -- 1818 - 0x71a  :   87 - 0x57
    "01001111", -- 1819 - 0x71b  :   79 - 0x4f
    "01010111", -- 1820 - 0x71c  :   87 - 0x57
    "00100111", -- 1821 - 0x71d  :   39 - 0x27
    "11000001", -- 1822 - 0x71e  :  193 - 0xc1
    "00100001", -- 1823 - 0x71f  :   33 - 0x21
    "00011101", -- 1824 - 0x720  :   29 - 0x1d
    "00001111", -- 1825 - 0x721  :   15 - 0xf
    "00001111", -- 1826 - 0x722  :   15 - 0xf
    "00011111", -- 1827 - 0x723  :   31 - 0x1f
    "00011111", -- 1828 - 0x724  :   31 - 0x1f
    "00011110", -- 1829 - 0x725  :   30 - 0x1e
    "00111000", -- 1830 - 0x726  :   56 - 0x38
    "00110000", -- 1831 - 0x727  :   48 - 0x30
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00111000", -- 1834 - 0x72a  :   56 - 0x38
    "00010000", -- 1835 - 0x72b  :   16 - 0x10
    "01001100", -- 1836 - 0x72c  :   76 - 0x4c
    "00011000", -- 1837 - 0x72d  :   24 - 0x18
    "10000110", -- 1838 - 0x72e  :  134 - 0x86
    "00100100", -- 1839 - 0x72f  :   36 - 0x24
    "00000000", -- 1840 - 0x730  :    0 - 0x0
    "01000010", -- 1841 - 0x731  :   66 - 0x42
    "00001010", -- 1842 - 0x732  :   10 - 0xa
    "01000000", -- 1843 - 0x733  :   64 - 0x40
    "00010000", -- 1844 - 0x734  :   16 - 0x10
    "00000010", -- 1845 - 0x735  :    2 - 0x2
    "00001000", -- 1846 - 0x736  :    8 - 0x8
    "00000010", -- 1847 - 0x737  :    2 - 0x2
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "10000000", -- 1850 - 0x73a  :  128 - 0x80
    "01000000", -- 1851 - 0x73b  :   64 - 0x40
    "00001000", -- 1852 - 0x73c  :    8 - 0x8
    "00001100", -- 1853 - 0x73d  :   12 - 0xc
    "00001010", -- 1854 - 0x73e  :   10 - 0xa
    "10000100", -- 1855 - 0x73f  :  132 - 0x84
    "00000000", -- 1856 - 0x740  :    0 - 0x0
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "11001111", -- 1858 - 0x742  :  207 - 0xcf
    "00100000", -- 1859 - 0x743  :   32 - 0x20
    "00100000", -- 1860 - 0x744  :   32 - 0x20
    "00100000", -- 1861 - 0x745  :   32 - 0x20
    "00100110", -- 1862 - 0x746  :   38 - 0x26
    "00101110", -- 1863 - 0x747  :   46 - 0x2e
    "11100000", -- 1864 - 0x748  :  224 - 0xe0
    "11100000", -- 1865 - 0x749  :  224 - 0xe0
    "11000000", -- 1866 - 0x74a  :  192 - 0xc0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00101111", -- 1872 - 0x750  :   47 - 0x2f
    "00100011", -- 1873 - 0x751  :   35 - 0x23
    "00100001", -- 1874 - 0x752  :   33 - 0x21
    "00100000", -- 1875 - 0x753  :   32 - 0x20
    "00100000", -- 1876 - 0x754  :   32 - 0x20
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "11000001", -- 1880 - 0x758  :  193 - 0xc1
    "10110001", -- 1881 - 0x759  :  177 - 0xb1
    "01011001", -- 1882 - 0x75a  :   89 - 0x59
    "01101101", -- 1883 - 0x75b  :  109 - 0x6d
    "00110101", -- 1884 - 0x75c  :   53 - 0x35
    "00111011", -- 1885 - 0x75d  :   59 - 0x3b
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000011", -- 1887 - 0x75f  :    3 - 0x3
    "00000000", -- 1888 - 0x760  :    0 - 0x0
    "00000010", -- 1889 - 0x761  :    2 - 0x2
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00001000", -- 1891 - 0x763  :    8 - 0x8
    "00000010", -- 1892 - 0x764  :    2 - 0x2
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00101000", -- 1894 - 0x766  :   40 - 0x28
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000100", -- 1896 - 0x768  :    4 - 0x4
    "00010000", -- 1897 - 0x769  :   16 - 0x10
    "00000010", -- 1898 - 0x76a  :    2 - 0x2
    "00010000", -- 1899 - 0x76b  :   16 - 0x10
    "00000100", -- 1900 - 0x76c  :    4 - 0x4
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00001010", -- 1902 - 0x76e  :   10 - 0xa
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "11000001", -- 1904 - 0x770  :  193 - 0xc1
    "10110001", -- 1905 - 0x771  :  177 - 0xb1
    "01011001", -- 1906 - 0x772  :   89 - 0x59
    "01101101", -- 1907 - 0x773  :  109 - 0x6d
    "00110101", -- 1908 - 0x774  :   53 - 0x35
    "00111011", -- 1909 - 0x775  :   59 - 0x3b
    "00011111", -- 1910 - 0x776  :   31 - 0x1f
    "00000011", -- 1911 - 0x777  :    3 - 0x3
    "00000000", -- 1912 - 0x778  :    0 - 0x0
    "00001111", -- 1913 - 0x779  :   15 - 0xf
    "00011111", -- 1914 - 0x77a  :   31 - 0x1f
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111100", -- 1916 - 0x77c  :  252 - 0xfc
    "01100011", -- 1917 - 0x77d  :   99 - 0x63
    "00011111", -- 1918 - 0x77e  :   31 - 0x1f
    "00000011", -- 1919 - 0x77f  :    3 - 0x3
    "00000000", -- 1920 - 0x780  :    0 - 0x0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "11111110", -- 1922 - 0x782  :  254 - 0xfe
    "11000110", -- 1923 - 0x783  :  198 - 0xc6
    "11000110", -- 1924 - 0x784  :  198 - 0xc6
    "11111110", -- 1925 - 0x785  :  254 - 0xfe
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000110", -- 1930 - 0x78a  :    6 - 0x6
    "00000110", -- 1931 - 0x78b  :    6 - 0x6
    "00001100", -- 1932 - 0x78c  :   12 - 0xc
    "00011000", -- 1933 - 0x78d  :   24 - 0x18
    "01110000", -- 1934 - 0x78e  :  112 - 0x70
    "01100000", -- 1935 - 0x78f  :   96 - 0x60
    "00000000", -- 1936 - 0x790  :    0 - 0x0
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000110", -- 1938 - 0x792  :    6 - 0x6
    "00000110", -- 1939 - 0x793  :    6 - 0x6
    "00000100", -- 1940 - 0x794  :    4 - 0x4
    "00000100", -- 1941 - 0x795  :    4 - 0x4
    "00001000", -- 1942 - 0x796  :    8 - 0x8
    "00001000", -- 1943 - 0x797  :    8 - 0x8
    "00001000", -- 1944 - 0x798  :    8 - 0x8
    "00010000", -- 1945 - 0x799  :   16 - 0x10
    "00110000", -- 1946 - 0x79a  :   48 - 0x30
    "00110000", -- 1947 - 0x79b  :   48 - 0x30
    "00110000", -- 1948 - 0x79c  :   48 - 0x30
    "00110000", -- 1949 - 0x79d  :   48 - 0x30
    "00010000", -- 1950 - 0x79e  :   16 - 0x10
    "00001000", -- 1951 - 0x79f  :    8 - 0x8
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000001", -- 1954 - 0x7a2  :    1 - 0x1
    "00000011", -- 1955 - 0x7a3  :    3 - 0x3
    "00000001", -- 1956 - 0x7a4  :    1 - 0x1
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000011", -- 1960 - 0x7a8  :    3 - 0x3
    "00001110", -- 1961 - 0x7a9  :   14 - 0xe
    "11111000", -- 1962 - 0x7aa  :  248 - 0xf8
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00100010", -- 1968 - 0x7b0  :   34 - 0x22
    "01100101", -- 1969 - 0x7b1  :  101 - 0x65
    "00100101", -- 1970 - 0x7b2  :   37 - 0x25
    "00100101", -- 1971 - 0x7b3  :   37 - 0x25
    "00100101", -- 1972 - 0x7b4  :   37 - 0x25
    "00100101", -- 1973 - 0x7b5  :   37 - 0x25
    "01110111", -- 1974 - 0x7b6  :  119 - 0x77
    "01110010", -- 1975 - 0x7b7  :  114 - 0x72
    "01100010", -- 1976 - 0x7b8  :   98 - 0x62
    "10010101", -- 1977 - 0x7b9  :  149 - 0x95
    "00010101", -- 1978 - 0x7ba  :   21 - 0x15
    "00100101", -- 1979 - 0x7bb  :   37 - 0x25
    "01000101", -- 1980 - 0x7bc  :   69 - 0x45
    "10000101", -- 1981 - 0x7bd  :  133 - 0x85
    "11110111", -- 1982 - 0x7be  :  247 - 0xf7
    "11110010", -- 1983 - 0x7bf  :  242 - 0xf2
    "10100010", -- 1984 - 0x7c0  :  162 - 0xa2
    "10100101", -- 1985 - 0x7c1  :  165 - 0xa5
    "10100101", -- 1986 - 0x7c2  :  165 - 0xa5
    "10100101", -- 1987 - 0x7c3  :  165 - 0xa5
    "11110101", -- 1988 - 0x7c4  :  245 - 0xf5
    "11110101", -- 1989 - 0x7c5  :  245 - 0xf5
    "00100111", -- 1990 - 0x7c6  :   39 - 0x27
    "00100010", -- 1991 - 0x7c7  :   34 - 0x22
    "11110010", -- 1992 - 0x7c8  :  242 - 0xf2
    "10000101", -- 1993 - 0x7c9  :  133 - 0x85
    "10000101", -- 1994 - 0x7ca  :  133 - 0x85
    "11100101", -- 1995 - 0x7cb  :  229 - 0xe5
    "00010101", -- 1996 - 0x7cc  :   21 - 0x15
    "00010101", -- 1997 - 0x7cd  :   21 - 0x15
    "11110111", -- 1998 - 0x7ce  :  247 - 0xf7
    "11100010", -- 1999 - 0x7cf  :  226 - 0xe2
    "01100010", -- 2000 - 0x7d0  :   98 - 0x62
    "10010101", -- 2001 - 0x7d1  :  149 - 0x95
    "01010101", -- 2002 - 0x7d2  :   85 - 0x55
    "01100101", -- 2003 - 0x7d3  :  101 - 0x65
    "10110101", -- 2004 - 0x7d4  :  181 - 0xb5
    "10010101", -- 2005 - 0x7d5  :  149 - 0x95
    "10010111", -- 2006 - 0x7d6  :  151 - 0x97
    "01100010", -- 2007 - 0x7d7  :   98 - 0x62
    "00100000", -- 2008 - 0x7d8  :   32 - 0x20
    "01010000", -- 2009 - 0x7d9  :   80 - 0x50
    "01010000", -- 2010 - 0x7da  :   80 - 0x50
    "01010000", -- 2011 - 0x7db  :   80 - 0x50
    "01010000", -- 2012 - 0x7dc  :   80 - 0x50
    "01010000", -- 2013 - 0x7dd  :   80 - 0x50
    "01110000", -- 2014 - 0x7de  :  112 - 0x70
    "00100000", -- 2015 - 0x7df  :   32 - 0x20
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "01100110", -- 2024 - 0x7e8  :  102 - 0x66
    "11100110", -- 2025 - 0x7e9  :  230 - 0xe6
    "01100110", -- 2026 - 0x7ea  :  102 - 0x66
    "01100110", -- 2027 - 0x7eb  :  102 - 0x66
    "01100110", -- 2028 - 0x7ec  :  102 - 0x66
    "01100111", -- 2029 - 0x7ed  :  103 - 0x67
    "11110011", -- 2030 - 0x7ee  :  243 - 0xf3
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "01011110", -- 2032 - 0x7f0  :   94 - 0x5e
    "01011001", -- 2033 - 0x7f1  :   89 - 0x59
    "01011001", -- 2034 - 0x7f2  :   89 - 0x59
    "01011001", -- 2035 - 0x7f3  :   89 - 0x59
    "01011110", -- 2036 - 0x7f4  :   94 - 0x5e
    "11011000", -- 2037 - 0x7f5  :  216 - 0xd8
    "10011000", -- 2038 - 0x7f6  :  152 - 0x98
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000100", -- 2045 - 0x7fd  :    4 - 0x4
    "00001000", -- 2046 - 0x7fe  :    8 - 0x8
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "00000000", -- 2048 - 0x800  :    0 - 0x0
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000000", -- 2050 - 0x802  :    0 - 0x0
    "00000000", -- 2051 - 0x803  :    0 - 0x0
    "00000000", -- 2052 - 0x804  :    0 - 0x0
    "00000000", -- 2053 - 0x805  :    0 - 0x0
    "00000000", -- 2054 - 0x806  :    0 - 0x0
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00000000", -- 2056 - 0x808  :    0 - 0x0
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000000", -- 2059 - 0x80b  :    0 - 0x0
    "00000000", -- 2060 - 0x80c  :    0 - 0x0
    "00000000", -- 2061 - 0x80d  :    0 - 0x0
    "00000000", -- 2062 - 0x80e  :    0 - 0x0
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "00000000", -- 2064 - 0x810  :    0 - 0x0
    "00000000", -- 2065 - 0x811  :    0 - 0x0
    "00000000", -- 2066 - 0x812  :    0 - 0x0
    "00000000", -- 2067 - 0x813  :    0 - 0x0
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00000000", -- 2072 - 0x818  :    0 - 0x0
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00000000", -- 2075 - 0x81b  :    0 - 0x0
    "00000000", -- 2076 - 0x81c  :    0 - 0x0
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00000000", -- 2080 - 0x820  :    0 - 0x0
    "00000000", -- 2081 - 0x821  :    0 - 0x0
    "00000000", -- 2082 - 0x822  :    0 - 0x0
    "00000000", -- 2083 - 0x823  :    0 - 0x0
    "00000000", -- 2084 - 0x824  :    0 - 0x0
    "00000000", -- 2085 - 0x825  :    0 - 0x0
    "00000000", -- 2086 - 0x826  :    0 - 0x0
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "00000000", -- 2088 - 0x828  :    0 - 0x0
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "00000000", -- 2092 - 0x82c  :    0 - 0x0
    "00000000", -- 2093 - 0x82d  :    0 - 0x0
    "00000000", -- 2094 - 0x82e  :    0 - 0x0
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00000000", -- 2096 - 0x830  :    0 - 0x0
    "00000000", -- 2097 - 0x831  :    0 - 0x0
    "00000000", -- 2098 - 0x832  :    0 - 0x0
    "00000000", -- 2099 - 0x833  :    0 - 0x0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "00000000", -- 2104 - 0x838  :    0 - 0x0
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0
    "00000000", -- 2113 - 0x841  :    0 - 0x0
    "00000000", -- 2114 - 0x842  :    0 - 0x0
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000000", -- 2116 - 0x844  :    0 - 0x0
    "00000000", -- 2117 - 0x845  :    0 - 0x0
    "00000000", -- 2118 - 0x846  :    0 - 0x0
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "00000000", -- 2120 - 0x848  :    0 - 0x0
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "00000000", -- 2124 - 0x84c  :    0 - 0x0
    "00000000", -- 2125 - 0x84d  :    0 - 0x0
    "00000000", -- 2126 - 0x84e  :    0 - 0x0
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00000000", -- 2128 - 0x850  :    0 - 0x0
    "00000000", -- 2129 - 0x851  :    0 - 0x0
    "00000000", -- 2130 - 0x852  :    0 - 0x0
    "00000000", -- 2131 - 0x853  :    0 - 0x0
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00000000", -- 2136 - 0x858  :    0 - 0x0
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "00000000", -- 2148 - 0x864  :    0 - 0x0
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00000000", -- 2150 - 0x866  :    0 - 0x0
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "00000000", -- 2152 - 0x868  :    0 - 0x0
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "00000000", -- 2157 - 0x86d  :    0 - 0x0
    "00000000", -- 2158 - 0x86e  :    0 - 0x0
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0
    "00000000", -- 2161 - 0x871  :    0 - 0x0
    "00000000", -- 2162 - 0x872  :    0 - 0x0
    "00000000", -- 2163 - 0x873  :    0 - 0x0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "00000000", -- 2168 - 0x878  :    0 - 0x0
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0
    "00000000", -- 2177 - 0x881  :    0 - 0x0
    "00000000", -- 2178 - 0x882  :    0 - 0x0
    "00000000", -- 2179 - 0x883  :    0 - 0x0
    "00000000", -- 2180 - 0x884  :    0 - 0x0
    "00000000", -- 2181 - 0x885  :    0 - 0x0
    "00000000", -- 2182 - 0x886  :    0 - 0x0
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "00000000", -- 2184 - 0x888  :    0 - 0x0
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "00000000", -- 2190 - 0x88e  :    0 - 0x0
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "00000000", -- 2192 - 0x890  :    0 - 0x0
    "00000000", -- 2193 - 0x891  :    0 - 0x0
    "00000000", -- 2194 - 0x892  :    0 - 0x0
    "00000000", -- 2195 - 0x893  :    0 - 0x0
    "00000000", -- 2196 - 0x894  :    0 - 0x0
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000000", -- 2200 - 0x898  :    0 - 0x0
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000000", -- 2203 - 0x89b  :    0 - 0x0
    "00000000", -- 2204 - 0x89c  :    0 - 0x0
    "00000000", -- 2205 - 0x89d  :    0 - 0x0
    "00000000", -- 2206 - 0x89e  :    0 - 0x0
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "00000000", -- 2212 - 0x8a4  :    0 - 0x0
    "00000000", -- 2213 - 0x8a5  :    0 - 0x0
    "00000000", -- 2214 - 0x8a6  :    0 - 0x0
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00000000", -- 2222 - 0x8ae  :    0 - 0x0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "00000000", -- 2224 - 0x8b0  :    0 - 0x0
    "00000000", -- 2225 - 0x8b1  :    0 - 0x0
    "00000000", -- 2226 - 0x8b2  :    0 - 0x0
    "00000000", -- 2227 - 0x8b3  :    0 - 0x0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "00000000", -- 2230 - 0x8b6  :    0 - 0x0
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00000000", -- 2232 - 0x8b8  :    0 - 0x0
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00000000", -- 2234 - 0x8ba  :    0 - 0x0
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00000000", -- 2236 - 0x8bc  :    0 - 0x0
    "00000000", -- 2237 - 0x8bd  :    0 - 0x0
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000000", -- 2244 - 0x8c4  :    0 - 0x0
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "00000000", -- 2246 - 0x8c6  :    0 - 0x0
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "00000000", -- 2256 - 0x8d0  :    0 - 0x0
    "00000000", -- 2257 - 0x8d1  :    0 - 0x0
    "00000000", -- 2258 - 0x8d2  :    0 - 0x0
    "00000000", -- 2259 - 0x8d3  :    0 - 0x0
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "00000000", -- 2267 - 0x8db  :    0 - 0x0
    "00000000", -- 2268 - 0x8dc  :    0 - 0x0
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000000", -- 2270 - 0x8de  :    0 - 0x0
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "00000000", -- 2276 - 0x8e4  :    0 - 0x0
    "00000000", -- 2277 - 0x8e5  :    0 - 0x0
    "00000000", -- 2278 - 0x8e6  :    0 - 0x0
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "00000000", -- 2283 - 0x8eb  :    0 - 0x0
    "00000000", -- 2284 - 0x8ec  :    0 - 0x0
    "00000000", -- 2285 - 0x8ed  :    0 - 0x0
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "00000000", -- 2288 - 0x8f0  :    0 - 0x0
    "00000000", -- 2289 - 0x8f1  :    0 - 0x0
    "00000000", -- 2290 - 0x8f2  :    0 - 0x0
    "00000000", -- 2291 - 0x8f3  :    0 - 0x0
    "00000000", -- 2292 - 0x8f4  :    0 - 0x0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00000000", -- 2298 - 0x8fa  :    0 - 0x0
    "00000000", -- 2299 - 0x8fb  :    0 - 0x0
    "00000000", -- 2300 - 0x8fc  :    0 - 0x0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000000", -- 2308 - 0x904  :    0 - 0x0
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "00000000", -- 2310 - 0x906  :    0 - 0x0
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00000000", -- 2316 - 0x90c  :    0 - 0x0
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "00000000", -- 2318 - 0x90e  :    0 - 0x0
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "00000000", -- 2320 - 0x910  :    0 - 0x0
    "00000000", -- 2321 - 0x911  :    0 - 0x0
    "00000000", -- 2322 - 0x912  :    0 - 0x0
    "00000000", -- 2323 - 0x913  :    0 - 0x0
    "00000000", -- 2324 - 0x914  :    0 - 0x0
    "00000000", -- 2325 - 0x915  :    0 - 0x0
    "00000000", -- 2326 - 0x916  :    0 - 0x0
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "00000000", -- 2328 - 0x918  :    0 - 0x0
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00000000", -- 2331 - 0x91b  :    0 - 0x0
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00000000", -- 2344 - 0x928  :    0 - 0x0
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "00000000", -- 2349 - 0x92d  :    0 - 0x0
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "11111111", -- 2352 - 0x930  :  255 - 0xff
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "11111111", -- 2354 - 0x932  :  255 - 0xff
    "11111111", -- 2355 - 0x933  :  255 - 0xff
    "11111111", -- 2356 - 0x934  :  255 - 0xff
    "11111111", -- 2357 - 0x935  :  255 - 0xff
    "11111111", -- 2358 - 0x936  :  255 - 0xff
    "11111111", -- 2359 - 0x937  :  255 - 0xff
    "11111111", -- 2360 - 0x938  :  255 - 0xff
    "11111111", -- 2361 - 0x939  :  255 - 0xff
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "11111111", -- 2363 - 0x93b  :  255 - 0xff
    "11111111", -- 2364 - 0x93c  :  255 - 0xff
    "11111111", -- 2365 - 0x93d  :  255 - 0xff
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "11111111", -- 2367 - 0x93f  :  255 - 0xff
    "00000000", -- 2368 - 0x940  :    0 - 0x0
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00000000", -- 2372 - 0x944  :    0 - 0x0
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00000000", -- 2376 - 0x948  :    0 - 0x0
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00000000", -- 2380 - 0x94c  :    0 - 0x0
    "00000000", -- 2381 - 0x94d  :    0 - 0x0
    "00000000", -- 2382 - 0x94e  :    0 - 0x0
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "01111111", -- 2384 - 0x950  :  127 - 0x7f
    "01111111", -- 2385 - 0x951  :  127 - 0x7f
    "01111111", -- 2386 - 0x952  :  127 - 0x7f
    "01111111", -- 2387 - 0x953  :  127 - 0x7f
    "01111111", -- 2388 - 0x954  :  127 - 0x7f
    "01111111", -- 2389 - 0x955  :  127 - 0x7f
    "01111111", -- 2390 - 0x956  :  127 - 0x7f
    "01111111", -- 2391 - 0x957  :  127 - 0x7f
    "00000000", -- 2392 - 0x958  :    0 - 0x0
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "11111111", -- 2400 - 0x960  :  255 - 0xff
    "10000000", -- 2401 - 0x961  :  128 - 0x80
    "10000000", -- 2402 - 0x962  :  128 - 0x80
    "10000000", -- 2403 - 0x963  :  128 - 0x80
    "10000000", -- 2404 - 0x964  :  128 - 0x80
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00011100", -- 2406 - 0x966  :   28 - 0x1c
    "00111110", -- 2407 - 0x967  :   62 - 0x3e
    "01111111", -- 2408 - 0x968  :  127 - 0x7f
    "01111111", -- 2409 - 0x969  :  127 - 0x7f
    "01111111", -- 2410 - 0x96a  :  127 - 0x7f
    "00111110", -- 2411 - 0x96b  :   62 - 0x3e
    "00011100", -- 2412 - 0x96c  :   28 - 0x1c
    "00000000", -- 2413 - 0x96d  :    0 - 0x0
    "00000000", -- 2414 - 0x96e  :    0 - 0x0
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00001000", -- 2416 - 0x970  :    8 - 0x8
    "00000100", -- 2417 - 0x971  :    4 - 0x4
    "00000100", -- 2418 - 0x972  :    4 - 0x4
    "00000100", -- 2419 - 0x973  :    4 - 0x4
    "00000100", -- 2420 - 0x974  :    4 - 0x4
    "00000100", -- 2421 - 0x975  :    4 - 0x4
    "00001000", -- 2422 - 0x976  :    8 - 0x8
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000011", -- 2424 - 0x978  :    3 - 0x3
    "00000101", -- 2425 - 0x979  :    5 - 0x5
    "00001011", -- 2426 - 0x97a  :   11 - 0xb
    "00001011", -- 2427 - 0x97b  :   11 - 0xb
    "00001111", -- 2428 - 0x97c  :   15 - 0xf
    "00001111", -- 2429 - 0x97d  :   15 - 0xf
    "00000111", -- 2430 - 0x97e  :    7 - 0x7
    "00000011", -- 2431 - 0x97f  :    3 - 0x3
    "00000001", -- 2432 - 0x980  :    1 - 0x1
    "00000011", -- 2433 - 0x981  :    3 - 0x3
    "00000111", -- 2434 - 0x982  :    7 - 0x7
    "00001111", -- 2435 - 0x983  :   15 - 0xf
    "00011111", -- 2436 - 0x984  :   31 - 0x1f
    "00111111", -- 2437 - 0x985  :   63 - 0x3f
    "01111111", -- 2438 - 0x986  :  127 - 0x7f
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "00000000", -- 2440 - 0x988  :    0 - 0x0
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000111", -- 2445 - 0x98d  :    7 - 0x7
    "00111111", -- 2446 - 0x98e  :   63 - 0x3f
    "11111111", -- 2447 - 0x98f  :  255 - 0xff
    "00000000", -- 2448 - 0x990  :    0 - 0x0
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "11100000", -- 2453 - 0x995  :  224 - 0xe0
    "11111100", -- 2454 - 0x996  :  252 - 0xfc
    "11111111", -- 2455 - 0x997  :  255 - 0xff
    "10000000", -- 2456 - 0x998  :  128 - 0x80
    "11000000", -- 2457 - 0x999  :  192 - 0xc0
    "11100000", -- 2458 - 0x99a  :  224 - 0xe0
    "11110000", -- 2459 - 0x99b  :  240 - 0xf0
    "11111000", -- 2460 - 0x99c  :  248 - 0xf8
    "11111100", -- 2461 - 0x99d  :  252 - 0xfc
    "11111110", -- 2462 - 0x99e  :  254 - 0xfe
    "11111111", -- 2463 - 0x99f  :  255 - 0xff
    "11111111", -- 2464 - 0x9a0  :  255 - 0xff
    "11111111", -- 2465 - 0x9a1  :  255 - 0xff
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "11111111", -- 2467 - 0x9a3  :  255 - 0xff
    "11111111", -- 2468 - 0x9a4  :  255 - 0xff
    "11111111", -- 2469 - 0x9a5  :  255 - 0xff
    "11111111", -- 2470 - 0x9a6  :  255 - 0xff
    "11111111", -- 2471 - 0x9a7  :  255 - 0xff
    "00000111", -- 2472 - 0x9a8  :    7 - 0x7
    "00001000", -- 2473 - 0x9a9  :    8 - 0x8
    "00010000", -- 2474 - 0x9aa  :   16 - 0x10
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "01100000", -- 2476 - 0x9ac  :   96 - 0x60
    "10000000", -- 2477 - 0x9ad  :  128 - 0x80
    "10000000", -- 2478 - 0x9ae  :  128 - 0x80
    "01000000", -- 2479 - 0x9af  :   64 - 0x40
    "00000011", -- 2480 - 0x9b0  :    3 - 0x3
    "00000100", -- 2481 - 0x9b1  :    4 - 0x4
    "00011000", -- 2482 - 0x9b2  :   24 - 0x18
    "00100000", -- 2483 - 0x9b3  :   32 - 0x20
    "00100000", -- 2484 - 0x9b4  :   32 - 0x20
    "00100000", -- 2485 - 0x9b5  :   32 - 0x20
    "01000110", -- 2486 - 0x9b6  :   70 - 0x46
    "10001000", -- 2487 - 0x9b7  :  136 - 0x88
    "11000000", -- 2488 - 0x9b8  :  192 - 0xc0
    "00100000", -- 2489 - 0x9b9  :   32 - 0x20
    "00010000", -- 2490 - 0x9ba  :   16 - 0x10
    "00010100", -- 2491 - 0x9bb  :   20 - 0x14
    "00001010", -- 2492 - 0x9bc  :   10 - 0xa
    "01000001", -- 2493 - 0x9bd  :   65 - 0x41
    "00100001", -- 2494 - 0x9be  :   33 - 0x21
    "00000001", -- 2495 - 0x9bf  :    1 - 0x1
    "10010000", -- 2496 - 0x9c0  :  144 - 0x90
    "10101000", -- 2497 - 0x9c1  :  168 - 0xa8
    "01001000", -- 2498 - 0x9c2  :   72 - 0x48
    "00001010", -- 2499 - 0x9c3  :   10 - 0xa
    "00000101", -- 2500 - 0x9c4  :    5 - 0x5
    "00000001", -- 2501 - 0x9c5  :    1 - 0x1
    "00000001", -- 2502 - 0x9c6  :    1 - 0x1
    "00000010", -- 2503 - 0x9c7  :    2 - 0x2
    "00100100", -- 2504 - 0x9c8  :   36 - 0x24
    "00010010", -- 2505 - 0x9c9  :   18 - 0x12
    "00001001", -- 2506 - 0x9ca  :    9 - 0x9
    "00001000", -- 2507 - 0x9cb  :    8 - 0x8
    "00000111", -- 2508 - 0x9cc  :    7 - 0x7
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0
    "01000000", -- 2513 - 0x9d1  :   64 - 0x40
    "11100011", -- 2514 - 0x9d2  :  227 - 0xe3
    "00111111", -- 2515 - 0x9d3  :   63 - 0x3f
    "00001100", -- 2516 - 0x9d4  :   12 - 0xc
    "10000001", -- 2517 - 0x9d5  :  129 - 0x81
    "01100010", -- 2518 - 0x9d6  :   98 - 0x62
    "00011100", -- 2519 - 0x9d7  :   28 - 0x1c
    "01000000", -- 2520 - 0x9d8  :   64 - 0x40
    "10000000", -- 2521 - 0x9d9  :  128 - 0x80
    "11000010", -- 2522 - 0x9da  :  194 - 0xc2
    "01111100", -- 2523 - 0x9db  :  124 - 0x7c
    "00111000", -- 2524 - 0x9dc  :   56 - 0x38
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "11000011", -- 2526 - 0x9de  :  195 - 0xc3
    "00111100", -- 2527 - 0x9df  :   60 - 0x3c
    "00000100", -- 2528 - 0x9e0  :    4 - 0x4
    "00000010", -- 2529 - 0x9e1  :    2 - 0x2
    "00000001", -- 2530 - 0x9e2  :    1 - 0x1
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000110", -- 2532 - 0x9e4  :    6 - 0x6
    "10011000", -- 2533 - 0x9e5  :  152 - 0x98
    "01100000", -- 2534 - 0x9e6  :   96 - 0x60
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "11000000", -- 2536 - 0x9e8  :  192 - 0xc0
    "11100000", -- 2537 - 0x9e9  :  224 - 0xe0
    "11110000", -- 2538 - 0x9ea  :  240 - 0xf0
    "11110000", -- 2539 - 0x9eb  :  240 - 0xf0
    "11110000", -- 2540 - 0x9ec  :  240 - 0xf0
    "11110000", -- 2541 - 0x9ed  :  240 - 0xf0
    "11100000", -- 2542 - 0x9ee  :  224 - 0xe0
    "11000000", -- 2543 - 0x9ef  :  192 - 0xc0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00011100", -- 2550 - 0x9f6  :   28 - 0x1c
    "00111110", -- 2551 - 0x9f7  :   62 - 0x3e
    "01111111", -- 2552 - 0x9f8  :  127 - 0x7f
    "01111111", -- 2553 - 0x9f9  :  127 - 0x7f
    "01111111", -- 2554 - 0x9fa  :  127 - 0x7f
    "00111110", -- 2555 - 0x9fb  :   62 - 0x3e
    "00011100", -- 2556 - 0x9fc  :   28 - 0x1c
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "11111111", -- 2560 - 0xa00  :  255 - 0xff
    "11111111", -- 2561 - 0xa01  :  255 - 0xff
    "11111111", -- 2562 - 0xa02  :  255 - 0xff
    "11111111", -- 2563 - 0xa03  :  255 - 0xff
    "11111111", -- 2564 - 0xa04  :  255 - 0xff
    "11111111", -- 2565 - 0xa05  :  255 - 0xff
    "11111111", -- 2566 - 0xa06  :  255 - 0xff
    "11111111", -- 2567 - 0xa07  :  255 - 0xff
    "00000000", -- 2568 - 0xa08  :    0 - 0x0
    "00001000", -- 2569 - 0xa09  :    8 - 0x8
    "00011000", -- 2570 - 0xa0a  :   24 - 0x18
    "00111000", -- 2571 - 0xa0b  :   56 - 0x38
    "11111100", -- 2572 - 0xa0c  :  252 - 0xfc
    "10111111", -- 2573 - 0xa0d  :  191 - 0xbf
    "01011110", -- 2574 - 0xa0e  :   94 - 0x5e
    "11011001", -- 2575 - 0xa0f  :  217 - 0xd9
    "10000001", -- 2576 - 0xa10  :  129 - 0x81
    "10000001", -- 2577 - 0xa11  :  129 - 0x81
    "10000001", -- 2578 - 0xa12  :  129 - 0x81
    "10000001", -- 2579 - 0xa13  :  129 - 0x81
    "10000001", -- 2580 - 0xa14  :  129 - 0x81
    "10000001", -- 2581 - 0xa15  :  129 - 0x81
    "10000001", -- 2582 - 0xa16  :  129 - 0x81
    "10000001", -- 2583 - 0xa17  :  129 - 0x81
    "00000001", -- 2584 - 0xa18  :    1 - 0x1
    "00000001", -- 2585 - 0xa19  :    1 - 0x1
    "00000001", -- 2586 - 0xa1a  :    1 - 0x1
    "00000001", -- 2587 - 0xa1b  :    1 - 0x1
    "00000001", -- 2588 - 0xa1c  :    1 - 0x1
    "00000001", -- 2589 - 0xa1d  :    1 - 0x1
    "00000001", -- 2590 - 0xa1e  :    1 - 0x1
    "00000001", -- 2591 - 0xa1f  :    1 - 0x1
    "00000000", -- 2592 - 0xa20  :    0 - 0x0
    "01111111", -- 2593 - 0xa21  :  127 - 0x7f
    "01111111", -- 2594 - 0xa22  :  127 - 0x7f
    "01100111", -- 2595 - 0xa23  :  103 - 0x67
    "01100111", -- 2596 - 0xa24  :  103 - 0x67
    "01111111", -- 2597 - 0xa25  :  127 - 0x7f
    "01111111", -- 2598 - 0xa26  :  127 - 0x7f
    "01111111", -- 2599 - 0xa27  :  127 - 0x7f
    "00000000", -- 2600 - 0xa28  :    0 - 0x0
    "11111111", -- 2601 - 0xa29  :  255 - 0xff
    "11111111", -- 2602 - 0xa2a  :  255 - 0xff
    "11111111", -- 2603 - 0xa2b  :  255 - 0xff
    "11111111", -- 2604 - 0xa2c  :  255 - 0xff
    "11111111", -- 2605 - 0xa2d  :  255 - 0xff
    "11111111", -- 2606 - 0xa2e  :  255 - 0xff
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "01111111", -- 2608 - 0xa30  :  127 - 0x7f
    "01111111", -- 2609 - 0xa31  :  127 - 0x7f
    "01111111", -- 2610 - 0xa32  :  127 - 0x7f
    "01111111", -- 2611 - 0xa33  :  127 - 0x7f
    "01111111", -- 2612 - 0xa34  :  127 - 0x7f
    "01111111", -- 2613 - 0xa35  :  127 - 0x7f
    "01111111", -- 2614 - 0xa36  :  127 - 0x7f
    "01111111", -- 2615 - 0xa37  :  127 - 0x7f
    "11111111", -- 2616 - 0xa38  :  255 - 0xff
    "11111111", -- 2617 - 0xa39  :  255 - 0xff
    "11111111", -- 2618 - 0xa3a  :  255 - 0xff
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "00000000", -- 2624 - 0xa40  :    0 - 0x0
    "11111111", -- 2625 - 0xa41  :  255 - 0xff
    "11111111", -- 2626 - 0xa42  :  255 - 0xff
    "11111111", -- 2627 - 0xa43  :  255 - 0xff
    "11111111", -- 2628 - 0xa44  :  255 - 0xff
    "11111111", -- 2629 - 0xa45  :  255 - 0xff
    "11111111", -- 2630 - 0xa46  :  255 - 0xff
    "11111111", -- 2631 - 0xa47  :  255 - 0xff
    "00000000", -- 2632 - 0xa48  :    0 - 0x0
    "11111111", -- 2633 - 0xa49  :  255 - 0xff
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11100111", -- 2635 - 0xa4b  :  231 - 0xe7
    "11100111", -- 2636 - 0xa4c  :  231 - 0xe7
    "11111111", -- 2637 - 0xa4d  :  255 - 0xff
    "11111111", -- 2638 - 0xa4e  :  255 - 0xff
    "11111111", -- 2639 - 0xa4f  :  255 - 0xff
    "11111111", -- 2640 - 0xa50  :  255 - 0xff
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "11111111", -- 2643 - 0xa53  :  255 - 0xff
    "11111111", -- 2644 - 0xa54  :  255 - 0xff
    "11111111", -- 2645 - 0xa55  :  255 - 0xff
    "11111111", -- 2646 - 0xa56  :  255 - 0xff
    "11111111", -- 2647 - 0xa57  :  255 - 0xff
    "00111111", -- 2648 - 0xa58  :   63 - 0x3f
    "01100000", -- 2649 - 0xa59  :   96 - 0x60
    "01000000", -- 2650 - 0xa5a  :   64 - 0x40
    "11000000", -- 2651 - 0xa5b  :  192 - 0xc0
    "10000000", -- 2652 - 0xa5c  :  128 - 0x80
    "10000000", -- 2653 - 0xa5d  :  128 - 0x80
    "10000000", -- 2654 - 0xa5e  :  128 - 0x80
    "10000000", -- 2655 - 0xa5f  :  128 - 0x80
    "10000000", -- 2656 - 0xa60  :  128 - 0x80
    "10000000", -- 2657 - 0xa61  :  128 - 0x80
    "10000000", -- 2658 - 0xa62  :  128 - 0x80
    "10000000", -- 2659 - 0xa63  :  128 - 0x80
    "10000000", -- 2660 - 0xa64  :  128 - 0x80
    "10000001", -- 2661 - 0xa65  :  129 - 0x81
    "01000010", -- 2662 - 0xa66  :   66 - 0x42
    "00111100", -- 2663 - 0xa67  :   60 - 0x3c
    "11111111", -- 2664 - 0xa68  :  255 - 0xff
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0
    "00000000", -- 2673 - 0xa71  :    0 - 0x0
    "00000000", -- 2674 - 0xa72  :    0 - 0x0
    "00000000", -- 2675 - 0xa73  :    0 - 0x0
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "00000001", -- 2677 - 0xa75  :    1 - 0x1
    "10000010", -- 2678 - 0xa76  :  130 - 0x82
    "01111100", -- 2679 - 0xa77  :  124 - 0x7c
    "00000000", -- 2680 - 0xa78  :    0 - 0x0
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000001", -- 2685 - 0xa7d  :    1 - 0x1
    "10000011", -- 2686 - 0xa7e  :  131 - 0x83
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "11111000", -- 2688 - 0xa80  :  248 - 0xf8
    "00000100", -- 2689 - 0xa81  :    4 - 0x4
    "00000010", -- 2690 - 0xa82  :    2 - 0x2
    "00000010", -- 2691 - 0xa83  :    2 - 0x2
    "00000001", -- 2692 - 0xa84  :    1 - 0x1
    "00000001", -- 2693 - 0xa85  :    1 - 0x1
    "00000001", -- 2694 - 0xa86  :    1 - 0x1
    "00000001", -- 2695 - 0xa87  :    1 - 0x1
    "00000001", -- 2696 - 0xa88  :    1 - 0x1
    "00000001", -- 2697 - 0xa89  :    1 - 0x1
    "00000001", -- 2698 - 0xa8a  :    1 - 0x1
    "00000001", -- 2699 - 0xa8b  :    1 - 0x1
    "00000001", -- 2700 - 0xa8c  :    1 - 0x1
    "10000001", -- 2701 - 0xa8d  :  129 - 0x81
    "01000010", -- 2702 - 0xa8e  :   66 - 0x42
    "00111100", -- 2703 - 0xa8f  :   60 - 0x3c
    "11111111", -- 2704 - 0xa90  :  255 - 0xff
    "11111111", -- 2705 - 0xa91  :  255 - 0xff
    "11111111", -- 2706 - 0xa92  :  255 - 0xff
    "11111111", -- 2707 - 0xa93  :  255 - 0xff
    "11111111", -- 2708 - 0xa94  :  255 - 0xff
    "11111111", -- 2709 - 0xa95  :  255 - 0xff
    "11111111", -- 2710 - 0xa96  :  255 - 0xff
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "01111111", -- 2712 - 0xa98  :  127 - 0x7f
    "10000000", -- 2713 - 0xa99  :  128 - 0x80
    "10100000", -- 2714 - 0xa9a  :  160 - 0xa0
    "10000111", -- 2715 - 0xa9b  :  135 - 0x87
    "10001111", -- 2716 - 0xa9c  :  143 - 0x8f
    "10001110", -- 2717 - 0xa9d  :  142 - 0x8e
    "10001110", -- 2718 - 0xa9e  :  142 - 0x8e
    "10000110", -- 2719 - 0xa9f  :  134 - 0x86
    "11111110", -- 2720 - 0xaa0  :  254 - 0xfe
    "00000001", -- 2721 - 0xaa1  :    1 - 0x1
    "00000101", -- 2722 - 0xaa2  :    5 - 0x5
    "11000001", -- 2723 - 0xaa3  :  193 - 0xc1
    "11100001", -- 2724 - 0xaa4  :  225 - 0xe1
    "01110001", -- 2725 - 0xaa5  :  113 - 0x71
    "01110001", -- 2726 - 0xaa6  :  113 - 0x71
    "11110001", -- 2727 - 0xaa7  :  241 - 0xf1
    "10000001", -- 2728 - 0xaa8  :  129 - 0x81
    "10000001", -- 2729 - 0xaa9  :  129 - 0x81
    "10000000", -- 2730 - 0xaaa  :  128 - 0x80
    "10000001", -- 2731 - 0xaab  :  129 - 0x81
    "10000001", -- 2732 - 0xaac  :  129 - 0x81
    "10100000", -- 2733 - 0xaad  :  160 - 0xa0
    "10000000", -- 2734 - 0xaae  :  128 - 0x80
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "11110001", -- 2736 - 0xab0  :  241 - 0xf1
    "11000001", -- 2737 - 0xab1  :  193 - 0xc1
    "11000001", -- 2738 - 0xab2  :  193 - 0xc1
    "10000001", -- 2739 - 0xab3  :  129 - 0x81
    "11000001", -- 2740 - 0xab4  :  193 - 0xc1
    "11000101", -- 2741 - 0xab5  :  197 - 0xc5
    "00000001", -- 2742 - 0xab6  :    1 - 0x1
    "11111111", -- 2743 - 0xab7  :  255 - 0xff
    "01111111", -- 2744 - 0xab8  :  127 - 0x7f
    "11111111", -- 2745 - 0xab9  :  255 - 0xff
    "11111111", -- 2746 - 0xaba  :  255 - 0xff
    "11111111", -- 2747 - 0xabb  :  255 - 0xff
    "11111111", -- 2748 - 0xabc  :  255 - 0xff
    "11111111", -- 2749 - 0xabd  :  255 - 0xff
    "11111111", -- 2750 - 0xabe  :  255 - 0xff
    "11111111", -- 2751 - 0xabf  :  255 - 0xff
    "11111110", -- 2752 - 0xac0  :  254 - 0xfe
    "11111111", -- 2753 - 0xac1  :  255 - 0xff
    "11111111", -- 2754 - 0xac2  :  255 - 0xff
    "11111111", -- 2755 - 0xac3  :  255 - 0xff
    "11111111", -- 2756 - 0xac4  :  255 - 0xff
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "11111111", -- 2758 - 0xac6  :  255 - 0xff
    "11111111", -- 2759 - 0xac7  :  255 - 0xff
    "11111111", -- 2760 - 0xac8  :  255 - 0xff
    "11111111", -- 2761 - 0xac9  :  255 - 0xff
    "11111111", -- 2762 - 0xaca  :  255 - 0xff
    "11111111", -- 2763 - 0xacb  :  255 - 0xff
    "11111111", -- 2764 - 0xacc  :  255 - 0xff
    "11111111", -- 2765 - 0xacd  :  255 - 0xff
    "11111111", -- 2766 - 0xace  :  255 - 0xff
    "01111111", -- 2767 - 0xacf  :  127 - 0x7f
    "11111111", -- 2768 - 0xad0  :  255 - 0xff
    "11111111", -- 2769 - 0xad1  :  255 - 0xff
    "11111111", -- 2770 - 0xad2  :  255 - 0xff
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "11111111", -- 2772 - 0xad4  :  255 - 0xff
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111110", -- 2775 - 0xad7  :  254 - 0xfe
    "00000000", -- 2776 - 0xad8  :    0 - 0x0
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00111000", -- 2782 - 0xade  :   56 - 0x38
    "01111100", -- 2783 - 0xadf  :  124 - 0x7c
    "11111110", -- 2784 - 0xae0  :  254 - 0xfe
    "11111110", -- 2785 - 0xae1  :  254 - 0xfe
    "11111110", -- 2786 - 0xae2  :  254 - 0xfe
    "01111100", -- 2787 - 0xae3  :  124 - 0x7c
    "00111000", -- 2788 - 0xae4  :   56 - 0x38
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00100000", -- 2792 - 0xae8  :   32 - 0x20
    "11100111", -- 2793 - 0xae9  :  231 - 0xe7
    "11100111", -- 2794 - 0xaea  :  231 - 0xe7
    "11100111", -- 2795 - 0xaeb  :  231 - 0xe7
    "11100111", -- 2796 - 0xaec  :  231 - 0xe7
    "11100111", -- 2797 - 0xaed  :  231 - 0xe7
    "11101111", -- 2798 - 0xaee  :  239 - 0xef
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000010", -- 2800 - 0xaf0  :    2 - 0x2
    "01111110", -- 2801 - 0xaf1  :  126 - 0x7e
    "01111110", -- 2802 - 0xaf2  :  126 - 0x7e
    "01111110", -- 2803 - 0xaf3  :  126 - 0x7e
    "01111110", -- 2804 - 0xaf4  :  126 - 0x7e
    "01111110", -- 2805 - 0xaf5  :  126 - 0x7e
    "11111110", -- 2806 - 0xaf6  :  254 - 0xfe
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "01111111", -- 2808 - 0xaf8  :  127 - 0x7f
    "01111111", -- 2809 - 0xaf9  :  127 - 0x7f
    "01111111", -- 2810 - 0xafa  :  127 - 0x7f
    "01100111", -- 2811 - 0xafb  :  103 - 0x67
    "01100111", -- 2812 - 0xafc  :  103 - 0x67
    "01111111", -- 2813 - 0xafd  :  127 - 0x7f
    "01111111", -- 2814 - 0xafe  :  127 - 0x7f
    "01111111", -- 2815 - 0xaff  :  127 - 0x7f
    "11111111", -- 2816 - 0xb00  :  255 - 0xff
    "10000000", -- 2817 - 0xb01  :  128 - 0x80
    "11111100", -- 2818 - 0xb02  :  252 - 0xfc
    "10001100", -- 2819 - 0xb03  :  140 - 0x8c
    "10001100", -- 2820 - 0xb04  :  140 - 0x8c
    "10001100", -- 2821 - 0xb05  :  140 - 0x8c
    "10001100", -- 2822 - 0xb06  :  140 - 0x8c
    "10001100", -- 2823 - 0xb07  :  140 - 0x8c
    "11111111", -- 2824 - 0xb08  :  255 - 0xff
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00001111", -- 2826 - 0xb0a  :   15 - 0xf
    "00001001", -- 2827 - 0xb0b  :    9 - 0x9
    "00001001", -- 2828 - 0xb0c  :    9 - 0x9
    "00001001", -- 2829 - 0xb0d  :    9 - 0x9
    "00001001", -- 2830 - 0xb0e  :    9 - 0x9
    "00001001", -- 2831 - 0xb0f  :    9 - 0x9
    "11111111", -- 2832 - 0xb10  :  255 - 0xff
    "00000000", -- 2833 - 0xb11  :    0 - 0x0
    "11111111", -- 2834 - 0xb12  :  255 - 0xff
    "11111111", -- 2835 - 0xb13  :  255 - 0xff
    "11111111", -- 2836 - 0xb14  :  255 - 0xff
    "11111111", -- 2837 - 0xb15  :  255 - 0xff
    "11111111", -- 2838 - 0xb16  :  255 - 0xff
    "11111111", -- 2839 - 0xb17  :  255 - 0xff
    "11111111", -- 2840 - 0xb18  :  255 - 0xff
    "00000001", -- 2841 - 0xb19  :    1 - 0x1
    "11111111", -- 2842 - 0xb1a  :  255 - 0xff
    "10101001", -- 2843 - 0xb1b  :  169 - 0xa9
    "11010001", -- 2844 - 0xb1c  :  209 - 0xd1
    "10101001", -- 2845 - 0xb1d  :  169 - 0xa9
    "11010001", -- 2846 - 0xb1e  :  209 - 0xd1
    "10101001", -- 2847 - 0xb1f  :  169 - 0xa9
    "10001100", -- 2848 - 0xb20  :  140 - 0x8c
    "10001100", -- 2849 - 0xb21  :  140 - 0x8c
    "10001100", -- 2850 - 0xb22  :  140 - 0x8c
    "10001100", -- 2851 - 0xb23  :  140 - 0x8c
    "10001100", -- 2852 - 0xb24  :  140 - 0x8c
    "10001100", -- 2853 - 0xb25  :  140 - 0x8c
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "00111111", -- 2855 - 0xb27  :   63 - 0x3f
    "00001001", -- 2856 - 0xb28  :    9 - 0x9
    "00001001", -- 2857 - 0xb29  :    9 - 0x9
    "00001001", -- 2858 - 0xb2a  :    9 - 0x9
    "00001001", -- 2859 - 0xb2b  :    9 - 0x9
    "00001001", -- 2860 - 0xb2c  :    9 - 0x9
    "00001001", -- 2861 - 0xb2d  :    9 - 0x9
    "11111111", -- 2862 - 0xb2e  :  255 - 0xff
    "11111111", -- 2863 - 0xb2f  :  255 - 0xff
    "11111111", -- 2864 - 0xb30  :  255 - 0xff
    "11111111", -- 2865 - 0xb31  :  255 - 0xff
    "11111111", -- 2866 - 0xb32  :  255 - 0xff
    "11111111", -- 2867 - 0xb33  :  255 - 0xff
    "11111111", -- 2868 - 0xb34  :  255 - 0xff
    "11111111", -- 2869 - 0xb35  :  255 - 0xff
    "11111111", -- 2870 - 0xb36  :  255 - 0xff
    "11111111", -- 2871 - 0xb37  :  255 - 0xff
    "11010001", -- 2872 - 0xb38  :  209 - 0xd1
    "10101001", -- 2873 - 0xb39  :  169 - 0xa9
    "11010001", -- 2874 - 0xb3a  :  209 - 0xd1
    "10101001", -- 2875 - 0xb3b  :  169 - 0xa9
    "11010001", -- 2876 - 0xb3c  :  209 - 0xd1
    "10101001", -- 2877 - 0xb3d  :  169 - 0xa9
    "11111111", -- 2878 - 0xb3e  :  255 - 0xff
    "11111100", -- 2879 - 0xb3f  :  252 - 0xfc
    "00100011", -- 2880 - 0xb40  :   35 - 0x23
    "00100011", -- 2881 - 0xb41  :   35 - 0x23
    "00100011", -- 2882 - 0xb42  :   35 - 0x23
    "00100011", -- 2883 - 0xb43  :   35 - 0x23
    "00100011", -- 2884 - 0xb44  :   35 - 0x23
    "00100011", -- 2885 - 0xb45  :   35 - 0x23
    "00100011", -- 2886 - 0xb46  :   35 - 0x23
    "00100011", -- 2887 - 0xb47  :   35 - 0x23
    "00000100", -- 2888 - 0xb48  :    4 - 0x4
    "00000100", -- 2889 - 0xb49  :    4 - 0x4
    "00000100", -- 2890 - 0xb4a  :    4 - 0x4
    "00000100", -- 2891 - 0xb4b  :    4 - 0x4
    "00000100", -- 2892 - 0xb4c  :    4 - 0x4
    "00000100", -- 2893 - 0xb4d  :    4 - 0x4
    "00000100", -- 2894 - 0xb4e  :    4 - 0x4
    "00000100", -- 2895 - 0xb4f  :    4 - 0x4
    "01000100", -- 2896 - 0xb50  :   68 - 0x44
    "10100100", -- 2897 - 0xb51  :  164 - 0xa4
    "01000100", -- 2898 - 0xb52  :   68 - 0x44
    "10100100", -- 2899 - 0xb53  :  164 - 0xa4
    "01000100", -- 2900 - 0xb54  :   68 - 0x44
    "10100100", -- 2901 - 0xb55  :  164 - 0xa4
    "01000100", -- 2902 - 0xb56  :   68 - 0x44
    "10100100", -- 2903 - 0xb57  :  164 - 0xa4
    "00011111", -- 2904 - 0xb58  :   31 - 0x1f
    "00111111", -- 2905 - 0xb59  :   63 - 0x3f
    "01111111", -- 2906 - 0xb5a  :  127 - 0x7f
    "01111111", -- 2907 - 0xb5b  :  127 - 0x7f
    "11111111", -- 2908 - 0xb5c  :  255 - 0xff
    "11111111", -- 2909 - 0xb5d  :  255 - 0xff
    "11111111", -- 2910 - 0xb5e  :  255 - 0xff
    "11111110", -- 2911 - 0xb5f  :  254 - 0xfe
    "11111111", -- 2912 - 0xb60  :  255 - 0xff
    "01111111", -- 2913 - 0xb61  :  127 - 0x7f
    "01111111", -- 2914 - 0xb62  :  127 - 0x7f
    "00111111", -- 2915 - 0xb63  :   63 - 0x3f
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000001", -- 2918 - 0xb66  :    1 - 0x1
    "00000001", -- 2919 - 0xb67  :    1 - 0x1
    "11111111", -- 2920 - 0xb68  :  255 - 0xff
    "10000000", -- 2921 - 0xb69  :  128 - 0x80
    "10000000", -- 2922 - 0xb6a  :  128 - 0x80
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "11111000", -- 2925 - 0xb6d  :  248 - 0xf8
    "11111100", -- 2926 - 0xb6e  :  252 - 0xfc
    "11111100", -- 2927 - 0xb6f  :  252 - 0xfc
    "11111111", -- 2928 - 0xb70  :  255 - 0xff
    "11111111", -- 2929 - 0xb71  :  255 - 0xff
    "11111111", -- 2930 - 0xb72  :  255 - 0xff
    "11111111", -- 2931 - 0xb73  :  255 - 0xff
    "11111111", -- 2932 - 0xb74  :  255 - 0xff
    "01111110", -- 2933 - 0xb75  :  126 - 0x7e
    "00111100", -- 2934 - 0xb76  :   60 - 0x3c
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "11111000", -- 2936 - 0xb78  :  248 - 0xf8
    "00000100", -- 2937 - 0xb79  :    4 - 0x4
    "00000010", -- 2938 - 0xb7a  :    2 - 0x2
    "00000010", -- 2939 - 0xb7b  :    2 - 0x2
    "00011101", -- 2940 - 0xb7c  :   29 - 0x1d
    "00111111", -- 2941 - 0xb7d  :   63 - 0x3f
    "01111111", -- 2942 - 0xb7e  :  127 - 0x7f
    "01111111", -- 2943 - 0xb7f  :  127 - 0x7f
    "11111100", -- 2944 - 0xb80  :  252 - 0xfc
    "10000000", -- 2945 - 0xb81  :  128 - 0x80
    "10000000", -- 2946 - 0xb82  :  128 - 0x80
    "10000000", -- 2947 - 0xb83  :  128 - 0x80
    "10000000", -- 2948 - 0xb84  :  128 - 0x80
    "10000000", -- 2949 - 0xb85  :  128 - 0x80
    "01100000", -- 2950 - 0xb86  :   96 - 0x60
    "00011111", -- 2951 - 0xb87  :   31 - 0x1f
    "00000011", -- 2952 - 0xb88  :    3 - 0x3
    "00000011", -- 2953 - 0xb89  :    3 - 0x3
    "00000011", -- 2954 - 0xb8a  :    3 - 0x3
    "00000011", -- 2955 - 0xb8b  :    3 - 0x3
    "00000001", -- 2956 - 0xb8c  :    1 - 0x1
    "00000001", -- 2957 - 0xb8d  :    1 - 0x1
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "11111111", -- 2959 - 0xb8f  :  255 - 0xff
    "11111110", -- 2960 - 0xb90  :  254 - 0xfe
    "11111110", -- 2961 - 0xb91  :  254 - 0xfe
    "11111110", -- 2962 - 0xb92  :  254 - 0xfe
    "11111110", -- 2963 - 0xb93  :  254 - 0xfe
    "11111100", -- 2964 - 0xb94  :  252 - 0xfc
    "11111100", -- 2965 - 0xb95  :  252 - 0xfc
    "11111000", -- 2966 - 0xb96  :  248 - 0xf8
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "00000000", -- 2968 - 0xb98  :    0 - 0x0
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "11111111", -- 2975 - 0xb9f  :  255 - 0xff
    "01111111", -- 2976 - 0xba0  :  127 - 0x7f
    "00111111", -- 2977 - 0xba1  :   63 - 0x3f
    "00011101", -- 2978 - 0xba2  :   29 - 0x1d
    "00000001", -- 2979 - 0xba3  :    1 - 0x1
    "00000001", -- 2980 - 0xba4  :    1 - 0x1
    "00000001", -- 2981 - 0xba5  :    1 - 0x1
    "00000011", -- 2982 - 0xba6  :    3 - 0x3
    "11111110", -- 2983 - 0xba7  :  254 - 0xfe
    "10000000", -- 2984 - 0xba8  :  128 - 0x80
    "10000000", -- 2985 - 0xba9  :  128 - 0x80
    "10000000", -- 2986 - 0xbaa  :  128 - 0x80
    "10000000", -- 2987 - 0xbab  :  128 - 0x80
    "10000000", -- 2988 - 0xbac  :  128 - 0x80
    "10000100", -- 2989 - 0xbad  :  132 - 0x84
    "11001010", -- 2990 - 0xbae  :  202 - 0xca
    "10110001", -- 2991 - 0xbaf  :  177 - 0xb1
    "00000001", -- 2992 - 0xbb0  :    1 - 0x1
    "00000001", -- 2993 - 0xbb1  :    1 - 0x1
    "00000001", -- 2994 - 0xbb2  :    1 - 0x1
    "00000001", -- 2995 - 0xbb3  :    1 - 0x1
    "00000001", -- 2996 - 0xbb4  :    1 - 0x1
    "00100001", -- 2997 - 0xbb5  :   33 - 0x21
    "01010011", -- 2998 - 0xbb6  :   83 - 0x53
    "10001101", -- 2999 - 0xbb7  :  141 - 0x8d
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "01110111", -- 3004 - 0xbbc  :  119 - 0x77
    "11111111", -- 3005 - 0xbbd  :  255 - 0xff
    "11111111", -- 3006 - 0xbbe  :  255 - 0xff
    "11111111", -- 3007 - 0xbbf  :  255 - 0xff
    "11111111", -- 3008 - 0xbc0  :  255 - 0xff
    "11111111", -- 3009 - 0xbc1  :  255 - 0xff
    "11111111", -- 3010 - 0xbc2  :  255 - 0xff
    "11111111", -- 3011 - 0xbc3  :  255 - 0xff
    "11111111", -- 3012 - 0xbc4  :  255 - 0xff
    "11111111", -- 3013 - 0xbc5  :  255 - 0xff
    "11111111", -- 3014 - 0xbc6  :  255 - 0xff
    "11111111", -- 3015 - 0xbc7  :  255 - 0xff
    "11111111", -- 3016 - 0xbc8  :  255 - 0xff
    "11111111", -- 3017 - 0xbc9  :  255 - 0xff
    "11111111", -- 3018 - 0xbca  :  255 - 0xff
    "01110111", -- 3019 - 0xbcb  :  119 - 0x77
    "01110111", -- 3020 - 0xbcc  :  119 - 0x77
    "01110111", -- 3021 - 0xbcd  :  119 - 0x77
    "01110111", -- 3022 - 0xbce  :  119 - 0x77
    "01110111", -- 3023 - 0xbcf  :  119 - 0x77
    "11111111", -- 3024 - 0xbd0  :  255 - 0xff
    "11111111", -- 3025 - 0xbd1  :  255 - 0xff
    "11111111", -- 3026 - 0xbd2  :  255 - 0xff
    "11100111", -- 3027 - 0xbd3  :  231 - 0xe7
    "11100111", -- 3028 - 0xbd4  :  231 - 0xe7
    "11111111", -- 3029 - 0xbd5  :  255 - 0xff
    "11111111", -- 3030 - 0xbd6  :  255 - 0xff
    "11111110", -- 3031 - 0xbd7  :  254 - 0xfe
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0
    "00100001", -- 3033 - 0xbd9  :   33 - 0x21
    "00100001", -- 3034 - 0xbda  :   33 - 0x21
    "01000001", -- 3035 - 0xbdb  :   65 - 0x41
    "01000001", -- 3036 - 0xbdc  :   65 - 0x41
    "01000001", -- 3037 - 0xbdd  :   65 - 0x41
    "01000001", -- 3038 - 0xbde  :   65 - 0x41
    "01000001", -- 3039 - 0xbdf  :   65 - 0x41
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0
    "10000000", -- 3041 - 0xbe1  :  128 - 0x80
    "10000000", -- 3042 - 0xbe2  :  128 - 0x80
    "10000000", -- 3043 - 0xbe3  :  128 - 0x80
    "10000000", -- 3044 - 0xbe4  :  128 - 0x80
    "10000000", -- 3045 - 0xbe5  :  128 - 0x80
    "10000000", -- 3046 - 0xbe6  :  128 - 0x80
    "10000000", -- 3047 - 0xbe7  :  128 - 0x80
    "00100001", -- 3048 - 0xbe8  :   33 - 0x21
    "00100001", -- 3049 - 0xbe9  :   33 - 0x21
    "00000001", -- 3050 - 0xbea  :    1 - 0x1
    "00000001", -- 3051 - 0xbeb  :    1 - 0x1
    "00000001", -- 3052 - 0xbec  :    1 - 0x1
    "00000001", -- 3053 - 0xbed  :    1 - 0x1
    "00000001", -- 3054 - 0xbee  :    1 - 0x1
    "00000001", -- 3055 - 0xbef  :    1 - 0x1
    "10000000", -- 3056 - 0xbf0  :  128 - 0x80
    "10000000", -- 3057 - 0xbf1  :  128 - 0x80
    "10000000", -- 3058 - 0xbf2  :  128 - 0x80
    "10000000", -- 3059 - 0xbf3  :  128 - 0x80
    "10000000", -- 3060 - 0xbf4  :  128 - 0x80
    "10000000", -- 3061 - 0xbf5  :  128 - 0x80
    "10000000", -- 3062 - 0xbf6  :  128 - 0x80
    "10000000", -- 3063 - 0xbf7  :  128 - 0x80
    "00000001", -- 3064 - 0xbf8  :    1 - 0x1
    "00000001", -- 3065 - 0xbf9  :    1 - 0x1
    "00000110", -- 3066 - 0xbfa  :    6 - 0x6
    "00001000", -- 3067 - 0xbfb  :    8 - 0x8
    "00011000", -- 3068 - 0xbfc  :   24 - 0x18
    "00100000", -- 3069 - 0xbfd  :   32 - 0x20
    "00100000", -- 3070 - 0xbfe  :   32 - 0x20
    "11000000", -- 3071 - 0xbff  :  192 - 0xc0
    "00000100", -- 3072 - 0xc00  :    4 - 0x4
    "00000100", -- 3073 - 0xc01  :    4 - 0x4
    "11000100", -- 3074 - 0xc02  :  196 - 0xc4
    "11110100", -- 3075 - 0xc03  :  244 - 0xf4
    "11110100", -- 3076 - 0xc04  :  244 - 0xf4
    "00000100", -- 3077 - 0xc05  :    4 - 0x4
    "00000100", -- 3078 - 0xc06  :    4 - 0x4
    "00000101", -- 3079 - 0xc07  :    5 - 0x5
    "01110000", -- 3080 - 0xc08  :  112 - 0x70
    "11110000", -- 3081 - 0xc09  :  240 - 0xf0
    "11110000", -- 3082 - 0xc0a  :  240 - 0xf0
    "11111111", -- 3083 - 0xc0b  :  255 - 0xff
    "11111111", -- 3084 - 0xc0c  :  255 - 0xff
    "11110000", -- 3085 - 0xc0d  :  240 - 0xf0
    "11110000", -- 3086 - 0xc0e  :  240 - 0xf0
    "01110000", -- 3087 - 0xc0f  :  112 - 0x70
    "11000000", -- 3088 - 0xc10  :  192 - 0xc0
    "10000111", -- 3089 - 0xc11  :  135 - 0x87
    "00011000", -- 3090 - 0xc12  :   24 - 0x18
    "10110000", -- 3091 - 0xc13  :  176 - 0xb0
    "11100111", -- 3092 - 0xc14  :  231 - 0xe7
    "11100111", -- 3093 - 0xc15  :  231 - 0xe7
    "11101111", -- 3094 - 0xc16  :  239 - 0xef
    "11101111", -- 3095 - 0xc17  :  239 - 0xef
    "01101111", -- 3096 - 0xc18  :  111 - 0x6f
    "01000011", -- 3097 - 0xc19  :   67 - 0x43
    "01011101", -- 3098 - 0xc1a  :   93 - 0x5d
    "00111111", -- 3099 - 0xc1b  :   63 - 0x3f
    "00111111", -- 3100 - 0xc1c  :   63 - 0x3f
    "01111111", -- 3101 - 0xc1d  :  127 - 0x7f
    "01111111", -- 3102 - 0xc1e  :  127 - 0x7f
    "11111111", -- 3103 - 0xc1f  :  255 - 0xff
    "00000011", -- 3104 - 0xc20  :    3 - 0x3
    "11111111", -- 3105 - 0xc21  :  255 - 0xff
    "11110001", -- 3106 - 0xc22  :  241 - 0xf1
    "01101110", -- 3107 - 0xc23  :  110 - 0x6e
    "11001111", -- 3108 - 0xc24  :  207 - 0xcf
    "11011111", -- 3109 - 0xc25  :  223 - 0xdf
    "11111111", -- 3110 - 0xc26  :  255 - 0xff
    "11111111", -- 3111 - 0xc27  :  255 - 0xff
    "11111101", -- 3112 - 0xc28  :  253 - 0xfd
    "11111011", -- 3113 - 0xc29  :  251 - 0xfb
    "11111011", -- 3114 - 0xc2a  :  251 - 0xfb
    "11110111", -- 3115 - 0xc2b  :  247 - 0xf7
    "11110111", -- 3116 - 0xc2c  :  247 - 0xf7
    "00001111", -- 3117 - 0xc2d  :   15 - 0xf
    "01111111", -- 3118 - 0xc2e  :  127 - 0x7f
    "11111111", -- 3119 - 0xc2f  :  255 - 0xff
    "11111111", -- 3120 - 0xc30  :  255 - 0xff
    "10000000", -- 3121 - 0xc31  :  128 - 0x80
    "10000000", -- 3122 - 0xc32  :  128 - 0x80
    "10000000", -- 3123 - 0xc33  :  128 - 0x80
    "10000000", -- 3124 - 0xc34  :  128 - 0x80
    "11111111", -- 3125 - 0xc35  :  255 - 0xff
    "11111111", -- 3126 - 0xc36  :  255 - 0xff
    "10000000", -- 3127 - 0xc37  :  128 - 0x80
    "11111110", -- 3128 - 0xc38  :  254 - 0xfe
    "00000011", -- 3129 - 0xc39  :    3 - 0x3
    "00000011", -- 3130 - 0xc3a  :    3 - 0x3
    "00000011", -- 3131 - 0xc3b  :    3 - 0x3
    "00000011", -- 3132 - 0xc3c  :    3 - 0x3
    "11111111", -- 3133 - 0xc3d  :  255 - 0xff
    "11111111", -- 3134 - 0xc3e  :  255 - 0xff
    "00000011", -- 3135 - 0xc3f  :    3 - 0x3
    "00000000", -- 3136 - 0xc40  :    0 - 0x0
    "11111111", -- 3137 - 0xc41  :  255 - 0xff
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "11111111", -- 3142 - 0xc46  :  255 - 0xff
    "11111111", -- 3143 - 0xc47  :  255 - 0xff
    "00100011", -- 3144 - 0xc48  :   35 - 0x23
    "11110011", -- 3145 - 0xc49  :  243 - 0xf3
    "00001011", -- 3146 - 0xc4a  :   11 - 0xb
    "00001011", -- 3147 - 0xc4b  :   11 - 0xb
    "00001011", -- 3148 - 0xc4c  :   11 - 0xb
    "00000111", -- 3149 - 0xc4d  :    7 - 0x7
    "11111111", -- 3150 - 0xc4e  :  255 - 0xff
    "11111111", -- 3151 - 0xc4f  :  255 - 0xff
    "10000000", -- 3152 - 0xc50  :  128 - 0x80
    "10000000", -- 3153 - 0xc51  :  128 - 0x80
    "10000000", -- 3154 - 0xc52  :  128 - 0x80
    "10000000", -- 3155 - 0xc53  :  128 - 0x80
    "11111111", -- 3156 - 0xc54  :  255 - 0xff
    "10000000", -- 3157 - 0xc55  :  128 - 0x80
    "10000000", -- 3158 - 0xc56  :  128 - 0x80
    "10000000", -- 3159 - 0xc57  :  128 - 0x80
    "00000011", -- 3160 - 0xc58  :    3 - 0x3
    "00000011", -- 3161 - 0xc59  :    3 - 0x3
    "00000011", -- 3162 - 0xc5a  :    3 - 0x3
    "00000011", -- 3163 - 0xc5b  :    3 - 0x3
    "11111111", -- 3164 - 0xc5c  :  255 - 0xff
    "00000011", -- 3165 - 0xc5d  :    3 - 0x3
    "00000011", -- 3166 - 0xc5e  :    3 - 0x3
    "00000011", -- 3167 - 0xc5f  :    3 - 0x3
    "00000000", -- 3168 - 0xc60  :    0 - 0x0
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "11111111", -- 3173 - 0xc65  :  255 - 0xff
    "00000000", -- 3174 - 0xc66  :    0 - 0x0
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000111", -- 3176 - 0xc68  :    7 - 0x7
    "00000111", -- 3177 - 0xc69  :    7 - 0x7
    "00000011", -- 3178 - 0xc6a  :    3 - 0x3
    "00000011", -- 3179 - 0xc6b  :    3 - 0x3
    "00000011", -- 3180 - 0xc6c  :    3 - 0x3
    "11111111", -- 3181 - 0xc6d  :  255 - 0xff
    "00000011", -- 3182 - 0xc6e  :    3 - 0x3
    "00000011", -- 3183 - 0xc6f  :    3 - 0x3
    "10000000", -- 3184 - 0xc70  :  128 - 0x80
    "11111111", -- 3185 - 0xc71  :  255 - 0xff
    "11111111", -- 3186 - 0xc72  :  255 - 0xff
    "11111111", -- 3187 - 0xc73  :  255 - 0xff
    "11111111", -- 3188 - 0xc74  :  255 - 0xff
    "11111111", -- 3189 - 0xc75  :  255 - 0xff
    "11111111", -- 3190 - 0xc76  :  255 - 0xff
    "11111111", -- 3191 - 0xc77  :  255 - 0xff
    "00000011", -- 3192 - 0xc78  :    3 - 0x3
    "11111111", -- 3193 - 0xc79  :  255 - 0xff
    "11111111", -- 3194 - 0xc7a  :  255 - 0xff
    "11111111", -- 3195 - 0xc7b  :  255 - 0xff
    "11111111", -- 3196 - 0xc7c  :  255 - 0xff
    "11111111", -- 3197 - 0xc7d  :  255 - 0xff
    "11111111", -- 3198 - 0xc7e  :  255 - 0xff
    "11111111", -- 3199 - 0xc7f  :  255 - 0xff
    "11111111", -- 3200 - 0xc80  :  255 - 0xff
    "11111111", -- 3201 - 0xc81  :  255 - 0xff
    "11111111", -- 3202 - 0xc82  :  255 - 0xff
    "11111111", -- 3203 - 0xc83  :  255 - 0xff
    "11111111", -- 3204 - 0xc84  :  255 - 0xff
    "11111111", -- 3205 - 0xc85  :  255 - 0xff
    "11111111", -- 3206 - 0xc86  :  255 - 0xff
    "11111111", -- 3207 - 0xc87  :  255 - 0xff
    "11111111", -- 3208 - 0xc88  :  255 - 0xff
    "11111111", -- 3209 - 0xc89  :  255 - 0xff
    "11010101", -- 3210 - 0xc8a  :  213 - 0xd5
    "10101010", -- 3211 - 0xc8b  :  170 - 0xaa
    "11010101", -- 3212 - 0xc8c  :  213 - 0xd5
    "10000000", -- 3213 - 0xc8d  :  128 - 0x80
    "10000000", -- 3214 - 0xc8e  :  128 - 0x80
    "11111111", -- 3215 - 0xc8f  :  255 - 0xff
    "11111111", -- 3216 - 0xc90  :  255 - 0xff
    "11111111", -- 3217 - 0xc91  :  255 - 0xff
    "01010111", -- 3218 - 0xc92  :   87 - 0x57
    "10101011", -- 3219 - 0xc93  :  171 - 0xab
    "01010111", -- 3220 - 0xc94  :   87 - 0x57
    "00000011", -- 3221 - 0xc95  :    3 - 0x3
    "00000011", -- 3222 - 0xc96  :    3 - 0x3
    "11111110", -- 3223 - 0xc97  :  254 - 0xfe
    "11111111", -- 3224 - 0xc98  :  255 - 0xff
    "10101010", -- 3225 - 0xc99  :  170 - 0xaa
    "01010101", -- 3226 - 0xc9a  :   85 - 0x55
    "10101010", -- 3227 - 0xc9b  :  170 - 0xaa
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "11111111", -- 3230 - 0xc9e  :  255 - 0xff
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "11111111", -- 3232 - 0xca0  :  255 - 0xff
    "10101111", -- 3233 - 0xca1  :  175 - 0xaf
    "01010111", -- 3234 - 0xca2  :   87 - 0x57
    "10101011", -- 3235 - 0xca3  :  171 - 0xab
    "00001011", -- 3236 - 0xca4  :   11 - 0xb
    "00001011", -- 3237 - 0xca5  :   11 - 0xb
    "11110011", -- 3238 - 0xca6  :  243 - 0xf3
    "00100011", -- 3239 - 0xca7  :   35 - 0x23
    "11111111", -- 3240 - 0xca8  :  255 - 0xff
    "11111111", -- 3241 - 0xca9  :  255 - 0xff
    "11111111", -- 3242 - 0xcaa  :  255 - 0xff
    "11111111", -- 3243 - 0xcab  :  255 - 0xff
    "11111111", -- 3244 - 0xcac  :  255 - 0xff
    "11111111", -- 3245 - 0xcad  :  255 - 0xff
    "11111111", -- 3246 - 0xcae  :  255 - 0xff
    "11111111", -- 3247 - 0xcaf  :  255 - 0xff
    "11111111", -- 3248 - 0xcb0  :  255 - 0xff
    "11111111", -- 3249 - 0xcb1  :  255 - 0xff
    "11111111", -- 3250 - 0xcb2  :  255 - 0xff
    "11111111", -- 3251 - 0xcb3  :  255 - 0xff
    "11111111", -- 3252 - 0xcb4  :  255 - 0xff
    "11111111", -- 3253 - 0xcb5  :  255 - 0xff
    "11111111", -- 3254 - 0xcb6  :  255 - 0xff
    "11111111", -- 3255 - 0xcb7  :  255 - 0xff
    "11111111", -- 3256 - 0xcb8  :  255 - 0xff
    "11111111", -- 3257 - 0xcb9  :  255 - 0xff
    "11111111", -- 3258 - 0xcba  :  255 - 0xff
    "11111111", -- 3259 - 0xcbb  :  255 - 0xff
    "11111111", -- 3260 - 0xcbc  :  255 - 0xff
    "11111111", -- 3261 - 0xcbd  :  255 - 0xff
    "11111111", -- 3262 - 0xcbe  :  255 - 0xff
    "11111111", -- 3263 - 0xcbf  :  255 - 0xff
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff
    "11111111", -- 3265 - 0xcc1  :  255 - 0xff
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111111", -- 3267 - 0xcc3  :  255 - 0xff
    "11111111", -- 3268 - 0xcc4  :  255 - 0xff
    "11111111", -- 3269 - 0xcc5  :  255 - 0xff
    "11111111", -- 3270 - 0xcc6  :  255 - 0xff
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "11111111", -- 3288 - 0xcd8  :  255 - 0xff
    "11111111", -- 3289 - 0xcd9  :  255 - 0xff
    "11111111", -- 3290 - 0xcda  :  255 - 0xff
    "11111111", -- 3291 - 0xcdb  :  255 - 0xff
    "11111111", -- 3292 - 0xcdc  :  255 - 0xff
    "11111111", -- 3293 - 0xcdd  :  255 - 0xff
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "11111111", -- 3296 - 0xce0  :  255 - 0xff
    "11111111", -- 3297 - 0xce1  :  255 - 0xff
    "11111111", -- 3298 - 0xce2  :  255 - 0xff
    "11111111", -- 3299 - 0xce3  :  255 - 0xff
    "11111111", -- 3300 - 0xce4  :  255 - 0xff
    "11111111", -- 3301 - 0xce5  :  255 - 0xff
    "11111111", -- 3302 - 0xce6  :  255 - 0xff
    "11111111", -- 3303 - 0xce7  :  255 - 0xff
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "11100000", -- 3305 - 0xce9  :  224 - 0xe0
    "11100000", -- 3306 - 0xcea  :  224 - 0xe0
    "11100000", -- 3307 - 0xceb  :  224 - 0xe0
    "11100000", -- 3308 - 0xcec  :  224 - 0xe0
    "11100000", -- 3309 - 0xced  :  224 - 0xe0
    "11100000", -- 3310 - 0xcee  :  224 - 0xe0
    "11100000", -- 3311 - 0xcef  :  224 - 0xe0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0
    "00001111", -- 3313 - 0xcf1  :   15 - 0xf
    "00001111", -- 3314 - 0xcf2  :   15 - 0xf
    "00001111", -- 3315 - 0xcf3  :   15 - 0xf
    "00001111", -- 3316 - 0xcf4  :   15 - 0xf
    "00001111", -- 3317 - 0xcf5  :   15 - 0xf
    "00001111", -- 3318 - 0xcf6  :   15 - 0xf
    "00001111", -- 3319 - 0xcf7  :   15 - 0xf
    "01001000", -- 3320 - 0xcf8  :   72 - 0x48
    "01001000", -- 3321 - 0xcf9  :   72 - 0x48
    "01101100", -- 3322 - 0xcfa  :  108 - 0x6c
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "11111110", -- 3326 - 0xcfe  :  254 - 0xfe
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000101", -- 3328 - 0xd00  :    5 - 0x5
    "00000101", -- 3329 - 0xd01  :    5 - 0x5
    "11000101", -- 3330 - 0xd02  :  197 - 0xc5
    "11110101", -- 3331 - 0xd03  :  245 - 0xf5
    "11110100", -- 3332 - 0xd04  :  244 - 0xf4
    "00000100", -- 3333 - 0xd05  :    4 - 0x4
    "00000100", -- 3334 - 0xd06  :    4 - 0x4
    "00000100", -- 3335 - 0xd07  :    4 - 0x4
    "01110000", -- 3336 - 0xd08  :  112 - 0x70
    "01110000", -- 3337 - 0xd09  :  112 - 0x70
    "01110000", -- 3338 - 0xd0a  :  112 - 0x70
    "01111111", -- 3339 - 0xd0b  :  127 - 0x7f
    "01111111", -- 3340 - 0xd0c  :  127 - 0x7f
    "01110000", -- 3341 - 0xd0d  :  112 - 0x70
    "01110000", -- 3342 - 0xd0e  :  112 - 0x70
    "01110000", -- 3343 - 0xd0f  :  112 - 0x70
    "00000000", -- 3344 - 0xd10  :    0 - 0x0
    "00000000", -- 3345 - 0xd11  :    0 - 0x0
    "00000000", -- 3346 - 0xd12  :    0 - 0x0
    "00000000", -- 3347 - 0xd13  :    0 - 0x0
    "00000000", -- 3348 - 0xd14  :    0 - 0x0
    "00000000", -- 3349 - 0xd15  :    0 - 0x0
    "00000000", -- 3350 - 0xd16  :    0 - 0x0
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "11111111", -- 3360 - 0xd20  :  255 - 0xff
    "11111111", -- 3361 - 0xd21  :  255 - 0xff
    "11111111", -- 3362 - 0xd22  :  255 - 0xff
    "11111111", -- 3363 - 0xd23  :  255 - 0xff
    "11111111", -- 3364 - 0xd24  :  255 - 0xff
    "11111110", -- 3365 - 0xd25  :  254 - 0xfe
    "10111110", -- 3366 - 0xd26  :  190 - 0xbe
    "11001110", -- 3367 - 0xd27  :  206 - 0xce
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000011", -- 3372 - 0xd2c  :    3 - 0x3
    "00000100", -- 3373 - 0xd2d  :    4 - 0x4
    "00000100", -- 3374 - 0xd2e  :    4 - 0x4
    "00000100", -- 3375 - 0xd2f  :    4 - 0x4
    "00000000", -- 3376 - 0xd30  :    0 - 0x0
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "01100000", -- 3378 - 0xd32  :   96 - 0x60
    "00110000", -- 3379 - 0xd33  :   48 - 0x30
    "00110000", -- 3380 - 0xd34  :   48 - 0x30
    "10011000", -- 3381 - 0xd35  :  152 - 0x98
    "10011000", -- 3382 - 0xd36  :  152 - 0x98
    "10011000", -- 3383 - 0xd37  :  152 - 0x98
    "00000100", -- 3384 - 0xd38  :    4 - 0x4
    "00000100", -- 3385 - 0xd39  :    4 - 0x4
    "00000100", -- 3386 - 0xd3a  :    4 - 0x4
    "00000100", -- 3387 - 0xd3b  :    4 - 0x4
    "00000100", -- 3388 - 0xd3c  :    4 - 0x4
    "00000011", -- 3389 - 0xd3d  :    3 - 0x3
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "10011000", -- 3392 - 0xd40  :  152 - 0x98
    "10011000", -- 3393 - 0xd41  :  152 - 0x98
    "10011000", -- 3394 - 0xd42  :  152 - 0x98
    "10011000", -- 3395 - 0xd43  :  152 - 0x98
    "10011000", -- 3396 - 0xd44  :  152 - 0x98
    "00110000", -- 3397 - 0xd45  :   48 - 0x30
    "00110000", -- 3398 - 0xd46  :   48 - 0x30
    "01100000", -- 3399 - 0xd47  :   96 - 0x60
    "00001111", -- 3400 - 0xd48  :   15 - 0xf
    "11101111", -- 3401 - 0xd49  :  239 - 0xef
    "11101111", -- 3402 - 0xd4a  :  239 - 0xef
    "11101111", -- 3403 - 0xd4b  :  239 - 0xef
    "11101111", -- 3404 - 0xd4c  :  239 - 0xef
    "11101111", -- 3405 - 0xd4d  :  239 - 0xef
    "11101111", -- 3406 - 0xd4e  :  239 - 0xef
    "11100000", -- 3407 - 0xd4f  :  224 - 0xe0
    "11100000", -- 3408 - 0xd50  :  224 - 0xe0
    "11101111", -- 3409 - 0xd51  :  239 - 0xef
    "11101111", -- 3410 - 0xd52  :  239 - 0xef
    "11101111", -- 3411 - 0xd53  :  239 - 0xef
    "11101111", -- 3412 - 0xd54  :  239 - 0xef
    "11101111", -- 3413 - 0xd55  :  239 - 0xef
    "11101111", -- 3414 - 0xd56  :  239 - 0xef
    "00001111", -- 3415 - 0xd57  :   15 - 0xf
    "10000000", -- 3416 - 0xd58  :  128 - 0x80
    "01000000", -- 3417 - 0xd59  :   64 - 0x40
    "00100000", -- 3418 - 0xd5a  :   32 - 0x20
    "00010000", -- 3419 - 0xd5b  :   16 - 0x10
    "00001111", -- 3420 - 0xd5c  :   15 - 0xf
    "00001111", -- 3421 - 0xd5d  :   15 - 0xf
    "00001111", -- 3422 - 0xd5e  :   15 - 0xf
    "00001111", -- 3423 - 0xd5f  :   15 - 0xf
    "00001111", -- 3424 - 0xd60  :   15 - 0xf
    "00001111", -- 3425 - 0xd61  :   15 - 0xf
    "00001111", -- 3426 - 0xd62  :   15 - 0xf
    "00001111", -- 3427 - 0xd63  :   15 - 0xf
    "00011111", -- 3428 - 0xd64  :   31 - 0x1f
    "00111111", -- 3429 - 0xd65  :   63 - 0x3f
    "01111111", -- 3430 - 0xd66  :  127 - 0x7f
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "00000001", -- 3432 - 0xd68  :    1 - 0x1
    "00000011", -- 3433 - 0xd69  :    3 - 0x3
    "00000111", -- 3434 - 0xd6a  :    7 - 0x7
    "00001111", -- 3435 - 0xd6b  :   15 - 0xf
    "11111111", -- 3436 - 0xd6c  :  255 - 0xff
    "11111111", -- 3437 - 0xd6d  :  255 - 0xff
    "11111111", -- 3438 - 0xd6e  :  255 - 0xff
    "11111111", -- 3439 - 0xd6f  :  255 - 0xff
    "11111111", -- 3440 - 0xd70  :  255 - 0xff
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "11111111", -- 3442 - 0xd72  :  255 - 0xff
    "11111111", -- 3443 - 0xd73  :  255 - 0xff
    "11111111", -- 3444 - 0xd74  :  255 - 0xff
    "11111111", -- 3445 - 0xd75  :  255 - 0xff
    "11111111", -- 3446 - 0xd76  :  255 - 0xff
    "11111111", -- 3447 - 0xd77  :  255 - 0xff
    "00000000", -- 3448 - 0xd78  :    0 - 0x0
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "00000000", -- 3451 - 0xd7b  :    0 - 0x0
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "00011111", -- 3456 - 0xd80  :   31 - 0x1f
    "00100000", -- 3457 - 0xd81  :   32 - 0x20
    "01000000", -- 3458 - 0xd82  :   64 - 0x40
    "01000000", -- 3459 - 0xd83  :   64 - 0x40
    "01000000", -- 3460 - 0xd84  :   64 - 0x40
    "10000000", -- 3461 - 0xd85  :  128 - 0x80
    "10000010", -- 3462 - 0xd86  :  130 - 0x82
    "10000010", -- 3463 - 0xd87  :  130 - 0x82
    "10000010", -- 3464 - 0xd88  :  130 - 0x82
    "10000000", -- 3465 - 0xd89  :  128 - 0x80
    "10100000", -- 3466 - 0xd8a  :  160 - 0xa0
    "01000100", -- 3467 - 0xd8b  :   68 - 0x44
    "01000011", -- 3468 - 0xd8c  :   67 - 0x43
    "01000000", -- 3469 - 0xd8d  :   64 - 0x40
    "00100001", -- 3470 - 0xd8e  :   33 - 0x21
    "00011110", -- 3471 - 0xd8f  :   30 - 0x1e
    "11111000", -- 3472 - 0xd90  :  248 - 0xf8
    "00000100", -- 3473 - 0xd91  :    4 - 0x4
    "00000010", -- 3474 - 0xd92  :    2 - 0x2
    "00000010", -- 3475 - 0xd93  :    2 - 0x2
    "00000010", -- 3476 - 0xd94  :    2 - 0x2
    "00000001", -- 3477 - 0xd95  :    1 - 0x1
    "01000001", -- 3478 - 0xd96  :   65 - 0x41
    "01000001", -- 3479 - 0xd97  :   65 - 0x41
    "01000001", -- 3480 - 0xd98  :   65 - 0x41
    "00000001", -- 3481 - 0xd99  :    1 - 0x1
    "00000101", -- 3482 - 0xd9a  :    5 - 0x5
    "00100010", -- 3483 - 0xd9b  :   34 - 0x22
    "11000010", -- 3484 - 0xd9c  :  194 - 0xc2
    "00000010", -- 3485 - 0xd9d  :    2 - 0x2
    "10000100", -- 3486 - 0xd9e  :  132 - 0x84
    "01111000", -- 3487 - 0xd9f  :  120 - 0x78
    "10000000", -- 3488 - 0xda0  :  128 - 0x80
    "01111111", -- 3489 - 0xda1  :  127 - 0x7f
    "01111111", -- 3490 - 0xda2  :  127 - 0x7f
    "01111111", -- 3491 - 0xda3  :  127 - 0x7f
    "01111111", -- 3492 - 0xda4  :  127 - 0x7f
    "01111111", -- 3493 - 0xda5  :  127 - 0x7f
    "01111111", -- 3494 - 0xda6  :  127 - 0x7f
    "01111111", -- 3495 - 0xda7  :  127 - 0x7f
    "01100001", -- 3496 - 0xda8  :   97 - 0x61
    "11011111", -- 3497 - 0xda9  :  223 - 0xdf
    "11011111", -- 3498 - 0xdaa  :  223 - 0xdf
    "11011111", -- 3499 - 0xdab  :  223 - 0xdf
    "11011111", -- 3500 - 0xdac  :  223 - 0xdf
    "11111111", -- 3501 - 0xdad  :  255 - 0xff
    "11000001", -- 3502 - 0xdae  :  193 - 0xc1
    "11011111", -- 3503 - 0xdaf  :  223 - 0xdf
    "01111111", -- 3504 - 0xdb0  :  127 - 0x7f
    "01111111", -- 3505 - 0xdb1  :  127 - 0x7f
    "11111111", -- 3506 - 0xdb2  :  255 - 0xff
    "00111111", -- 3507 - 0xdb3  :   63 - 0x3f
    "01001111", -- 3508 - 0xdb4  :   79 - 0x4f
    "01110001", -- 3509 - 0xdb5  :  113 - 0x71
    "01111111", -- 3510 - 0xdb6  :  127 - 0x7f
    "11111111", -- 3511 - 0xdb7  :  255 - 0xff
    "11011111", -- 3512 - 0xdb8  :  223 - 0xdf
    "11011111", -- 3513 - 0xdb9  :  223 - 0xdf
    "10111111", -- 3514 - 0xdba  :  191 - 0xbf
    "10111111", -- 3515 - 0xdbb  :  191 - 0xbf
    "01111111", -- 3516 - 0xdbc  :  127 - 0x7f
    "01111111", -- 3517 - 0xdbd  :  127 - 0x7f
    "01111111", -- 3518 - 0xdbe  :  127 - 0x7f
    "01111111", -- 3519 - 0xdbf  :  127 - 0x7f
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000011", -- 3522 - 0xdc2  :    3 - 0x3
    "00001100", -- 3523 - 0xdc3  :   12 - 0xc
    "00010000", -- 3524 - 0xdc4  :   16 - 0x10
    "00100000", -- 3525 - 0xdc5  :   32 - 0x20
    "01000000", -- 3526 - 0xdc6  :   64 - 0x40
    "01000000", -- 3527 - 0xdc7  :   64 - 0x40
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "11000000", -- 3530 - 0xdca  :  192 - 0xc0
    "00110000", -- 3531 - 0xdcb  :   48 - 0x30
    "00001000", -- 3532 - 0xdcc  :    8 - 0x8
    "00000100", -- 3533 - 0xdcd  :    4 - 0x4
    "00000010", -- 3534 - 0xdce  :    2 - 0x2
    "00000010", -- 3535 - 0xdcf  :    2 - 0x2
    "10000000", -- 3536 - 0xdd0  :  128 - 0x80
    "10000000", -- 3537 - 0xdd1  :  128 - 0x80
    "10000000", -- 3538 - 0xdd2  :  128 - 0x80
    "10000000", -- 3539 - 0xdd3  :  128 - 0x80
    "10000000", -- 3540 - 0xdd4  :  128 - 0x80
    "10000000", -- 3541 - 0xdd5  :  128 - 0x80
    "10000000", -- 3542 - 0xdd6  :  128 - 0x80
    "10000000", -- 3543 - 0xdd7  :  128 - 0x80
    "00000001", -- 3544 - 0xdd8  :    1 - 0x1
    "00000001", -- 3545 - 0xdd9  :    1 - 0x1
    "00000001", -- 3546 - 0xdda  :    1 - 0x1
    "00000001", -- 3547 - 0xddb  :    1 - 0x1
    "00000001", -- 3548 - 0xddc  :    1 - 0x1
    "00000001", -- 3549 - 0xddd  :    1 - 0x1
    "00000001", -- 3550 - 0xdde  :    1 - 0x1
    "00000001", -- 3551 - 0xddf  :    1 - 0x1
    "01000000", -- 3552 - 0xde0  :   64 - 0x40
    "01000000", -- 3553 - 0xde1  :   64 - 0x40
    "01000000", -- 3554 - 0xde2  :   64 - 0x40
    "00100000", -- 3555 - 0xde3  :   32 - 0x20
    "00110000", -- 3556 - 0xde4  :   48 - 0x30
    "00011100", -- 3557 - 0xde5  :   28 - 0x1c
    "00001111", -- 3558 - 0xde6  :   15 - 0xf
    "00000111", -- 3559 - 0xde7  :    7 - 0x7
    "00000010", -- 3560 - 0xde8  :    2 - 0x2
    "00000010", -- 3561 - 0xde9  :    2 - 0x2
    "00000010", -- 3562 - 0xdea  :    2 - 0x2
    "00000100", -- 3563 - 0xdeb  :    4 - 0x4
    "00001100", -- 3564 - 0xdec  :   12 - 0xc
    "00111000", -- 3565 - 0xded  :   56 - 0x38
    "11110000", -- 3566 - 0xdee  :  240 - 0xf0
    "11110000", -- 3567 - 0xdef  :  240 - 0xf0
    "00001000", -- 3568 - 0xdf0  :    8 - 0x8
    "00001000", -- 3569 - 0xdf1  :    8 - 0x8
    "00001000", -- 3570 - 0xdf2  :    8 - 0x8
    "00001000", -- 3571 - 0xdf3  :    8 - 0x8
    "00001000", -- 3572 - 0xdf4  :    8 - 0x8
    "00001100", -- 3573 - 0xdf5  :   12 - 0xc
    "00000101", -- 3574 - 0xdf6  :    5 - 0x5
    "00001010", -- 3575 - 0xdf7  :   10 - 0xa
    "00010000", -- 3576 - 0xdf8  :   16 - 0x10
    "01010000", -- 3577 - 0xdf9  :   80 - 0x50
    "01010000", -- 3578 - 0xdfa  :   80 - 0x50
    "01010000", -- 3579 - 0xdfb  :   80 - 0x50
    "01010000", -- 3580 - 0xdfc  :   80 - 0x50
    "00110000", -- 3581 - 0xdfd  :   48 - 0x30
    "10100000", -- 3582 - 0xdfe  :  160 - 0xa0
    "01010000", -- 3583 - 0xdff  :   80 - 0x50
    "00000000", -- 3584 - 0xe00  :    0 - 0x0
    "01000001", -- 3585 - 0xe01  :   65 - 0x41
    "00100010", -- 3586 - 0xe02  :   34 - 0x22
    "00100010", -- 3587 - 0xe03  :   34 - 0x22
    "00011100", -- 3588 - 0xe04  :   28 - 0x1c
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "11100011", -- 3592 - 0xe08  :  227 - 0xe3
    "00010100", -- 3593 - 0xe09  :   20 - 0x14
    "00111110", -- 3594 - 0xe0a  :   62 - 0x3e
    "00111110", -- 3595 - 0xe0b  :   62 - 0x3e
    "00111110", -- 3596 - 0xe0c  :   62 - 0x3e
    "00111110", -- 3597 - 0xe0d  :   62 - 0x3e
    "00010100", -- 3598 - 0xe0e  :   20 - 0x14
    "11100011", -- 3599 - 0xe0f  :  227 - 0xe3
    "11111111", -- 3600 - 0xe10  :  255 - 0xff
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "11111000", -- 3602 - 0xe12  :  248 - 0xf8
    "11110000", -- 3603 - 0xe13  :  240 - 0xf0
    "11110000", -- 3604 - 0xe14  :  240 - 0xf0
    "11100000", -- 3605 - 0xe15  :  224 - 0xe0
    "11100000", -- 3606 - 0xe16  :  224 - 0xe0
    "11100000", -- 3607 - 0xe17  :  224 - 0xe0
    "11111111", -- 3608 - 0xe18  :  255 - 0xff
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "01111111", -- 3610 - 0xe1a  :  127 - 0x7f
    "00111111", -- 3611 - 0xe1b  :   63 - 0x3f
    "00111111", -- 3612 - 0xe1c  :   63 - 0x3f
    "10011111", -- 3613 - 0xe1d  :  159 - 0x9f
    "10011111", -- 3614 - 0xe1e  :  159 - 0x9f
    "10011111", -- 3615 - 0xe1f  :  159 - 0x9f
    "11100000", -- 3616 - 0xe20  :  224 - 0xe0
    "11100000", -- 3617 - 0xe21  :  224 - 0xe0
    "11100000", -- 3618 - 0xe22  :  224 - 0xe0
    "11100000", -- 3619 - 0xe23  :  224 - 0xe0
    "11100000", -- 3620 - 0xe24  :  224 - 0xe0
    "11110011", -- 3621 - 0xe25  :  243 - 0xf3
    "11110000", -- 3622 - 0xe26  :  240 - 0xf0
    "11111000", -- 3623 - 0xe27  :  248 - 0xf8
    "10011111", -- 3624 - 0xe28  :  159 - 0x9f
    "10011111", -- 3625 - 0xe29  :  159 - 0x9f
    "10011111", -- 3626 - 0xe2a  :  159 - 0x9f
    "10011111", -- 3627 - 0xe2b  :  159 - 0x9f
    "10011111", -- 3628 - 0xe2c  :  159 - 0x9f
    "00111111", -- 3629 - 0xe2d  :   63 - 0x3f
    "00111111", -- 3630 - 0xe2e  :   63 - 0x3f
    "01111111", -- 3631 - 0xe2f  :  127 - 0x7f
    "00000000", -- 3632 - 0xe30  :    0 - 0x0
    "01110000", -- 3633 - 0xe31  :  112 - 0x70
    "00011111", -- 3634 - 0xe32  :   31 - 0x1f
    "00010000", -- 3635 - 0xe33  :   16 - 0x10
    "01110000", -- 3636 - 0xe34  :  112 - 0x70
    "01111111", -- 3637 - 0xe35  :  127 - 0x7f
    "01111111", -- 3638 - 0xe36  :  127 - 0x7f
    "01111111", -- 3639 - 0xe37  :  127 - 0x7f
    "00000000", -- 3640 - 0xe38  :    0 - 0x0
    "00000011", -- 3641 - 0xe39  :    3 - 0x3
    "11111000", -- 3642 - 0xe3a  :  248 - 0xf8
    "00000000", -- 3643 - 0xe3b  :    0 - 0x0
    "00000011", -- 3644 - 0xe3c  :    3 - 0x3
    "11111011", -- 3645 - 0xe3d  :  251 - 0xfb
    "11111011", -- 3646 - 0xe3e  :  251 - 0xfb
    "11111011", -- 3647 - 0xe3f  :  251 - 0xfb
    "01111100", -- 3648 - 0xe40  :  124 - 0x7c
    "01111011", -- 3649 - 0xe41  :  123 - 0x7b
    "01110110", -- 3650 - 0xe42  :  118 - 0x76
    "01110101", -- 3651 - 0xe43  :  117 - 0x75
    "01110101", -- 3652 - 0xe44  :  117 - 0x75
    "01110111", -- 3653 - 0xe45  :  119 - 0x77
    "00010111", -- 3654 - 0xe46  :   23 - 0x17
    "01100111", -- 3655 - 0xe47  :  103 - 0x67
    "00111011", -- 3656 - 0xe48  :   59 - 0x3b
    "11111011", -- 3657 - 0xe49  :  251 - 0xfb
    "01111011", -- 3658 - 0xe4a  :  123 - 0x7b
    "11111011", -- 3659 - 0xe4b  :  251 - 0xfb
    "11111011", -- 3660 - 0xe4c  :  251 - 0xfb
    "11110011", -- 3661 - 0xe4d  :  243 - 0xf3
    "11111000", -- 3662 - 0xe4e  :  248 - 0xf8
    "11110011", -- 3663 - 0xe4f  :  243 - 0xf3
    "00001111", -- 3664 - 0xe50  :   15 - 0xf
    "00001111", -- 3665 - 0xe51  :   15 - 0xf
    "00011111", -- 3666 - 0xe52  :   31 - 0x1f
    "00011111", -- 3667 - 0xe53  :   31 - 0x1f
    "00111111", -- 3668 - 0xe54  :   63 - 0x3f
    "00111100", -- 3669 - 0xe55  :   60 - 0x3c
    "01111000", -- 3670 - 0xe56  :  120 - 0x78
    "01111010", -- 3671 - 0xe57  :  122 - 0x7a
    "11111000", -- 3672 - 0xe58  :  248 - 0xf8
    "11111000", -- 3673 - 0xe59  :  248 - 0xf8
    "11111100", -- 3674 - 0xe5a  :  252 - 0xfc
    "11111100", -- 3675 - 0xe5b  :  252 - 0xfc
    "11111110", -- 3676 - 0xe5c  :  254 - 0xfe
    "00111110", -- 3677 - 0xe5d  :   62 - 0x3e
    "00011110", -- 3678 - 0xe5e  :   30 - 0x1e
    "01011111", -- 3679 - 0xe5f  :   95 - 0x5f
    "01110110", -- 3680 - 0xe60  :  118 - 0x76
    "01110110", -- 3681 - 0xe61  :  118 - 0x76
    "01110110", -- 3682 - 0xe62  :  118 - 0x76
    "01110000", -- 3683 - 0xe63  :  112 - 0x70
    "01111101", -- 3684 - 0xe64  :  125 - 0x7d
    "01111100", -- 3685 - 0xe65  :  124 - 0x7c
    "01111111", -- 3686 - 0xe66  :  127 - 0x7f
    "01111111", -- 3687 - 0xe67  :  127 - 0x7f
    "01101111", -- 3688 - 0xe68  :  111 - 0x6f
    "01101111", -- 3689 - 0xe69  :  111 - 0x6f
    "01101111", -- 3690 - 0xe6a  :  111 - 0x6f
    "00001111", -- 3691 - 0xe6b  :   15 - 0xf
    "10111111", -- 3692 - 0xe6c  :  191 - 0xbf
    "00111111", -- 3693 - 0xe6d  :   63 - 0x3f
    "11111111", -- 3694 - 0xe6e  :  255 - 0xff
    "11111111", -- 3695 - 0xe6f  :  255 - 0xff
    "00111100", -- 3696 - 0xe70  :   60 - 0x3c
    "01111110", -- 3697 - 0xe71  :  126 - 0x7e
    "01111110", -- 3698 - 0xe72  :  126 - 0x7e
    "11111111", -- 3699 - 0xe73  :  255 - 0xff
    "11111111", -- 3700 - 0xe74  :  255 - 0xff
    "11111111", -- 3701 - 0xe75  :  255 - 0xff
    "01000010", -- 3702 - 0xe76  :   66 - 0x42
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00000000", -- 3704 - 0xe78  :    0 - 0x0
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "11110000", -- 3712 - 0xe80  :  240 - 0xf0
    "11100000", -- 3713 - 0xe81  :  224 - 0xe0
    "11100000", -- 3714 - 0xe82  :  224 - 0xe0
    "11000000", -- 3715 - 0xe83  :  192 - 0xc0
    "11000000", -- 3716 - 0xe84  :  192 - 0xc0
    "10000000", -- 3717 - 0xe85  :  128 - 0x80
    "10000000", -- 3718 - 0xe86  :  128 - 0x80
    "10000000", -- 3719 - 0xe87  :  128 - 0x80
    "00001111", -- 3720 - 0xe88  :   15 - 0xf
    "00000111", -- 3721 - 0xe89  :    7 - 0x7
    "00000111", -- 3722 - 0xe8a  :    7 - 0x7
    "00000011", -- 3723 - 0xe8b  :    3 - 0x3
    "00000011", -- 3724 - 0xe8c  :    3 - 0x3
    "00000001", -- 3725 - 0xe8d  :    1 - 0x1
    "00000001", -- 3726 - 0xe8e  :    1 - 0x1
    "00000001", -- 3727 - 0xe8f  :    1 - 0x1
    "10000000", -- 3728 - 0xe90  :  128 - 0x80
    "10000000", -- 3729 - 0xe91  :  128 - 0x80
    "11000000", -- 3730 - 0xe92  :  192 - 0xc0
    "11000000", -- 3731 - 0xe93  :  192 - 0xc0
    "11100000", -- 3732 - 0xe94  :  224 - 0xe0
    "11111000", -- 3733 - 0xe95  :  248 - 0xf8
    "11111110", -- 3734 - 0xe96  :  254 - 0xfe
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111111", -- 3736 - 0xe98  :  255 - 0xff
    "01111111", -- 3737 - 0xe99  :  127 - 0x7f
    "00011111", -- 3738 - 0xe9a  :   31 - 0x1f
    "00000111", -- 3739 - 0xe9b  :    7 - 0x7
    "00000011", -- 3740 - 0xe9c  :    3 - 0x3
    "00000011", -- 3741 - 0xe9d  :    3 - 0x3
    "00000001", -- 3742 - 0xe9e  :    1 - 0x1
    "10000001", -- 3743 - 0xe9f  :  129 - 0x81
    "10000000", -- 3744 - 0xea0  :  128 - 0x80
    "10000000", -- 3745 - 0xea1  :  128 - 0x80
    "10000000", -- 3746 - 0xea2  :  128 - 0x80
    "11000000", -- 3747 - 0xea3  :  192 - 0xc0
    "11000000", -- 3748 - 0xea4  :  192 - 0xc0
    "11100000", -- 3749 - 0xea5  :  224 - 0xe0
    "11100000", -- 3750 - 0xea6  :  224 - 0xe0
    "11110000", -- 3751 - 0xea7  :  240 - 0xf0
    "00000001", -- 3752 - 0xea8  :    1 - 0x1
    "00000001", -- 3753 - 0xea9  :    1 - 0x1
    "00000001", -- 3754 - 0xeaa  :    1 - 0x1
    "00000011", -- 3755 - 0xeab  :    3 - 0x3
    "00000011", -- 3756 - 0xeac  :    3 - 0x3
    "00000111", -- 3757 - 0xead  :    7 - 0x7
    "00000111", -- 3758 - 0xeae  :    7 - 0x7
    "00001111", -- 3759 - 0xeaf  :   15 - 0xf
    "11111111", -- 3760 - 0xeb0  :  255 - 0xff
    "11111111", -- 3761 - 0xeb1  :  255 - 0xff
    "11111111", -- 3762 - 0xeb2  :  255 - 0xff
    "11111111", -- 3763 - 0xeb3  :  255 - 0xff
    "11111111", -- 3764 - 0xeb4  :  255 - 0xff
    "11111111", -- 3765 - 0xeb5  :  255 - 0xff
    "11111111", -- 3766 - 0xeb6  :  255 - 0xff
    "11111111", -- 3767 - 0xeb7  :  255 - 0xff
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "11111111", -- 3772 - 0xebc  :  255 - 0xff
    "11111111", -- 3773 - 0xebd  :  255 - 0xff
    "11111111", -- 3774 - 0xebe  :  255 - 0xff
    "11111111", -- 3775 - 0xebf  :  255 - 0xff
    "10000001", -- 3776 - 0xec0  :  129 - 0x81
    "10000001", -- 3777 - 0xec1  :  129 - 0x81
    "10000001", -- 3778 - 0xec2  :  129 - 0x81
    "10000001", -- 3779 - 0xec3  :  129 - 0x81
    "10000001", -- 3780 - 0xec4  :  129 - 0x81
    "10000001", -- 3781 - 0xec5  :  129 - 0x81
    "10000001", -- 3782 - 0xec6  :  129 - 0x81
    "10000001", -- 3783 - 0xec7  :  129 - 0x81
    "00000001", -- 3784 - 0xec8  :    1 - 0x1
    "00000001", -- 3785 - 0xec9  :    1 - 0x1
    "00000001", -- 3786 - 0xeca  :    1 - 0x1
    "00000011", -- 3787 - 0xecb  :    3 - 0x3
    "00000011", -- 3788 - 0xecc  :    3 - 0x3
    "00000111", -- 3789 - 0xecd  :    7 - 0x7
    "00000111", -- 3790 - 0xece  :    7 - 0x7
    "00001111", -- 3791 - 0xecf  :   15 - 0xf
    "00000001", -- 3792 - 0xed0  :    1 - 0x1
    "00000001", -- 3793 - 0xed1  :    1 - 0x1
    "00000001", -- 3794 - 0xed2  :    1 - 0x1
    "00000001", -- 3795 - 0xed3  :    1 - 0x1
    "00000001", -- 3796 - 0xed4  :    1 - 0x1
    "00000001", -- 3797 - 0xed5  :    1 - 0x1
    "00000001", -- 3798 - 0xed6  :    1 - 0x1
    "00000001", -- 3799 - 0xed7  :    1 - 0x1
    "10000001", -- 3800 - 0xed8  :  129 - 0x81
    "10000001", -- 3801 - 0xed9  :  129 - 0x81
    "10000001", -- 3802 - 0xeda  :  129 - 0x81
    "10000001", -- 3803 - 0xedb  :  129 - 0x81
    "10000001", -- 3804 - 0xedc  :  129 - 0x81
    "10000001", -- 3805 - 0xedd  :  129 - 0x81
    "10000001", -- 3806 - 0xede  :  129 - 0x81
    "10000001", -- 3807 - 0xedf  :  129 - 0x81
    "11111111", -- 3808 - 0xee0  :  255 - 0xff
    "00000011", -- 3809 - 0xee1  :    3 - 0x3
    "00000011", -- 3810 - 0xee2  :    3 - 0x3
    "00000011", -- 3811 - 0xee3  :    3 - 0x3
    "00000011", -- 3812 - 0xee4  :    3 - 0x3
    "00000011", -- 3813 - 0xee5  :    3 - 0x3
    "00000011", -- 3814 - 0xee6  :    3 - 0x3
    "11111111", -- 3815 - 0xee7  :  255 - 0xff
    "11111111", -- 3816 - 0xee8  :  255 - 0xff
    "11111111", -- 3817 - 0xee9  :  255 - 0xff
    "11111111", -- 3818 - 0xeea  :  255 - 0xff
    "11111111", -- 3819 - 0xeeb  :  255 - 0xff
    "11111111", -- 3820 - 0xeec  :  255 - 0xff
    "11111111", -- 3821 - 0xeed  :  255 - 0xff
    "11111111", -- 3822 - 0xeee  :  255 - 0xff
    "11111111", -- 3823 - 0xeef  :  255 - 0xff
    "10000000", -- 3824 - 0xef0  :  128 - 0x80
    "10000000", -- 3825 - 0xef1  :  128 - 0x80
    "10000000", -- 3826 - 0xef2  :  128 - 0x80
    "10000000", -- 3827 - 0xef3  :  128 - 0x80
    "10000000", -- 3828 - 0xef4  :  128 - 0x80
    "10000000", -- 3829 - 0xef5  :  128 - 0x80
    "10000000", -- 3830 - 0xef6  :  128 - 0x80
    "10000000", -- 3831 - 0xef7  :  128 - 0x80
    "00000001", -- 3832 - 0xef8  :    1 - 0x1
    "00000001", -- 3833 - 0xef9  :    1 - 0x1
    "00000001", -- 3834 - 0xefa  :    1 - 0x1
    "00000011", -- 3835 - 0xefb  :    3 - 0x3
    "00000111", -- 3836 - 0xefc  :    7 - 0x7
    "00000011", -- 3837 - 0xefd  :    3 - 0x3
    "00000001", -- 3838 - 0xefe  :    1 - 0x1
    "00000001", -- 3839 - 0xeff  :    1 - 0x1
    "10000001", -- 3840 - 0xf00  :  129 - 0x81
    "10000001", -- 3841 - 0xf01  :  129 - 0x81
    "10000001", -- 3842 - 0xf02  :  129 - 0x81
    "10000001", -- 3843 - 0xf03  :  129 - 0x81
    "10000001", -- 3844 - 0xf04  :  129 - 0x81
    "10000001", -- 3845 - 0xf05  :  129 - 0x81
    "10000001", -- 3846 - 0xf06  :  129 - 0x81
    "10000001", -- 3847 - 0xf07  :  129 - 0x81
    "11111111", -- 3848 - 0xf08  :  255 - 0xff
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "11111111", -- 3850 - 0xf0a  :  255 - 0xff
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "11111111", -- 3856 - 0xf10  :  255 - 0xff
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "11111111", -- 3860 - 0xf14  :  255 - 0xff
    "11111111", -- 3861 - 0xf15  :  255 - 0xff
    "11111111", -- 3862 - 0xf16  :  255 - 0xff
    "11111111", -- 3863 - 0xf17  :  255 - 0xff
    "10000001", -- 3864 - 0xf18  :  129 - 0x81
    "10000001", -- 3865 - 0xf19  :  129 - 0x81
    "10000001", -- 3866 - 0xf1a  :  129 - 0x81
    "10000001", -- 3867 - 0xf1b  :  129 - 0x81
    "10000001", -- 3868 - 0xf1c  :  129 - 0x81
    "10000001", -- 3869 - 0xf1d  :  129 - 0x81
    "10000001", -- 3870 - 0xf1e  :  129 - 0x81
    "10000001", -- 3871 - 0xf1f  :  129 - 0x81
    "10000000", -- 3872 - 0xf20  :  128 - 0x80
    "10000000", -- 3873 - 0xf21  :  128 - 0x80
    "11000000", -- 3874 - 0xf22  :  192 - 0xc0
    "11000000", -- 3875 - 0xf23  :  192 - 0xc0
    "11100000", -- 3876 - 0xf24  :  224 - 0xe0
    "11111000", -- 3877 - 0xf25  :  248 - 0xf8
    "11111110", -- 3878 - 0xf26  :  254 - 0xfe
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff
    "01111111", -- 3881 - 0xf29  :  127 - 0x7f
    "00011111", -- 3882 - 0xf2a  :   31 - 0x1f
    "00000111", -- 3883 - 0xf2b  :    7 - 0x7
    "00000011", -- 3884 - 0xf2c  :    3 - 0x3
    "00000011", -- 3885 - 0xf2d  :    3 - 0x3
    "00000001", -- 3886 - 0xf2e  :    1 - 0x1
    "10000001", -- 3887 - 0xf2f  :  129 - 0x81
    "10000001", -- 3888 - 0xf30  :  129 - 0x81
    "10000001", -- 3889 - 0xf31  :  129 - 0x81
    "10000001", -- 3890 - 0xf32  :  129 - 0x81
    "10000001", -- 3891 - 0xf33  :  129 - 0x81
    "10000001", -- 3892 - 0xf34  :  129 - 0x81
    "10000001", -- 3893 - 0xf35  :  129 - 0x81
    "10000001", -- 3894 - 0xf36  :  129 - 0x81
    "10000001", -- 3895 - 0xf37  :  129 - 0x81
    "10000001", -- 3896 - 0xf38  :  129 - 0x81
    "10000001", -- 3897 - 0xf39  :  129 - 0x81
    "10000001", -- 3898 - 0xf3a  :  129 - 0x81
    "10000001", -- 3899 - 0xf3b  :  129 - 0x81
    "10000001", -- 3900 - 0xf3c  :  129 - 0x81
    "10000001", -- 3901 - 0xf3d  :  129 - 0x81
    "10000001", -- 3902 - 0xf3e  :  129 - 0x81
    "10000001", -- 3903 - 0xf3f  :  129 - 0x81
    "01111110", -- 3904 - 0xf40  :  126 - 0x7e
    "00111100", -- 3905 - 0xf41  :   60 - 0x3c
    "00111100", -- 3906 - 0xf42  :   60 - 0x3c
    "00011000", -- 3907 - 0xf43  :   24 - 0x18
    "00011000", -- 3908 - 0xf44  :   24 - 0x18
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "11110010", -- 3912 - 0xf48  :  242 - 0xf2
    "11111110", -- 3913 - 0xf49  :  254 - 0xfe
    "11111110", -- 3914 - 0xf4a  :  254 - 0xfe
    "11111111", -- 3915 - 0xf4b  :  255 - 0xff
    "11111111", -- 3916 - 0xf4c  :  255 - 0xff
    "11101111", -- 3917 - 0xf4d  :  239 - 0xef
    "11110111", -- 3918 - 0xf4e  :  247 - 0xf7
    "11111000", -- 3919 - 0xf4f  :  248 - 0xf8
    "10111111", -- 3920 - 0xf50  :  191 - 0xbf
    "10111110", -- 3921 - 0xf51  :  190 - 0xbe
    "10111101", -- 3922 - 0xf52  :  189 - 0xbd
    "01111011", -- 3923 - 0xf53  :  123 - 0x7b
    "01111011", -- 3924 - 0xf54  :  123 - 0x7b
    "00000111", -- 3925 - 0xf55  :    7 - 0x7
    "11110011", -- 3926 - 0xf56  :  243 - 0xf3
    "11111101", -- 3927 - 0xf57  :  253 - 0xfd
    "11111111", -- 3928 - 0xf58  :  255 - 0xff
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "01100111", -- 3931 - 0xf5b  :  103 - 0x67
    "01011001", -- 3932 - 0xf5c  :   89 - 0x59
    "10011110", -- 3933 - 0xf5d  :  158 - 0x9e
    "10111111", -- 3934 - 0xf5e  :  191 - 0xbf
    "10111111", -- 3935 - 0xf5f  :  191 - 0xbf
    "00100000", -- 3936 - 0xf60  :   32 - 0x20
    "11100110", -- 3937 - 0xf61  :  230 - 0xe6
    "01010100", -- 3938 - 0xf62  :   84 - 0x54
    "00100110", -- 3939 - 0xf63  :   38 - 0x26
    "00100001", -- 3940 - 0xf64  :   33 - 0x21
    "00000110", -- 3941 - 0xf65  :    6 - 0x6
    "01010100", -- 3942 - 0xf66  :   84 - 0x54
    "00100110", -- 3943 - 0xf67  :   38 - 0x26
    "00100000", -- 3944 - 0xf68  :   32 - 0x20
    "10011010", -- 3945 - 0xf69  :  154 - 0x9a
    "00000001", -- 3946 - 0xf6a  :    1 - 0x1
    "01001001", -- 3947 - 0xf6b  :   73 - 0x49
    "00100000", -- 3948 - 0xf6c  :   32 - 0x20
    "10100101", -- 3949 - 0xf6d  :  165 - 0xa5
    "11001001", -- 3950 - 0xf6e  :  201 - 0xc9
    "01000110", -- 3951 - 0xf6f  :   70 - 0x46
    "11010001", -- 3952 - 0xf70  :  209 - 0xd1
    "11011000", -- 3953 - 0xf71  :  216 - 0xd8
    "11011000", -- 3954 - 0xf72  :  216 - 0xd8
    "11011110", -- 3955 - 0xf73  :  222 - 0xde
    "11010001", -- 3956 - 0xf74  :  209 - 0xd1
    "11010000", -- 3957 - 0xf75  :  208 - 0xd0
    "11011010", -- 3958 - 0xf76  :  218 - 0xda
    "11011110", -- 3959 - 0xf77  :  222 - 0xde
    "11011011", -- 3960 - 0xf78  :  219 - 0xdb
    "11011001", -- 3961 - 0xf79  :  217 - 0xd9
    "11011011", -- 3962 - 0xf7a  :  219 - 0xdb
    "11011100", -- 3963 - 0xf7b  :  220 - 0xdc
    "11011011", -- 3964 - 0xf7c  :  219 - 0xdb
    "11011111", -- 3965 - 0xf7d  :  223 - 0xdf
    "00100000", -- 3966 - 0xf7e  :   32 - 0x20
    "11100110", -- 3967 - 0xf7f  :  230 - 0xe6
    "11011010", -- 3968 - 0xf80  :  218 - 0xda
    "11011011", -- 3969 - 0xf81  :  219 - 0xdb
    "11100000", -- 3970 - 0xf82  :  224 - 0xe0
    "00100001", -- 3971 - 0xf83  :   33 - 0x21
    "00000110", -- 3972 - 0xf84  :    6 - 0x6
    "00001010", -- 3973 - 0xf85  :   10 - 0xa
    "11010110", -- 3974 - 0xf86  :  214 - 0xd6
    "11010111", -- 3975 - 0xf87  :  215 - 0xd7
    "00100001", -- 3976 - 0xf88  :   33 - 0x21
    "00100110", -- 3977 - 0xf89  :   38 - 0x26
    "00010100", -- 3978 - 0xf8a  :   20 - 0x14
    "11010000", -- 3979 - 0xf8b  :  208 - 0xd0
    "11101000", -- 3980 - 0xf8c  :  232 - 0xe8
    "11010001", -- 3981 - 0xf8d  :  209 - 0xd1
    "11010000", -- 3982 - 0xf8e  :  208 - 0xd0
    "11010001", -- 3983 - 0xf8f  :  209 - 0xd1
    "11011110", -- 3984 - 0xf90  :  222 - 0xde
    "11010001", -- 3985 - 0xf91  :  209 - 0xd1
    "11010000", -- 3986 - 0xf92  :  208 - 0xd0
    "11010001", -- 3987 - 0xf93  :  209 - 0xd1
    "11010000", -- 3988 - 0xf94  :  208 - 0xd0
    "11010001", -- 3989 - 0xf95  :  209 - 0xd1
    "00100110", -- 3990 - 0xf96  :   38 - 0x26
    "00100001", -- 3991 - 0xf97  :   33 - 0x21
    "01000010", -- 3992 - 0xf98  :   66 - 0x42
    "11011011", -- 3993 - 0xf99  :  219 - 0xdb
    "11011011", -- 3994 - 0xf9a  :  219 - 0xdb
    "01000010", -- 3995 - 0xf9b  :   66 - 0x42
    "00100110", -- 3996 - 0xf9c  :   38 - 0x26
    "11011011", -- 3997 - 0xf9d  :  219 - 0xdb
    "01000010", -- 3998 - 0xf9e  :   66 - 0x42
    "11011011", -- 3999 - 0xf9f  :  219 - 0xdb
    "01000110", -- 4000 - 0xfa0  :   70 - 0x46
    "11011011", -- 4001 - 0xfa1  :  219 - 0xdb
    "00100001", -- 4002 - 0xfa2  :   33 - 0x21
    "01101100", -- 4003 - 0xfa3  :  108 - 0x6c
    "00001110", -- 4004 - 0xfa4  :   14 - 0xe
    "11011111", -- 4005 - 0xfa5  :  223 - 0xdf
    "11011011", -- 4006 - 0xfa6  :  219 - 0xdb
    "11011011", -- 4007 - 0xfa7  :  219 - 0xdb
    "11100100", -- 4008 - 0xfa8  :  228 - 0xe4
    "11100101", -- 4009 - 0xfa9  :  229 - 0xe5
    "00100110", -- 4010 - 0xfaa  :   38 - 0x26
    "00100001", -- 4011 - 0xfab  :   33 - 0x21
    "10000110", -- 4012 - 0xfac  :  134 - 0x86
    "00010100", -- 4013 - 0xfad  :   20 - 0x14
    "11011011", -- 4014 - 0xfae  :  219 - 0xdb
    "11011011", -- 4015 - 0xfaf  :  219 - 0xdb
    "00100110", -- 4016 - 0xfb0  :   38 - 0x26
    "11011011", -- 4017 - 0xfb1  :  219 - 0xdb
    "11100011", -- 4018 - 0xfb2  :  227 - 0xe3
    "11011011", -- 4019 - 0xfb3  :  219 - 0xdb
    "11100000", -- 4020 - 0xfb4  :  224 - 0xe0
    "11011011", -- 4021 - 0xfb5  :  219 - 0xdb
    "11011011", -- 4022 - 0xfb6  :  219 - 0xdb
    "11100110", -- 4023 - 0xfb7  :  230 - 0xe6
    "11011011", -- 4024 - 0xfb8  :  219 - 0xdb
    "01000010", -- 4025 - 0xfb9  :   66 - 0x42
    "11011011", -- 4026 - 0xfba  :  219 - 0xdb
    "11011011", -- 4027 - 0xfbb  :  219 - 0xdb
    "11011011", -- 4028 - 0xfbc  :  219 - 0xdb
    "11010100", -- 4029 - 0xfbd  :  212 - 0xd4
    "11011001", -- 4030 - 0xfbe  :  217 - 0xd9
    "00100110", -- 4031 - 0xfbf  :   38 - 0x26
    "11100111", -- 4032 - 0xfc0  :  231 - 0xe7
    "00100001", -- 4033 - 0xfc1  :   33 - 0x21
    "11000101", -- 4034 - 0xfc2  :  197 - 0xc5
    "00010110", -- 4035 - 0xfc3  :   22 - 0x16
    "01011111", -- 4036 - 0xfc4  :   95 - 0x5f
    "10010101", -- 4037 - 0xfc5  :  149 - 0x95
    "10010101", -- 4038 - 0xfc6  :  149 - 0x95
    "10010101", -- 4039 - 0xfc7  :  149 - 0x95
    "10010101", -- 4040 - 0xfc8  :  149 - 0x95
    "10010110", -- 4041 - 0xfc9  :  150 - 0x96
    "10010101", -- 4042 - 0xfca  :  149 - 0x95
    "10010101", -- 4043 - 0xfcb  :  149 - 0x95
    "10010111", -- 4044 - 0xfcc  :  151 - 0x97
    "10011000", -- 4045 - 0xfcd  :  152 - 0x98
    "10010111", -- 4046 - 0xfce  :  151 - 0x97
    "10011000", -- 4047 - 0xfcf  :  152 - 0x98
    "00001000", -- 4048 - 0xfd0  :    8 - 0x8
    "00000101", -- 4049 - 0xfd1  :    5 - 0x5
    "00100100", -- 4050 - 0xfd2  :   36 - 0x24
    "00010111", -- 4051 - 0xfd3  :   23 - 0x17
    "00010010", -- 4052 - 0xfd4  :   18 - 0x12
    "00010111", -- 4053 - 0xfd5  :   23 - 0x17
    "00011101", -- 4054 - 0xfd6  :   29 - 0x1d
    "00001110", -- 4055 - 0xfd7  :   14 - 0xe
    "00011001", -- 4056 - 0xfd8  :   25 - 0x19
    "00010101", -- 4057 - 0xfd9  :   21 - 0x15
    "00001010", -- 4058 - 0xfda  :   10 - 0xa
    "00100010", -- 4059 - 0xfdb  :   34 - 0x22
    "00001110", -- 4060 - 0xfdc  :   14 - 0xe
    "00011011", -- 4061 - 0xfdd  :   27 - 0x1b
    "00100100", -- 4062 - 0xfde  :   36 - 0x24
    "00010000", -- 4063 - 0xfdf  :   16 - 0x10
    "00011001", -- 4064 - 0xfe0  :   25 - 0x19
    "00010101", -- 4065 - 0xfe1  :   21 - 0x15
    "00001010", -- 4066 - 0xfe2  :   10 - 0xa
    "00100010", -- 4067 - 0xfe3  :   34 - 0x22
    "00001110", -- 4068 - 0xfe4  :   14 - 0xe
    "00011011", -- 4069 - 0xfe5  :   27 - 0x1b
    "00100100", -- 4070 - 0xfe6  :   36 - 0x24
    "00010000", -- 4071 - 0xfe7  :   16 - 0x10
    "00011001", -- 4072 - 0xfe8  :   25 - 0x19
    "00101000", -- 4073 - 0xfe9  :   40 - 0x28
    "00100010", -- 4074 - 0xfea  :   34 - 0x22
    "11110110", -- 4075 - 0xfeb  :  246 - 0xf6
    "00000001", -- 4076 - 0xfec  :    1 - 0x1
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00100011", -- 4078 - 0xfee  :   35 - 0x23
    "11001001", -- 4079 - 0xfef  :  201 - 0xc9
    "10101010", -- 4080 - 0xff0  :  170 - 0xaa
    "00100011", -- 4081 - 0xff1  :   35 - 0x23
    "11101010", -- 4082 - 0xff2  :  234 - 0xea
    "00000100", -- 4083 - 0xff3  :    4 - 0x4
    "10011001", -- 4084 - 0xff4  :  153 - 0x99
    "10101010", -- 4085 - 0xff5  :  170 - 0xaa
    "10101010", -- 4086 - 0xff6  :  170 - 0xaa
    "10101010", -- 4087 - 0xff7  :  170 - 0xaa
    "11111111", -- 4088 - 0xff8  :  255 - 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111" -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= nametable_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
