--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_color1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_color1;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_color1 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000011", --    2 -  0x2  :    3 - 0x3
    "00000001", --    3 -  0x3  :    1 - 0x1
    "00000001", --    4 -  0x4  :    1 - 0x1
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000011", --    6 -  0x6  :    3 - 0x3
    "00000001", --    7 -  0x7  :    1 - 0x1
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00111000", --   10 -  0xa  :   56 - 0x38
    "10110100", --   11 -  0xb  :  180 - 0xb4
    "10101000", --   12 -  0xc  :  168 - 0xa8
    "11010100", --   13 -  0xd  :  212 - 0xd4
    "01110100", --   14 -  0xe  :  116 - 0x74
    "01111110", --   15 -  0xf  :  126 - 0x7e
    "00111000", --   16 - 0x10  :   56 - 0x38 -- Sprite 0x2
    "01111000", --   17 - 0x11  :  120 - 0x78
    "01111100", --   18 - 0x12  :  124 - 0x7c
    "01111110", --   19 - 0x13  :  126 - 0x7e
    "01111110", --   20 - 0x14  :  126 - 0x7e
    "01111110", --   21 - 0x15  :  126 - 0x7e
    "00111110", --   22 - 0x16  :   62 - 0x3e
    "00011110", --   23 - 0x17  :   30 - 0x1e
    "11110110", --   24 - 0x18  :  246 - 0xf6 -- Sprite 0x3
    "11110000", --   25 - 0x19  :  240 - 0xf0
    "00111000", --   26 - 0x1a  :   56 - 0x38
    "11010000", --   27 - 0x1b  :  208 - 0xd0
    "11100000", --   28 - 0x1c  :  224 - 0xe0
    "01110000", --   29 - 0x1d  :  112 - 0x70
    "10111000", --   30 - 0x1e  :  184 - 0xb8
    "01000000", --   31 - 0x1f  :   64 - 0x40
    "00011100", --   32 - 0x20  :   28 - 0x1c -- Sprite 0x4
    "00011100", --   33 - 0x21  :   28 - 0x1c
    "00011110", --   34 - 0x22  :   30 - 0x1e
    "00011111", --   35 - 0x23  :   31 - 0x1f
    "00001100", --   36 - 0x24  :   12 - 0xc
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "10101000", --   40 - 0x28  :  168 - 0xa8 -- Sprite 0x5
    "01010000", --   41 - 0x29  :   80 - 0x50
    "10101000", --   42 - 0x2a  :  168 - 0xa8
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "01100000", --   44 - 0x2c  :   96 - 0x60
    "01100000", --   45 - 0x2d  :   96 - 0x60
    "01110000", --   46 - 0x2e  :  112 - 0x70
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00011100", --   48 - 0x30  :   28 - 0x1c -- Sprite 0x6
    "00011100", --   49 - 0x31  :   28 - 0x1c
    "00011110", --   50 - 0x32  :   30 - 0x1e
    "00011111", --   51 - 0x33  :   31 - 0x1f
    "00001100", --   52 - 0x34  :   12 - 0xc
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000001", --   54 - 0x36  :    1 - 0x1
    "00000000", --   55 - 0x37  :    0 - 0x0
    "10101000", --   56 - 0x38  :  168 - 0xa8 -- Sprite 0x7
    "01010000", --   57 - 0x39  :   80 - 0x50
    "10101000", --   58 - 0x3a  :  168 - 0xa8
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "01011000", --   60 - 0x3c  :   88 - 0x58
    "11011000", --   61 - 0x3d  :  216 - 0xd8
    "10001100", --   62 - 0x3e  :  140 - 0x8c
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00011100", --   64 - 0x40  :   28 - 0x1c -- Sprite 0x8
    "00011100", --   65 - 0x41  :   28 - 0x1c
    "00011110", --   66 - 0x42  :   30 - 0x1e
    "00011111", --   67 - 0x43  :   31 - 0x1f
    "00001100", --   68 - 0x44  :   12 - 0xc
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "10101000", --   72 - 0x48  :  168 - 0xa8 -- Sprite 0x9
    "01010100", --   73 - 0x49  :   84 - 0x54
    "10101000", --   74 - 0x4a  :  168 - 0xa8
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "01101110", --   76 - 0x4c  :  110 - 0x6e
    "11000000", --   77 - 0x4d  :  192 - 0xc0
    "10000000", --   78 - 0x4e  :  128 - 0x80
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00011100", --   80 - 0x50  :   28 - 0x1c -- Sprite 0xa
    "00011100", --   81 - 0x51  :   28 - 0x1c
    "00011110", --   82 - 0x52  :   30 - 0x1e
    "00011111", --   83 - 0x53  :   31 - 0x1f
    "00001100", --   84 - 0x54  :   12 - 0xc
    "00000001", --   85 - 0x55  :    1 - 0x1
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "10101000", --   88 - 0x58  :  168 - 0xa8 -- Sprite 0xb
    "01010100", --   89 - 0x59  :   84 - 0x54
    "10101000", --   90 - 0x5a  :  168 - 0xa8
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "11011000", --   92 - 0x5c  :  216 - 0xd8
    "11011100", --   93 - 0x5d  :  220 - 0xdc
    "00001100", --   94 - 0x5e  :   12 - 0xc
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "11110110", --   96 - 0x60  :  246 - 0xf6 -- Sprite 0xc
    "11110000", --   97 - 0x61  :  240 - 0xf0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "11111100", --   99 - 0x63  :  252 - 0xfc
    "11111000", --  100 - 0x64  :  248 - 0xf8
    "00000000", --  101 - 0x65  :    0 - 0x0
    "10101000", --  102 - 0x66  :  168 - 0xa8
    "01010100", --  103 - 0x67  :   84 - 0x54
    "00111000", --  104 - 0x68  :   56 - 0x38 -- Sprite 0xd
    "01111000", --  105 - 0x69  :  120 - 0x78
    "01111100", --  106 - 0x6a  :  124 - 0x7c
    "01111101", --  107 - 0x6b  :  125 - 0x7d
    "01111101", --  108 - 0x6c  :  125 - 0x7d
    "01111011", --  109 - 0x6d  :  123 - 0x7b
    "00111011", --  110 - 0x6e  :   59 - 0x3b
    "00011011", --  111 - 0x6f  :   27 - 0x1b
    "11110110", --  112 - 0x70  :  246 - 0xf6 -- Sprite 0xe
    "11110000", --  113 - 0x71  :  240 - 0xf0
    "01111000", --  114 - 0x72  :  120 - 0x78
    "01110000", --  115 - 0x73  :  112 - 0x70
    "10100000", --  116 - 0x74  :  160 - 0xa0
    "10010000", --  117 - 0x75  :  144 - 0x90
    "00101000", --  118 - 0x76  :   40 - 0x28
    "01010100", --  119 - 0x77  :   84 - 0x54
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000011", --  122 - 0x7a  :    3 - 0x3
    "00000001", --  123 - 0x7b  :    1 - 0x1
    "00000001", --  124 - 0x7c  :    1 - 0x1
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000011", --  126 - 0x7e  :    3 - 0x3
    "00000001", --  127 - 0x7f  :    1 - 0x1
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  129 - 0x81  :    3 - 0x3
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00001111", --  131 - 0x83  :   15 - 0xf
    "00001111", --  132 - 0x84  :   15 - 0xf
    "00011111", --  133 - 0x85  :   31 - 0x1f
    "00011111", --  134 - 0x86  :   31 - 0x1f
    "00011110", --  135 - 0x87  :   30 - 0x1e
    "00110110", --  136 - 0x88  :   54 - 0x36 -- Sprite 0x11
    "10110000", --  137 - 0x89  :  176 - 0xb0
    "10111000", --  138 - 0x8a  :  184 - 0xb8
    "10010000", --  139 - 0x8b  :  144 - 0x90
    "10100000", --  140 - 0x8c  :  160 - 0xa0
    "01110000", --  141 - 0x8d  :  112 - 0x70
    "00111000", --  142 - 0x8e  :   56 - 0x38
    "01000000", --  143 - 0x8f  :   64 - 0x40
    "00011100", --  144 - 0x90  :   28 - 0x1c -- Sprite 0x12
    "00011100", --  145 - 0x91  :   28 - 0x1c
    "00011110", --  146 - 0x92  :   30 - 0x1e
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00001100", --  148 - 0x94  :   12 - 0xc
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000011", --  155 - 0x9b  :    3 - 0x3
    "00000111", --  156 - 0x9c  :    7 - 0x7
    "00001111", --  157 - 0x9d  :   15 - 0xf
    "00001111", --  158 - 0x9e  :   15 - 0xf
    "00011111", --  159 - 0x9f  :   31 - 0x1f
    "11110110", --  160 - 0xa0  :  246 - 0xf6 -- Sprite 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "11111000", --  162 - 0xa2  :  248 - 0xf8
    "11111110", --  163 - 0xa3  :  254 - 0xfe
    "11111110", --  164 - 0xa4  :  254 - 0xfe
    "11111110", --  165 - 0xa5  :  254 - 0xfe
    "11111000", --  166 - 0xa6  :  248 - 0xf8
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000011", --  168 - 0xa8  :    3 - 0x3 -- Sprite 0x15
    "00000011", --  169 - 0xa9  :    3 - 0x3
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000011", --  171 - 0xab  :    3 - 0x3
    "00000011", --  172 - 0xac  :    3 - 0x3
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00001111", --  174 - 0xae  :   15 - 0xf
    "00111111", --  175 - 0xaf  :   63 - 0x3f
    "11011000", --  176 - 0xb0  :  216 - 0xd8 -- Sprite 0x16
    "11000000", --  177 - 0xb1  :  192 - 0xc0
    "11100000", --  178 - 0xb2  :  224 - 0xe0
    "01000000", --  179 - 0xb3  :   64 - 0x40
    "10000000", --  180 - 0xb4  :  128 - 0x80
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "11100000", --  182 - 0xb6  :  224 - 0xe0
    "11111100", --  183 - 0xb7  :  252 - 0xfc
    "01111111", --  184 - 0xb8  :  127 - 0x7f -- Sprite 0x17
    "01111111", --  185 - 0xb9  :  127 - 0x7f
    "01111111", --  186 - 0xba  :  127 - 0x7f
    "01111100", --  187 - 0xbb  :  124 - 0x7c
    "00110000", --  188 - 0xbc  :   48 - 0x30
    "00000001", --  189 - 0xbd  :    1 - 0x1
    "00000001", --  190 - 0xbe  :    1 - 0x1
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "11111100", --  192 - 0xc0  :  252 - 0xfc -- Sprite 0x18
    "11111110", --  193 - 0xc1  :  254 - 0xfe
    "11111100", --  194 - 0xc2  :  252 - 0xfc
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "10000000", --  197 - 0xc5  :  128 - 0x80
    "11000000", --  198 - 0xc6  :  192 - 0xc0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000111", --  200 - 0xc8  :    7 - 0x7 -- Sprite 0x19
    "00000111", --  201 - 0xc9  :    7 - 0x7
    "00000001", --  202 - 0xca  :    1 - 0x1
    "00000110", --  203 - 0xcb  :    6 - 0x6
    "00000111", --  204 - 0xcc  :    7 - 0x7
    "00000110", --  205 - 0xcd  :    6 - 0x6
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00001111", --  207 - 0xcf  :   15 - 0xf
    "10110000", --  208 - 0xd0  :  176 - 0xb0 -- Sprite 0x1a
    "10000000", --  209 - 0xd1  :  128 - 0x80
    "11000000", --  210 - 0xd2  :  192 - 0xc0
    "10000000", --  211 - 0xd3  :  128 - 0x80
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "11100000", --  215 - 0xd7  :  224 - 0xe0
    "00111111", --  216 - 0xd8  :   63 - 0x3f -- Sprite 0x1b
    "00111111", --  217 - 0xd9  :   63 - 0x3f
    "01111111", --  218 - 0xda  :  127 - 0x7f
    "01111111", --  219 - 0xdb  :  127 - 0x7f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000011", --  222 - 0xde  :    3 - 0x3
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "11111111", --  224 - 0xe0  :  255 - 0xff -- Sprite 0x1c
    "11111111", --  225 - 0xe1  :  255 - 0xff
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111111", --  227 - 0xe3  :  255 - 0xff
    "11111111", --  228 - 0xe4  :  255 - 0xff
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "10000000", --  230 - 0xe6  :  128 - 0x80
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Sprite 0x1d
    "11000000", --  233 - 0xe9  :  192 - 0xc0
    "11000000", --  234 - 0xea  :  192 - 0xc0
    "11000000", --  235 - 0xeb  :  192 - 0xc0
    "10000000", --  236 - 0xec  :  128 - 0x80
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "11100000", --  240 - 0xf0  :  224 - 0xe0 -- Sprite 0x1e
    "10011100", --  241 - 0xf1  :  156 - 0x9c
    "00111000", --  242 - 0xf2  :   56 - 0x38
    "11100000", --  243 - 0xf3  :  224 - 0xe0
    "11001000", --  244 - 0xf4  :  200 - 0xc8
    "00010100", --  245 - 0xf5  :   20 - 0x14
    "10101000", --  246 - 0xf6  :  168 - 0xa8
    "01010100", --  247 - 0xf7  :   84 - 0x54
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00111000", --  250 - 0xfa  :   56 - 0x38
    "10110100", --  251 - 0xfb  :  180 - 0xb4
    "10101000", --  252 - 0xfc  :  168 - 0xa8
    "11010100", --  253 - 0xfd  :  212 - 0xd4
    "01110100", --  254 - 0xfe  :  116 - 0x74
    "00011110", --  255 - 0xff  :   30 - 0x1e
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00001100", --  258 - 0x102  :   12 - 0xc
    "00000111", --  259 - 0x103  :    7 - 0x7
    "00001111", --  260 - 0x104  :   15 - 0xf
    "00000111", --  261 - 0x105  :    7 - 0x7
    "00001111", --  262 - 0x106  :   15 - 0xf
    "00001111", --  263 - 0x107  :   15 - 0xf
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00110000", --  266 - 0x10a  :   48 - 0x30
    "11100000", --  267 - 0x10b  :  224 - 0xe0
    "11110000", --  268 - 0x10c  :  240 - 0xf0
    "11100000", --  269 - 0x10d  :  224 - 0xe0
    "11110000", --  270 - 0x10e  :  240 - 0xf0
    "11110000", --  271 - 0x10f  :  240 - 0xf0
    "00000111", --  272 - 0x110  :    7 - 0x7 -- Sprite 0x22
    "00000011", --  273 - 0x111  :    3 - 0x3
    "00011000", --  274 - 0x112  :   24 - 0x18
    "00010101", --  275 - 0x113  :   21 - 0x15
    "00000010", --  276 - 0x114  :    2 - 0x2
    "00000101", --  277 - 0x115  :    5 - 0x5
    "00000010", --  278 - 0x116  :    2 - 0x2
    "00000100", --  279 - 0x117  :    4 - 0x4
    "11100000", --  280 - 0x118  :  224 - 0xe0 -- Sprite 0x23
    "11000000", --  281 - 0x119  :  192 - 0xc0
    "00111100", --  282 - 0x11a  :   60 - 0x3c
    "01111100", --  283 - 0x11b  :  124 - 0x7c
    "01111100", --  284 - 0x11c  :  124 - 0x7c
    "01111100", --  285 - 0x11d  :  124 - 0x7c
    "11101100", --  286 - 0x11e  :  236 - 0xec
    "11100000", --  287 - 0x11f  :  224 - 0xe0
    "00000010", --  288 - 0x120  :    2 - 0x2 -- Sprite 0x24
    "00000101", --  289 - 0x121  :    5 - 0x5
    "00001011", --  290 - 0x122  :   11 - 0xb
    "00001011", --  291 - 0x123  :   11 - 0xb
    "00001101", --  292 - 0x124  :   13 - 0xd
    "00011000", --  293 - 0x125  :   24 - 0x18
    "00111000", --  294 - 0x126  :   56 - 0x38
    "00000000", --  295 - 0x127  :    0 - 0x0
    "11100000", --  296 - 0x128  :  224 - 0xe0 -- Sprite 0x25
    "11100000", --  297 - 0x129  :  224 - 0xe0
    "11100000", --  298 - 0x12a  :  224 - 0xe0
    "11010000", --  299 - 0x12b  :  208 - 0xd0
    "10111000", --  300 - 0x12c  :  184 - 0xb8
    "00111000", --  301 - 0x12d  :   56 - 0x38
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Sprite 0x27
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Sprite 0x29
    "00011111", --  329 - 0x149  :   31 - 0x1f
    "00011111", --  330 - 0x14a  :   31 - 0x1f
    "00011111", --  331 - 0x14b  :   31 - 0x1f
    "00001100", --  332 - 0x14c  :   12 - 0xc
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000001", --  334 - 0x14e  :    1 - 0x1
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00011111", --  336 - 0x150  :   31 - 0x1f -- Sprite 0x2a
    "00011111", --  337 - 0x151  :   31 - 0x1f
    "00011111", --  338 - 0x152  :   31 - 0x1f
    "00011111", --  339 - 0x153  :   31 - 0x1f
    "00001100", --  340 - 0x154  :   12 - 0xc
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Sprite 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Sprite 0x2d
    "01111110", --  361 - 0x169  :  126 - 0x7e
    "01000010", --  362 - 0x16a  :   66 - 0x42
    "01000010", --  363 - 0x16b  :   66 - 0x42
    "01000010", --  364 - 0x16c  :   66 - 0x42
    "01000010", --  365 - 0x16d  :   66 - 0x42
    "01111110", --  366 - 0x16e  :  126 - 0x7e
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "01100110", --  376 - 0x178  :  102 - 0x66 -- Sprite 0x2f
    "01100000", --  377 - 0x179  :   96 - 0x60
    "01101000", --  378 - 0x17a  :  104 - 0x68
    "11100000", --  379 - 0x17b  :  224 - 0xe0
    "11000000", --  380 - 0x17c  :  192 - 0xc0
    "00010000", --  381 - 0x17d  :   16 - 0x10
    "00101000", --  382 - 0x17e  :   40 - 0x28
    "01010000", --  383 - 0x17f  :   80 - 0x50
    "11110110", --  384 - 0x180  :  246 - 0xf6 -- Sprite 0x30
    "11110000", --  385 - 0x181  :  240 - 0xf0
    "00111000", --  386 - 0x182  :   56 - 0x38
    "11010000", --  387 - 0x183  :  208 - 0xd0
    "11000000", --  388 - 0x184  :  192 - 0xc0
    "11111000", --  389 - 0x185  :  248 - 0xf8
    "01111000", --  390 - 0x186  :  120 - 0x78
    "00000000", --  391 - 0x187  :    0 - 0x0
    "11110110", --  392 - 0x188  :  246 - 0xf6 -- Sprite 0x31
    "11110000", --  393 - 0x189  :  240 - 0xf0
    "00111000", --  394 - 0x18a  :   56 - 0x38
    "11010000", --  395 - 0x18b  :  208 - 0xd0
    "11000000", --  396 - 0x18c  :  192 - 0xc0
    "11100000", --  397 - 0x18d  :  224 - 0xe0
    "01111000", --  398 - 0x18e  :  120 - 0x78
    "00111000", --  399 - 0x18f  :   56 - 0x38
    "11110110", --  400 - 0x190  :  246 - 0xf6 -- Sprite 0x32
    "11110000", --  401 - 0x191  :  240 - 0xf0
    "00111000", --  402 - 0x192  :   56 - 0x38
    "11000000", --  403 - 0x193  :  192 - 0xc0
    "11011000", --  404 - 0x194  :  216 - 0xd8
    "11111000", --  405 - 0x195  :  248 - 0xf8
    "01100000", --  406 - 0x196  :   96 - 0x60
    "00010000", --  407 - 0x197  :   16 - 0x10
    "00011100", --  408 - 0x198  :   28 - 0x1c -- Sprite 0x33
    "00011100", --  409 - 0x199  :   28 - 0x1c
    "00011110", --  410 - 0x19a  :   30 - 0x1e
    "00011111", --  411 - 0x19b  :   31 - 0x1f
    "00001100", --  412 - 0x19c  :   12 - 0xc
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "10000000", --  416 - 0x1a0  :  128 - 0x80 -- Sprite 0x34
    "01010000", --  417 - 0x1a1  :   80 - 0x50
    "10101000", --  418 - 0x1a2  :  168 - 0xa8
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "01011000", --  420 - 0x1a4  :   88 - 0x58
    "11011000", --  421 - 0x1a5  :  216 - 0xd8
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00011100", --  424 - 0x1a8  :   28 - 0x1c -- Sprite 0x35
    "00011100", --  425 - 0x1a9  :   28 - 0x1c
    "00011110", --  426 - 0x1aa  :   30 - 0x1e
    "00011111", --  427 - 0x1ab  :   31 - 0x1f
    "00001100", --  428 - 0x1ac  :   12 - 0xc
    "00000001", --  429 - 0x1ad  :    1 - 0x1
    "00000001", --  430 - 0x1ae  :    1 - 0x1
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "10101000", --  432 - 0x1b0  :  168 - 0xa8 -- Sprite 0x36
    "01010000", --  433 - 0x1b1  :   80 - 0x50
    "10101000", --  434 - 0x1b2  :  168 - 0xa8
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "01011000", --  436 - 0x1b4  :   88 - 0x58
    "11001110", --  437 - 0x1b5  :  206 - 0xce
    "10000110", --  438 - 0x1b6  :  134 - 0x86
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "10101000", --  440 - 0x1b8  :  168 - 0xa8 -- Sprite 0x37
    "01010000", --  441 - 0x1b9  :   80 - 0x50
    "10101000", --  442 - 0x1ba  :  168 - 0xa8
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "01011000", --  444 - 0x1bc  :   88 - 0x58
    "11011000", --  445 - 0x1bd  :  216 - 0xd8
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00111100", --  512 - 0x200  :   60 - 0x3c -- Sprite 0x40
    "01111100", --  513 - 0x201  :  124 - 0x7c
    "11100110", --  514 - 0x202  :  230 - 0xe6
    "11101110", --  515 - 0x203  :  238 - 0xee
    "11110110", --  516 - 0x204  :  246 - 0xf6
    "11100110", --  517 - 0x205  :  230 - 0xe6
    "00111100", --  518 - 0x206  :   60 - 0x3c
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00111000", --  520 - 0x208  :   56 - 0x38 -- Sprite 0x41
    "01111000", --  521 - 0x209  :  120 - 0x78
    "00111000", --  522 - 0x20a  :   56 - 0x38
    "00111000", --  523 - 0x20b  :   56 - 0x38
    "00111000", --  524 - 0x20c  :   56 - 0x38
    "00111000", --  525 - 0x20d  :   56 - 0x38
    "00111000", --  526 - 0x20e  :   56 - 0x38
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01111100", --  528 - 0x210  :  124 - 0x7c -- Sprite 0x42
    "11111110", --  529 - 0x211  :  254 - 0xfe
    "11100110", --  530 - 0x212  :  230 - 0xe6
    "00011110", --  531 - 0x213  :   30 - 0x1e
    "01111100", --  532 - 0x214  :  124 - 0x7c
    "11100000", --  533 - 0x215  :  224 - 0xe0
    "11111110", --  534 - 0x216  :  254 - 0xfe
    "00000000", --  535 - 0x217  :    0 - 0x0
    "01111100", --  536 - 0x218  :  124 - 0x7c -- Sprite 0x43
    "11111100", --  537 - 0x219  :  252 - 0xfc
    "11100110", --  538 - 0x21a  :  230 - 0xe6
    "00011100", --  539 - 0x21b  :   28 - 0x1c
    "01100110", --  540 - 0x21c  :  102 - 0x66
    "11101110", --  541 - 0x21d  :  238 - 0xee
    "11111100", --  542 - 0x21e  :  252 - 0xfc
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00001100", --  544 - 0x220  :   12 - 0xc -- Sprite 0x44
    "00011100", --  545 - 0x221  :   28 - 0x1c
    "00111100", --  546 - 0x222  :   60 - 0x3c
    "01111100", --  547 - 0x223  :  124 - 0x7c
    "11101100", --  548 - 0x224  :  236 - 0xec
    "11111110", --  549 - 0x225  :  254 - 0xfe
    "00001100", --  550 - 0x226  :   12 - 0xc
    "00000000", --  551 - 0x227  :    0 - 0x0
    "11111110", --  552 - 0x228  :  254 - 0xfe -- Sprite 0x45
    "11111110", --  553 - 0x229  :  254 - 0xfe
    "11100000", --  554 - 0x22a  :  224 - 0xe0
    "11111110", --  555 - 0x22b  :  254 - 0xfe
    "00000110", --  556 - 0x22c  :    6 - 0x6
    "11101110", --  557 - 0x22d  :  238 - 0xee
    "11111100", --  558 - 0x22e  :  252 - 0xfc
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00111100", --  560 - 0x230  :   60 - 0x3c -- Sprite 0x46
    "01111100", --  561 - 0x231  :  124 - 0x7c
    "11100000", --  562 - 0x232  :  224 - 0xe0
    "11111110", --  563 - 0x233  :  254 - 0xfe
    "11100110", --  564 - 0x234  :  230 - 0xe6
    "11101110", --  565 - 0x235  :  238 - 0xee
    "00111100", --  566 - 0x236  :   60 - 0x3c
    "00000000", --  567 - 0x237  :    0 - 0x0
    "11111110", --  568 - 0x238  :  254 - 0xfe -- Sprite 0x47
    "11111100", --  569 - 0x239  :  252 - 0xfc
    "00001100", --  570 - 0x23a  :   12 - 0xc
    "00111000", --  571 - 0x23b  :   56 - 0x38
    "00111000", --  572 - 0x23c  :   56 - 0x38
    "01110000", --  573 - 0x23d  :  112 - 0x70
    "01110000", --  574 - 0x23e  :  112 - 0x70
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00111110", --  576 - 0x240  :   62 - 0x3e -- Sprite 0x48
    "01111100", --  577 - 0x241  :  124 - 0x7c
    "11100110", --  578 - 0x242  :  230 - 0xe6
    "10111100", --  579 - 0x243  :  188 - 0xbc
    "11100110", --  580 - 0x244  :  230 - 0xe6
    "11101110", --  581 - 0x245  :  238 - 0xee
    "00111100", --  582 - 0x246  :   60 - 0x3c
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00111100", --  584 - 0x248  :   60 - 0x3c -- Sprite 0x49
    "01111100", --  585 - 0x249  :  124 - 0x7c
    "11100110", --  586 - 0x24a  :  230 - 0xe6
    "11101110", --  587 - 0x24b  :  238 - 0xee
    "11111110", --  588 - 0x24c  :  254 - 0xfe
    "10000110", --  589 - 0x24d  :  134 - 0x86
    "01111100", --  590 - 0x24e  :  124 - 0x7c
    "01000000", --  591 - 0x24f  :   64 - 0x40
    "11101110", --  592 - 0x250  :  238 - 0xee -- Sprite 0x4a
    "11101110", --  593 - 0x251  :  238 - 0xee
    "11101110", --  594 - 0x252  :  238 - 0xee
    "11101110", --  595 - 0x253  :  238 - 0xee
    "11101110", --  596 - 0x254  :  238 - 0xee
    "11101110", --  597 - 0x255  :  238 - 0xee
    "11101110", --  598 - 0x256  :  238 - 0xee
    "10001000", --  599 - 0x257  :  136 - 0x88
    "11100000", --  600 - 0x258  :  224 - 0xe0 -- Sprite 0x4b
    "11100000", --  601 - 0x259  :  224 - 0xe0
    "11100000", --  602 - 0x25a  :  224 - 0xe0
    "11100000", --  603 - 0x25b  :  224 - 0xe0
    "11100000", --  604 - 0x25c  :  224 - 0xe0
    "11100000", --  605 - 0x25d  :  224 - 0xe0
    "11100000", --  606 - 0x25e  :  224 - 0xe0
    "10000000", --  607 - 0x25f  :  128 - 0x80
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x4c
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "01111111", --  610 - 0x262  :  127 - 0x7f
    "01111111", --  611 - 0x263  :  127 - 0x7f
    "01111111", --  612 - 0x264  :  127 - 0x7f
    "01111111", --  613 - 0x265  :  127 - 0x7f
    "01111111", --  614 - 0x266  :  127 - 0x7f
    "01111111", --  615 - 0x267  :  127 - 0x7f
    "01111111", --  616 - 0x268  :  127 - 0x7f -- Sprite 0x4d
    "01111111", --  617 - 0x269  :  127 - 0x7f
    "01111111", --  618 - 0x26a  :  127 - 0x7f
    "01111111", --  619 - 0x26b  :  127 - 0x7f
    "01111111", --  620 - 0x26c  :  127 - 0x7f
    "01111111", --  621 - 0x26d  :  127 - 0x7f
    "01111111", --  622 - 0x26e  :  127 - 0x7f
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x4e
    "11111110", --  625 - 0x271  :  254 - 0xfe
    "11111110", --  626 - 0x272  :  254 - 0xfe
    "11111110", --  627 - 0x273  :  254 - 0xfe
    "11111110", --  628 - 0x274  :  254 - 0xfe
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111110", --  631 - 0x277  :  254 - 0xfe
    "11111110", --  632 - 0x278  :  254 - 0xfe -- Sprite 0x4f
    "11111110", --  633 - 0x279  :  254 - 0xfe
    "11111110", --  634 - 0x27a  :  254 - 0xfe
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "11111110", --  636 - 0x27c  :  254 - 0xfe
    "11111110", --  637 - 0x27d  :  254 - 0xfe
    "11111110", --  638 - 0x27e  :  254 - 0xfe
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00010000", --  649 - 0x289  :   16 - 0x10
    "00010000", --  650 - 0x28a  :   16 - 0x10
    "01111100", --  651 - 0x28b  :  124 - 0x7c
    "00111000", --  652 - 0x28c  :   56 - 0x38
    "00111000", --  653 - 0x28d  :   56 - 0x38
    "01101100", --  654 - 0x28e  :  108 - 0x6c
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00010000", --  657 - 0x291  :   16 - 0x10
    "00010000", --  658 - 0x292  :   16 - 0x10
    "01111100", --  659 - 0x293  :  124 - 0x7c
    "00111000", --  660 - 0x294  :   56 - 0x38
    "00111000", --  661 - 0x295  :   56 - 0x38
    "01101100", --  662 - 0x296  :  108 - 0x6c
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "11111111", --  672 - 0x2a0  :  255 - 0xff -- Sprite 0x54
    "11111111", --  673 - 0x2a1  :  255 - 0xff
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111111", --  679 - 0x2a7  :  255 - 0xff
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Sprite 0x55
    "11111111", --  681 - 0x2a9  :  255 - 0xff
    "11111111", --  682 - 0x2aa  :  255 - 0xff
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11111111", --  684 - 0x2ac  :  255 - 0xff
    "11111111", --  685 - 0x2ad  :  255 - 0xff
    "11111111", --  686 - 0x2ae  :  255 - 0xff
    "11111111", --  687 - 0x2af  :  255 - 0xff
    "00000010", --  688 - 0x2b0  :    2 - 0x2 -- Sprite 0x56
    "00000101", --  689 - 0x2b1  :    5 - 0x5
    "10101010", --  690 - 0x2b2  :  170 - 0xaa
    "01010001", --  691 - 0x2b3  :   81 - 0x51
    "10101010", --  692 - 0x2b4  :  170 - 0xaa
    "01010001", --  693 - 0x2b5  :   81 - 0x51
    "10100010", --  694 - 0x2b6  :  162 - 0xa2
    "00000100", --  695 - 0x2b7  :    4 - 0x4
    "00001000", --  696 - 0x2b8  :    8 - 0x8 -- Sprite 0x57
    "01010101", --  697 - 0x2b9  :   85 - 0x55
    "00101010", --  698 - 0x2ba  :   42 - 0x2a
    "01010101", --  699 - 0x2bb  :   85 - 0x55
    "00101010", --  700 - 0x2bc  :   42 - 0x2a
    "01000101", --  701 - 0x2bd  :   69 - 0x45
    "00001010", --  702 - 0x2be  :   10 - 0xa
    "00010000", --  703 - 0x2bf  :   16 - 0x10
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x58
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "01011111", --  706 - 0x2c2  :   95 - 0x5f
    "01101111", --  707 - 0x2c3  :  111 - 0x6f
    "01110000", --  708 - 0x2c4  :  112 - 0x70
    "01110111", --  709 - 0x2c5  :  119 - 0x77
    "01110111", --  710 - 0x2c6  :  119 - 0x77
    "01110111", --  711 - 0x2c7  :  119 - 0x77
    "01110111", --  712 - 0x2c8  :  119 - 0x77 -- Sprite 0x59
    "01110111", --  713 - 0x2c9  :  119 - 0x77
    "01110111", --  714 - 0x2ca  :  119 - 0x77
    "01110000", --  715 - 0x2cb  :  112 - 0x70
    "01101111", --  716 - 0x2cc  :  111 - 0x6f
    "01011111", --  717 - 0x2cd  :   95 - 0x5f
    "00010101", --  718 - 0x2ce  :   21 - 0x15
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x5a
    "11111100", --  721 - 0x2d1  :  252 - 0xfc
    "11111000", --  722 - 0x2d2  :  248 - 0xf8
    "11110110", --  723 - 0x2d3  :  246 - 0xf6
    "00001100", --  724 - 0x2d4  :   12 - 0xc
    "11101110", --  725 - 0x2d5  :  238 - 0xee
    "11101100", --  726 - 0x2d6  :  236 - 0xec
    "11101110", --  727 - 0x2d7  :  238 - 0xee
    "11101100", --  728 - 0x2d8  :  236 - 0xec -- Sprite 0x5b
    "11101110", --  729 - 0x2d9  :  238 - 0xee
    "11101100", --  730 - 0x2da  :  236 - 0xec
    "00001110", --  731 - 0x2db  :   14 - 0xe
    "11110100", --  732 - 0x2dc  :  244 - 0xf4
    "11111010", --  733 - 0x2dd  :  250 - 0xfa
    "01010100", --  734 - 0x2de  :   84 - 0x54
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00011100", --  737 - 0x2e1  :   28 - 0x1c
    "00111110", --  738 - 0x2e2  :   62 - 0x3e
    "00111110", --  739 - 0x2e3  :   62 - 0x3e
    "00111110", --  740 - 0x2e4  :   62 - 0x3e
    "00011100", --  741 - 0x2e5  :   28 - 0x1c
    "00011100", --  742 - 0x2e6  :   28 - 0x1c
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Sprite 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "00010100", --  753 - 0x2f1  :   20 - 0x14
    "00110110", --  754 - 0x2f2  :   54 - 0x36
    "00111110", --  755 - 0x2f3  :   62 - 0x3e
    "00111110", --  756 - 0x2f4  :   62 - 0x3e
    "00011100", --  757 - 0x2f5  :   28 - 0x1c
    "00001000", --  758 - 0x2f6  :    8 - 0x8
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Sprite 0x5f
    "00010100", --  761 - 0x2f9  :   20 - 0x14
    "00011100", --  762 - 0x2fa  :   28 - 0x1c
    "00011100", --  763 - 0x2fb  :   28 - 0x1c
    "00011100", --  764 - 0x2fc  :   28 - 0x1c
    "00011100", --  765 - 0x2fd  :   28 - 0x1c
    "00011100", --  766 - 0x2fe  :   28 - 0x1c
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "01111111", --  769 - 0x301  :  127 - 0x7f
    "01111111", --  770 - 0x302  :  127 - 0x7f
    "01111111", --  771 - 0x303  :  127 - 0x7f
    "01111111", --  772 - 0x304  :  127 - 0x7f
    "01111111", --  773 - 0x305  :  127 - 0x7f
    "00101010", --  774 - 0x306  :   42 - 0x2a
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "10101010", --  782 - 0x30e  :  170 - 0xaa
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x62
    "11111110", --  785 - 0x311  :  254 - 0xfe
    "11111110", --  786 - 0x312  :  254 - 0xfe
    "11111110", --  787 - 0x313  :  254 - 0xfe
    "11111110", --  788 - 0x314  :  254 - 0xfe
    "11111110", --  789 - 0x315  :  254 - 0xfe
    "10101010", --  790 - 0x316  :  170 - 0xaa
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Sprite 0x63
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000001", --  802 - 0x322  :    1 - 0x1
    "00000001", --  803 - 0x323  :    1 - 0x1
    "00000011", --  804 - 0x324  :    3 - 0x3
    "00000011", --  805 - 0x325  :    3 - 0x3
    "00000111", --  806 - 0x326  :    7 - 0x7
    "00000111", --  807 - 0x327  :    7 - 0x7
    "00001111", --  808 - 0x328  :   15 - 0xf -- Sprite 0x65
    "00001111", --  809 - 0x329  :   15 - 0xf
    "00011111", --  810 - 0x32a  :   31 - 0x1f
    "00011111", --  811 - 0x32b  :   31 - 0x1f
    "00111111", --  812 - 0x32c  :   63 - 0x3f
    "00111111", --  813 - 0x32d  :   63 - 0x3f
    "01010101", --  814 - 0x32e  :   85 - 0x55
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "10000000", --  819 - 0x333  :  128 - 0x80
    "01000000", --  820 - 0x334  :   64 - 0x40
    "10000000", --  821 - 0x335  :  128 - 0x80
    "11000000", --  822 - 0x336  :  192 - 0xc0
    "11100000", --  823 - 0x337  :  224 - 0xe0
    "11010000", --  824 - 0x338  :  208 - 0xd0 -- Sprite 0x67
    "11100000", --  825 - 0x339  :  224 - 0xe0
    "11110000", --  826 - 0x33a  :  240 - 0xf0
    "11101000", --  827 - 0x33b  :  232 - 0xe8
    "11110100", --  828 - 0x33c  :  244 - 0xf4
    "11111000", --  829 - 0x33d  :  248 - 0xf8
    "01010100", --  830 - 0x33e  :   84 - 0x54
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- Sprite 0x6f
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Sprite 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Sprite 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Sprite 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Sprite 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Sprite 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x80
    "00000011", -- 1025 - 0x401  :    3 - 0x3
    "00001111", -- 1026 - 0x402  :   15 - 0xf
    "00011111", -- 1027 - 0x403  :   31 - 0x1f
    "00011111", -- 1028 - 0x404  :   31 - 0x1f
    "00111111", -- 1029 - 0x405  :   63 - 0x3f
    "00111111", -- 1030 - 0x406  :   63 - 0x3f
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Sprite 0x81
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x82
    "11000000", -- 1041 - 0x411  :  192 - 0xc0
    "11110000", -- 1042 - 0x412  :  240 - 0xf0
    "11110000", -- 1043 - 0x413  :  240 - 0xf0
    "11101100", -- 1044 - 0x414  :  236 - 0xec
    "11100000", -- 1045 - 0x415  :  224 - 0xe0
    "11111100", -- 1046 - 0x416  :  252 - 0xfc
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "11100000", -- 1054 - 0x41e  :  224 - 0xe0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Sprite 0x84
    "00000011", -- 1057 - 0x421  :    3 - 0x3
    "00001111", -- 1058 - 0x422  :   15 - 0xf
    "00011111", -- 1059 - 0x423  :   31 - 0x1f
    "00011111", -- 1060 - 0x424  :   31 - 0x1f
    "00111111", -- 1061 - 0x425  :   63 - 0x3f
    "00111111", -- 1062 - 0x426  :   63 - 0x3f
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Sprite 0x85
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00001000", -- 1069 - 0x42d  :    8 - 0x8
    "00001110", -- 1070 - 0x42e  :   14 - 0xe
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x86
    "11000000", -- 1073 - 0x431  :  192 - 0xc0
    "11110000", -- 1074 - 0x432  :  240 - 0xf0
    "11110000", -- 1075 - 0x433  :  240 - 0xf0
    "11101100", -- 1076 - 0x434  :  236 - 0xec
    "11100000", -- 1077 - 0x435  :  224 - 0xe0
    "11111100", -- 1078 - 0x436  :  252 - 0xfc
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Sprite 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000110", -- 1085 - 0x43d  :    6 - 0x6
    "00001100", -- 1086 - 0x43e  :   12 - 0xc
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x88
    "00000011", -- 1089 - 0x441  :    3 - 0x3
    "00000011", -- 1090 - 0x442  :    3 - 0x3
    "00000100", -- 1091 - 0x443  :    4 - 0x4
    "00001111", -- 1092 - 0x444  :   15 - 0xf
    "00011111", -- 1093 - 0x445  :   31 - 0x1f
    "01101111", -- 1094 - 0x446  :  111 - 0x6f
    "01101111", -- 1095 - 0x447  :  111 - 0x6f
    "01101111", -- 1096 - 0x448  :  111 - 0x6f -- Sprite 0x89
    "01101111", -- 1097 - 0x449  :  111 - 0x6f
    "00011111", -- 1098 - 0x44a  :   31 - 0x1f
    "00001111", -- 1099 - 0x44b  :   15 - 0xf
    "00000100", -- 1100 - 0x44c  :    4 - 0x4
    "00000011", -- 1101 - 0x44d  :    3 - 0x3
    "00000011", -- 1102 - 0x44e  :    3 - 0x3
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x8a
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00011000", -- 1106 - 0x452  :   24 - 0x18
    "00110111", -- 1107 - 0x453  :   55 - 0x37
    "00101111", -- 1108 - 0x454  :   47 - 0x2f
    "00011111", -- 1109 - 0x455  :   31 - 0x1f
    "00011111", -- 1110 - 0x456  :   31 - 0x1f
    "00011111", -- 1111 - 0x457  :   31 - 0x1f
    "00011111", -- 1112 - 0x458  :   31 - 0x1f -- Sprite 0x8b
    "00011111", -- 1113 - 0x459  :   31 - 0x1f
    "00011111", -- 1114 - 0x45a  :   31 - 0x1f
    "00101111", -- 1115 - 0x45b  :   47 - 0x2f
    "00110111", -- 1116 - 0x45c  :   55 - 0x37
    "00011000", -- 1117 - 0x45d  :   24 - 0x18
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x8c
    "00000011", -- 1121 - 0x461  :    3 - 0x3
    "00000001", -- 1122 - 0x462  :    1 - 0x1
    "00011001", -- 1123 - 0x463  :   25 - 0x19
    "00111001", -- 1124 - 0x464  :   57 - 0x39
    "00011011", -- 1125 - 0x465  :   27 - 0x1b
    "00001111", -- 1126 - 0x466  :   15 - 0xf
    "00001111", -- 1127 - 0x467  :   15 - 0xf
    "01111111", -- 1128 - 0x468  :  127 - 0x7f -- Sprite 0x8d
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "00111111", -- 1130 - 0x46a  :   63 - 0x3f
    "00010111", -- 1131 - 0x46b  :   23 - 0x17
    "00000110", -- 1132 - 0x46c  :    6 - 0x6
    "00000100", -- 1133 - 0x46d  :    4 - 0x4
    "00000111", -- 1134 - 0x46e  :    7 - 0x7
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Sprite 0x8e
    "11000000", -- 1137 - 0x471  :  192 - 0xc0
    "11110000", -- 1138 - 0x472  :  240 - 0xf0
    "10111000", -- 1139 - 0x473  :  184 - 0xb8
    "10011100", -- 1140 - 0x474  :  156 - 0x9c
    "11111100", -- 1141 - 0x475  :  252 - 0xfc
    "11111110", -- 1142 - 0x476  :  254 - 0xfe
    "11000000", -- 1143 - 0x477  :  192 - 0xc0
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- Sprite 0x8f
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111000", -- 1146 - 0x47a  :  248 - 0xf8
    "11110000", -- 1147 - 0x47b  :  240 - 0xf0
    "11000000", -- 1148 - 0x47c  :  192 - 0xc0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "10000000", -- 1151 - 0x47f  :  128 - 0x80
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000001", -- 1153 - 0x481  :    1 - 0x1
    "00001001", -- 1154 - 0x482  :    9 - 0x9
    "00011001", -- 1155 - 0x483  :   25 - 0x19
    "00011100", -- 1156 - 0x484  :   28 - 0x1c
    "00001101", -- 1157 - 0x485  :   13 - 0xd
    "00001111", -- 1158 - 0x486  :   15 - 0xf
    "00101111", -- 1159 - 0x487  :   47 - 0x2f
    "01111111", -- 1160 - 0x488  :  127 - 0x7f -- Sprite 0x91
    "01111111", -- 1161 - 0x489  :  127 - 0x7f
    "00111111", -- 1162 - 0x48a  :   63 - 0x3f
    "00011011", -- 1163 - 0x48b  :   27 - 0x1b
    "00000011", -- 1164 - 0x48c  :    3 - 0x3
    "00000011", -- 1165 - 0x48d  :    3 - 0x3
    "00000001", -- 1166 - 0x48e  :    1 - 0x1
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x92
    "11000000", -- 1169 - 0x491  :  192 - 0xc0
    "11110000", -- 1170 - 0x492  :  240 - 0xf0
    "11011000", -- 1171 - 0x493  :  216 - 0xd8
    "11001100", -- 1172 - 0x494  :  204 - 0xcc
    "11111100", -- 1173 - 0x495  :  252 - 0xfc
    "11111110", -- 1174 - 0x496  :  254 - 0xfe
    "11100000", -- 1175 - 0x497  :  224 - 0xe0
    "11111110", -- 1176 - 0x498  :  254 - 0xfe -- Sprite 0x93
    "11111110", -- 1177 - 0x499  :  254 - 0xfe
    "11111000", -- 1178 - 0x49a  :  248 - 0xf8
    "01110000", -- 1179 - 0x49b  :  112 - 0x70
    "01000000", -- 1180 - 0x49c  :   64 - 0x40
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "11000000", -- 1182 - 0x49e  :  192 - 0xc0
    "00100000", -- 1183 - 0x49f  :   32 - 0x20
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00001100", -- 1186 - 0x4a2  :   12 - 0xc
    "00001110", -- 1187 - 0x4a3  :   14 - 0xe
    "00000110", -- 1188 - 0x4a4  :    6 - 0x6
    "00100110", -- 1189 - 0x4a5  :   38 - 0x26
    "00110111", -- 1190 - 0x4a6  :   55 - 0x37
    "00110011", -- 1191 - 0x4a7  :   51 - 0x33
    "01111111", -- 1192 - 0x4a8  :  127 - 0x7f -- Sprite 0x95
    "01111111", -- 1193 - 0x4a9  :  127 - 0x7f
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00011111", -- 1195 - 0x4ab  :   31 - 0x1f
    "00001110", -- 1196 - 0x4ac  :   14 - 0xe
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "11000000", -- 1201 - 0x4b1  :  192 - 0xc0
    "11110000", -- 1202 - 0x4b2  :  240 - 0xf0
    "01101000", -- 1203 - 0x4b3  :  104 - 0x68
    "01100100", -- 1204 - 0x4b4  :  100 - 0x64
    "11111100", -- 1205 - 0x4b5  :  252 - 0xfc
    "11111110", -- 1206 - 0x4b6  :  254 - 0xfe
    "11110000", -- 1207 - 0x4b7  :  240 - 0xf0
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- Sprite 0x97
    "11111110", -- 1209 - 0x4b9  :  254 - 0xfe
    "11111100", -- 1210 - 0x4ba  :  252 - 0xfc
    "10110000", -- 1211 - 0x4bb  :  176 - 0xb0
    "11000000", -- 1212 - 0x4bc  :  192 - 0xc0
    "11000000", -- 1213 - 0x4bd  :  192 - 0xc0
    "01110000", -- 1214 - 0x4be  :  112 - 0x70
    "00001000", -- 1215 - 0x4bf  :    8 - 0x8
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x98
    "00000001", -- 1217 - 0x4c1  :    1 - 0x1
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000001", -- 1222 - 0x4c6  :    1 - 0x1
    "00000011", -- 1223 - 0x4c7  :    3 - 0x3
    "00000111", -- 1224 - 0x4c8  :    7 - 0x7 -- Sprite 0x99
    "00010111", -- 1225 - 0x4c9  :   23 - 0x17
    "00101111", -- 1226 - 0x4ca  :   47 - 0x2f
    "00011110", -- 1227 - 0x4cb  :   30 - 0x1e
    "00010001", -- 1228 - 0x4cc  :   17 - 0x11
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000001", -- 1230 - 0x4ce  :    1 - 0x1
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00010000", -- 1233 - 0x4d1  :   16 - 0x10
    "01111000", -- 1234 - 0x4d2  :  120 - 0x78
    "01110100", -- 1235 - 0x4d3  :  116 - 0x74
    "11111110", -- 1236 - 0x4d4  :  254 - 0xfe
    "11111000", -- 1237 - 0x4d5  :  248 - 0xf8
    "11111100", -- 1238 - 0x4d6  :  252 - 0xfc
    "11111000", -- 1239 - 0x4d7  :  248 - 0xf8
    "11111000", -- 1240 - 0x4d8  :  248 - 0xf8 -- Sprite 0x9b
    "11010000", -- 1241 - 0x4d9  :  208 - 0xd0
    "00110000", -- 1242 - 0x4da  :   48 - 0x30
    "01100000", -- 1243 - 0x4db  :   96 - 0x60
    "10000000", -- 1244 - 0x4dc  :  128 - 0x80
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Sprite 0x9c
    "00000001", -- 1249 - 0x4e1  :    1 - 0x1
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000001", -- 1254 - 0x4e6  :    1 - 0x1
    "00000011", -- 1255 - 0x4e7  :    3 - 0x3
    "00000111", -- 1256 - 0x4e8  :    7 - 0x7 -- Sprite 0x9d
    "00010111", -- 1257 - 0x4e9  :   23 - 0x17
    "00101111", -- 1258 - 0x4ea  :   47 - 0x2f
    "00011110", -- 1259 - 0x4eb  :   30 - 0x1e
    "00010000", -- 1260 - 0x4ec  :   16 - 0x10
    "00000100", -- 1261 - 0x4ed  :    4 - 0x4
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x9e
    "00010000", -- 1265 - 0x4f1  :   16 - 0x10
    "01111000", -- 1266 - 0x4f2  :  120 - 0x78
    "01110100", -- 1267 - 0x4f3  :  116 - 0x74
    "11111110", -- 1268 - 0x4f4  :  254 - 0xfe
    "11111000", -- 1269 - 0x4f5  :  248 - 0xf8
    "11111100", -- 1270 - 0x4f6  :  252 - 0xfc
    "11111000", -- 1271 - 0x4f7  :  248 - 0xf8
    "11111000", -- 1272 - 0x4f8  :  248 - 0xf8 -- Sprite 0x9f
    "11010000", -- 1273 - 0x4f9  :  208 - 0xd0
    "00110000", -- 1274 - 0x4fa  :   48 - 0x30
    "11000000", -- 1275 - 0x4fb  :  192 - 0xc0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0xa0
    "00000011", -- 1281 - 0x501  :    3 - 0x3
    "00001111", -- 1282 - 0x502  :   15 - 0xf
    "00011111", -- 1283 - 0x503  :   31 - 0x1f
    "00111111", -- 1284 - 0x504  :   63 - 0x3f
    "00111111", -- 1285 - 0x505  :   63 - 0x3f
    "01111111", -- 1286 - 0x506  :  127 - 0x7f
    "01111111", -- 1287 - 0x507  :  127 - 0x7f
    "01111111", -- 1288 - 0x508  :  127 - 0x7f -- Sprite 0xa1
    "01111111", -- 1289 - 0x509  :  127 - 0x7f
    "00111111", -- 1290 - 0x50a  :   63 - 0x3f
    "00111111", -- 1291 - 0x50b  :   63 - 0x3f
    "00011111", -- 1292 - 0x50c  :   31 - 0x1f
    "00000101", -- 1293 - 0x50d  :    5 - 0x5
    "00000010", -- 1294 - 0x50e  :    2 - 0x2
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Sprite 0xa2
    "11000000", -- 1297 - 0x511  :  192 - 0xc0
    "11110000", -- 1298 - 0x512  :  240 - 0xf0
    "11111000", -- 1299 - 0x513  :  248 - 0xf8
    "11111000", -- 1300 - 0x514  :  248 - 0xf8
    "11111100", -- 1301 - 0x515  :  252 - 0xfc
    "11111010", -- 1302 - 0x516  :  250 - 0xfa
    "11111100", -- 1303 - 0x517  :  252 - 0xfc
    "11111010", -- 1304 - 0x518  :  250 - 0xfa -- Sprite 0xa3
    "11110100", -- 1305 - 0x519  :  244 - 0xf4
    "11101000", -- 1306 - 0x51a  :  232 - 0xe8
    "11010100", -- 1307 - 0x51b  :  212 - 0xd4
    "10101000", -- 1308 - 0x51c  :  168 - 0xa8
    "01010000", -- 1309 - 0x51d  :   80 - 0x50
    "10000000", -- 1310 - 0x51e  :  128 - 0x80
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0xa4
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00001110", -- 1315 - 0x523  :   14 - 0xe
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00001010", -- 1317 - 0x525  :   10 - 0xa
    "01001010", -- 1318 - 0x526  :   74 - 0x4a
    "01100000", -- 1319 - 0x527  :   96 - 0x60
    "01111111", -- 1320 - 0x528  :  127 - 0x7f -- Sprite 0xa5
    "01111000", -- 1321 - 0x529  :  120 - 0x78
    "00110111", -- 1322 - 0x52a  :   55 - 0x37
    "00111011", -- 1323 - 0x52b  :   59 - 0x3b
    "00111100", -- 1324 - 0x52c  :   60 - 0x3c
    "00011111", -- 1325 - 0x52d  :   31 - 0x1f
    "00000111", -- 1326 - 0x52e  :    7 - 0x7
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "01110000", -- 1331 - 0x533  :  112 - 0x70
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "01010000", -- 1333 - 0x535  :   80 - 0x50
    "01010010", -- 1334 - 0x536  :   82 - 0x52
    "00000110", -- 1335 - 0x537  :    6 - 0x6
    "11111100", -- 1336 - 0x538  :  252 - 0xfc -- Sprite 0xa7
    "00011010", -- 1337 - 0x539  :   26 - 0x1a
    "11101100", -- 1338 - 0x53a  :  236 - 0xec
    "11011000", -- 1339 - 0x53b  :  216 - 0xd8
    "00110100", -- 1340 - 0x53c  :   52 - 0x34
    "11101000", -- 1341 - 0x53d  :  232 - 0xe8
    "11000000", -- 1342 - 0x53e  :  192 - 0xc0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00001110", -- 1347 - 0x543  :   14 - 0xe
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00001110", -- 1349 - 0x545  :   14 - 0xe
    "01001010", -- 1350 - 0x546  :   74 - 0x4a
    "01100000", -- 1351 - 0x547  :   96 - 0x60
    "01111111", -- 1352 - 0x548  :  127 - 0x7f -- Sprite 0xa9
    "01111100", -- 1353 - 0x549  :  124 - 0x7c
    "01111011", -- 1354 - 0x54a  :  123 - 0x7b
    "01110111", -- 1355 - 0x54b  :  119 - 0x77
    "01111000", -- 1356 - 0x54c  :  120 - 0x78
    "01111111", -- 1357 - 0x54d  :  127 - 0x7f
    "01111111", -- 1358 - 0x54e  :  127 - 0x7f
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "01110000", -- 1363 - 0x553  :  112 - 0x70
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "01110000", -- 1365 - 0x555  :  112 - 0x70
    "01010010", -- 1366 - 0x556  :   82 - 0x52
    "00000110", -- 1367 - 0x557  :    6 - 0x6
    "11111100", -- 1368 - 0x558  :  252 - 0xfc -- Sprite 0xab
    "00111010", -- 1369 - 0x559  :   58 - 0x3a
    "11011100", -- 1370 - 0x55a  :  220 - 0xdc
    "11101010", -- 1371 - 0x55b  :  234 - 0xea
    "00011100", -- 1372 - 0x55c  :   28 - 0x1c
    "11111010", -- 1373 - 0x55d  :  250 - 0xfa
    "11110100", -- 1374 - 0x55e  :  244 - 0xf4
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000011", -- 1377 - 0x561  :    3 - 0x3
    "00001111", -- 1378 - 0x562  :   15 - 0xf
    "00001111", -- 1379 - 0x563  :   15 - 0xf
    "00011111", -- 1380 - 0x564  :   31 - 0x1f
    "01011111", -- 1381 - 0x565  :   95 - 0x5f
    "01010000", -- 1382 - 0x566  :   80 - 0x50
    "00010000", -- 1383 - 0x567  :   16 - 0x10
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Sprite 0xad
    "11111010", -- 1385 - 0x569  :  250 - 0xfa
    "11111010", -- 1386 - 0x56a  :  250 - 0xfa
    "11111010", -- 1387 - 0x56b  :  250 - 0xfa
    "10111010", -- 1388 - 0x56c  :  186 - 0xba
    "10011010", -- 1389 - 0x56d  :  154 - 0x9a
    "00001010", -- 1390 - 0x56e  :   10 - 0xa
    "00000010", -- 1391 - 0x56f  :    2 - 0x2
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00001111", -- 1394 - 0x572  :   15 - 0xf
    "00001111", -- 1395 - 0x573  :   15 - 0xf
    "00011111", -- 1396 - 0x574  :   31 - 0x1f
    "01011111", -- 1397 - 0x575  :   95 - 0x5f
    "01010000", -- 1398 - 0x576  :   80 - 0x50
    "00010111", -- 1399 - 0x577  :   23 - 0x17
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "11111010", -- 1401 - 0x579  :  250 - 0xfa
    "11111010", -- 1402 - 0x57a  :  250 - 0xfa
    "11111010", -- 1403 - 0x57b  :  250 - 0xfa
    "00111010", -- 1404 - 0x57c  :   58 - 0x3a
    "01011010", -- 1405 - 0x57d  :   90 - 0x5a
    "01101010", -- 1406 - 0x57e  :  106 - 0x6a
    "11110010", -- 1407 - 0x57f  :  242 - 0xf2
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000011", -- 1410 - 0x582  :    3 - 0x3
    "00001111", -- 1411 - 0x583  :   15 - 0xf
    "00111011", -- 1412 - 0x584  :   59 - 0x3b
    "00111111", -- 1413 - 0x585  :   63 - 0x3f
    "01101111", -- 1414 - 0x586  :  111 - 0x6f
    "01111101", -- 1415 - 0x587  :  125 - 0x7d
    "00001111", -- 1416 - 0x588  :   15 - 0xf -- Sprite 0xb1
    "01110000", -- 1417 - 0x589  :  112 - 0x70
    "01111111", -- 1418 - 0x58a  :  127 - 0x7f
    "00001111", -- 1419 - 0x58b  :   15 - 0xf
    "01110000", -- 1420 - 0x58c  :  112 - 0x70
    "01111111", -- 1421 - 0x58d  :  127 - 0x7f
    "00001111", -- 1422 - 0x58e  :   15 - 0xf
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0xb2
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "11000000", -- 1426 - 0x592  :  192 - 0xc0
    "11110000", -- 1427 - 0x593  :  240 - 0xf0
    "10111100", -- 1428 - 0x594  :  188 - 0xbc
    "11110100", -- 1429 - 0x595  :  244 - 0xf4
    "11111110", -- 1430 - 0x596  :  254 - 0xfe
    "11011110", -- 1431 - 0x597  :  222 - 0xde
    "11110000", -- 1432 - 0x598  :  240 - 0xf0 -- Sprite 0xb3
    "00001110", -- 1433 - 0x599  :   14 - 0xe
    "11111110", -- 1434 - 0x59a  :  254 - 0xfe
    "11110000", -- 1435 - 0x59b  :  240 - 0xf0
    "00001110", -- 1436 - 0x59c  :   14 - 0xe
    "11111110", -- 1437 - 0x59d  :  254 - 0xfe
    "11110000", -- 1438 - 0x59e  :  240 - 0xf0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000011", -- 1442 - 0x5a2  :    3 - 0x3
    "00001111", -- 1443 - 0x5a3  :   15 - 0xf
    "00111011", -- 1444 - 0x5a4  :   59 - 0x3b
    "00111111", -- 1445 - 0x5a5  :   63 - 0x3f
    "01101111", -- 1446 - 0x5a6  :  111 - 0x6f
    "01111101", -- 1447 - 0x5a7  :  125 - 0x7d
    "00001111", -- 1448 - 0x5a8  :   15 - 0xf -- Sprite 0xb5
    "01110000", -- 1449 - 0x5a9  :  112 - 0x70
    "01111111", -- 1450 - 0x5aa  :  127 - 0x7f
    "00001111", -- 1451 - 0x5ab  :   15 - 0xf
    "01110000", -- 1452 - 0x5ac  :  112 - 0x70
    "01111111", -- 1453 - 0x5ad  :  127 - 0x7f
    "00001111", -- 1454 - 0x5ae  :   15 - 0xf
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "11000000", -- 1458 - 0x5b2  :  192 - 0xc0
    "11110000", -- 1459 - 0x5b3  :  240 - 0xf0
    "10111100", -- 1460 - 0x5b4  :  188 - 0xbc
    "11110100", -- 1461 - 0x5b5  :  244 - 0xf4
    "11111110", -- 1462 - 0x5b6  :  254 - 0xfe
    "11011110", -- 1463 - 0x5b7  :  222 - 0xde
    "11110000", -- 1464 - 0x5b8  :  240 - 0xf0 -- Sprite 0xb7
    "00001110", -- 1465 - 0x5b9  :   14 - 0xe
    "11111110", -- 1466 - 0x5ba  :  254 - 0xfe
    "11110000", -- 1467 - 0x5bb  :  240 - 0xf0
    "00001110", -- 1468 - 0x5bc  :   14 - 0xe
    "11111110", -- 1469 - 0x5bd  :  254 - 0xfe
    "11110000", -- 1470 - 0x5be  :  240 - 0xf0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0xb8
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000011", -- 1474 - 0x5c2  :    3 - 0x3
    "00001111", -- 1475 - 0x5c3  :   15 - 0xf
    "00111011", -- 1476 - 0x5c4  :   59 - 0x3b
    "00111111", -- 1477 - 0x5c5  :   63 - 0x3f
    "01101111", -- 1478 - 0x5c6  :  111 - 0x6f
    "01111101", -- 1479 - 0x5c7  :  125 - 0x7d
    "00001111", -- 1480 - 0x5c8  :   15 - 0xf -- Sprite 0xb9
    "00100000", -- 1481 - 0x5c9  :   32 - 0x20
    "01010101", -- 1482 - 0x5ca  :   85 - 0x55
    "00001010", -- 1483 - 0x5cb  :   10 - 0xa
    "01110000", -- 1484 - 0x5cc  :  112 - 0x70
    "01111111", -- 1485 - 0x5cd  :  127 - 0x7f
    "00001111", -- 1486 - 0x5ce  :   15 - 0xf
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0xba
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "11000000", -- 1490 - 0x5d2  :  192 - 0xc0
    "11110000", -- 1491 - 0x5d3  :  240 - 0xf0
    "10111100", -- 1492 - 0x5d4  :  188 - 0xbc
    "11110100", -- 1493 - 0x5d5  :  244 - 0xf4
    "11111110", -- 1494 - 0x5d6  :  254 - 0xfe
    "11011110", -- 1495 - 0x5d7  :  222 - 0xde
    "11110000", -- 1496 - 0x5d8  :  240 - 0xf0 -- Sprite 0xbb
    "00001010", -- 1497 - 0x5d9  :   10 - 0xa
    "01010100", -- 1498 - 0x5da  :   84 - 0x54
    "10100000", -- 1499 - 0x5db  :  160 - 0xa0
    "00001110", -- 1500 - 0x5dc  :   14 - 0xe
    "11111110", -- 1501 - 0x5dd  :  254 - 0xfe
    "11110000", -- 1502 - 0x5de  :  240 - 0xf0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0xbc
    "01110011", -- 1505 - 0x5e1  :  115 - 0x73
    "01111011", -- 1506 - 0x5e2  :  123 - 0x7b
    "01111111", -- 1507 - 0x5e3  :  127 - 0x7f
    "00111111", -- 1508 - 0x5e4  :   63 - 0x3f
    "00011100", -- 1509 - 0x5e5  :   28 - 0x1c
    "01111011", -- 1510 - 0x5e6  :  123 - 0x7b
    "01111011", -- 1511 - 0x5e7  :  123 - 0x7b
    "01111011", -- 1512 - 0x5e8  :  123 - 0x7b -- Sprite 0xbd
    "01111011", -- 1513 - 0x5e9  :  123 - 0x7b
    "00011100", -- 1514 - 0x5ea  :   28 - 0x1c
    "00111111", -- 1515 - 0x5eb  :   63 - 0x3f
    "01111111", -- 1516 - 0x5ec  :  127 - 0x7f
    "01111011", -- 1517 - 0x5ed  :  123 - 0x7b
    "01110011", -- 1518 - 0x5ee  :  115 - 0x73
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "11001110", -- 1521 - 0x5f1  :  206 - 0xce
    "11011110", -- 1522 - 0x5f2  :  222 - 0xde
    "11111110", -- 1523 - 0x5f3  :  254 - 0xfe
    "11111100", -- 1524 - 0x5f4  :  252 - 0xfc
    "00111000", -- 1525 - 0x5f5  :   56 - 0x38
    "11011110", -- 1526 - 0x5f6  :  222 - 0xde
    "11011110", -- 1527 - 0x5f7  :  222 - 0xde
    "11011110", -- 1528 - 0x5f8  :  222 - 0xde -- Sprite 0xbf
    "11011110", -- 1529 - 0x5f9  :  222 - 0xde
    "00111000", -- 1530 - 0x5fa  :   56 - 0x38
    "11111100", -- 1531 - 0x5fb  :  252 - 0xfc
    "11111110", -- 1532 - 0x5fc  :  254 - 0xfe
    "11011110", -- 1533 - 0x5fd  :  222 - 0xde
    "11001110", -- 1534 - 0x5fe  :  206 - 0xce
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "01000000", -- 1538 - 0x602  :   64 - 0x40
    "01100000", -- 1539 - 0x603  :   96 - 0x60
    "01100001", -- 1540 - 0x604  :   97 - 0x61
    "00000010", -- 1541 - 0x605  :    2 - 0x2
    "00000010", -- 1542 - 0x606  :    2 - 0x2
    "00000111", -- 1543 - 0x607  :    7 - 0x7
    "00000111", -- 1544 - 0x608  :    7 - 0x7 -- Sprite 0xc1
    "00000100", -- 1545 - 0x609  :    4 - 0x4
    "00000111", -- 1546 - 0x60a  :    7 - 0x7
    "00000001", -- 1547 - 0x60b  :    1 - 0x1
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00010000", -- 1549 - 0x60d  :   16 - 0x10
    "00101000", -- 1550 - 0x60e  :   40 - 0x28
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000010", -- 1554 - 0x612  :    2 - 0x2
    "00000110", -- 1555 - 0x613  :    6 - 0x6
    "11100110", -- 1556 - 0x614  :  230 - 0xe6
    "10100000", -- 1557 - 0x615  :  160 - 0xa0
    "10100000", -- 1558 - 0x616  :  160 - 0xa0
    "11110000", -- 1559 - 0x617  :  240 - 0xf0
    "11110000", -- 1560 - 0x618  :  240 - 0xf0 -- Sprite 0xc3
    "00110000", -- 1561 - 0x619  :   48 - 0x30
    "11000000", -- 1562 - 0x61a  :  192 - 0xc0
    "10000000", -- 1563 - 0x61b  :  128 - 0x80
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00001000", -- 1565 - 0x61d  :    8 - 0x8
    "00010100", -- 1566 - 0x61e  :   20 - 0x14
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000101", -- 1569 - 0x621  :    5 - 0x5
    "00000111", -- 1570 - 0x622  :    7 - 0x7
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000001", -- 1575 - 0x627  :    1 - 0x1
    "00000010", -- 1576 - 0x628  :    2 - 0x2 -- Sprite 0xc5
    "00000111", -- 1577 - 0x629  :    7 - 0x7
    "00100111", -- 1578 - 0x62a  :   39 - 0x27
    "01010011", -- 1579 - 0x62b  :   83 - 0x53
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000010", -- 1581 - 0x62d  :    2 - 0x2
    "00000101", -- 1582 - 0x62e  :    5 - 0x5
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "01100000", -- 1589 - 0x635  :   96 - 0x60
    "11011000", -- 1590 - 0x636  :  216 - 0xd8
    "10110000", -- 1591 - 0x637  :  176 - 0xb0
    "11101000", -- 1592 - 0x638  :  232 - 0xe8 -- Sprite 0xc7
    "01111000", -- 1593 - 0x639  :  120 - 0x78
    "10110110", -- 1594 - 0x63a  :  182 - 0xb6
    "11100100", -- 1595 - 0x63b  :  228 - 0xe4
    "00000110", -- 1596 - 0x63c  :    6 - 0x6
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "01000000", -- 1602 - 0x642  :   64 - 0x40
    "00100000", -- 1603 - 0x643  :   32 - 0x20
    "01000000", -- 1604 - 0x644  :   64 - 0x40
    "00000111", -- 1605 - 0x645  :    7 - 0x7
    "00000101", -- 1606 - 0x646  :    5 - 0x5
    "00001101", -- 1607 - 0x647  :   13 - 0xd
    "00001101", -- 1608 - 0x648  :   13 - 0xd -- Sprite 0xc9
    "00000101", -- 1609 - 0x649  :    5 - 0x5
    "00000011", -- 1610 - 0x64a  :    3 - 0x3
    "01000011", -- 1611 - 0x64b  :   67 - 0x43
    "00100000", -- 1612 - 0x64c  :   32 - 0x20
    "01000000", -- 1613 - 0x64d  :   64 - 0x40
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00011100", -- 1617 - 0x651  :   28 - 0x1c
    "00011000", -- 1618 - 0x652  :   24 - 0x18
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "10000000", -- 1621 - 0x655  :  128 - 0x80
    "11100000", -- 1622 - 0x656  :  224 - 0xe0
    "10010000", -- 1623 - 0x657  :  144 - 0x90
    "11110000", -- 1624 - 0x658  :  240 - 0xf0 -- Sprite 0xcb
    "10010000", -- 1625 - 0x659  :  144 - 0x90
    "11110000", -- 1626 - 0x65a  :  240 - 0xf0
    "10000000", -- 1627 - 0x65b  :  128 - 0x80
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00011000", -- 1629 - 0x65d  :   24 - 0x18
    "00011100", -- 1630 - 0x65e  :   28 - 0x1c
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00001000", -- 1633 - 0x661  :    8 - 0x8
    "00000100", -- 1634 - 0x662  :    4 - 0x4
    "00001000", -- 1635 - 0x663  :    8 - 0x8
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "01000110", -- 1637 - 0x665  :   70 - 0x46
    "00101111", -- 1638 - 0x666  :   47 - 0x2f
    "01001110", -- 1639 - 0x667  :   78 - 0x4e
    "00001101", -- 1640 - 0x668  :   13 - 0xd -- Sprite 0xcd
    "00001011", -- 1641 - 0x669  :   11 - 0xb
    "00001111", -- 1642 - 0x66a  :   15 - 0xf
    "00000110", -- 1643 - 0x66b  :    6 - 0x6
    "00000011", -- 1644 - 0x66c  :    3 - 0x3
    "00011100", -- 1645 - 0x66d  :   28 - 0x1c
    "00010100", -- 1646 - 0x66e  :   20 - 0x14
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000110", -- 1653 - 0x675  :    6 - 0x6
    "00000100", -- 1654 - 0x676  :    4 - 0x4
    "10000110", -- 1655 - 0x677  :  134 - 0x86
    "11000000", -- 1656 - 0x678  :  192 - 0xc0 -- Sprite 0xcf
    "01100000", -- 1657 - 0x679  :   96 - 0x60
    "10100000", -- 1658 - 0x67a  :  160 - 0xa0
    "11000000", -- 1659 - 0x67b  :  192 - 0xc0
    "01000000", -- 1660 - 0x67c  :   64 - 0x40
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000100", -- 1668 - 0x684  :    4 - 0x4
    "00001110", -- 1669 - 0x685  :   14 - 0xe
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111001", -- 1671 - 0x687  :   57 - 0x39
    "01110000", -- 1672 - 0x688  :  112 - 0x70 -- Sprite 0xd1
    "01111000", -- 1673 - 0x689  :  120 - 0x78
    "00111111", -- 1674 - 0x68a  :   63 - 0x3f
    "00111111", -- 1675 - 0x68b  :   63 - 0x3f
    "00000011", -- 1676 - 0x68c  :    3 - 0x3
    "00001100", -- 1677 - 0x68d  :   12 - 0xc
    "00001110", -- 1678 - 0x68e  :   14 - 0xe
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0xd2
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00001000", -- 1683 - 0x693  :    8 - 0x8
    "11011000", -- 1684 - 0x694  :  216 - 0xd8
    "11111100", -- 1685 - 0x695  :  252 - 0xfc
    "11111100", -- 1686 - 0x696  :  252 - 0xfc
    "10011100", -- 1687 - 0x697  :  156 - 0x9c
    "00001100", -- 1688 - 0x698  :   12 - 0xc -- Sprite 0xd3
    "10011100", -- 1689 - 0x699  :  156 - 0x9c
    "11111000", -- 1690 - 0x69a  :  248 - 0xf8
    "01111000", -- 1691 - 0x69b  :  120 - 0x78
    "10001000", -- 1692 - 0x69c  :  136 - 0x88
    "00110000", -- 1693 - 0x69d  :   48 - 0x30
    "00111000", -- 1694 - 0x69e  :   56 - 0x38
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000001", -- 1700 - 0x6a4  :    1 - 0x1
    "00001011", -- 1701 - 0x6a5  :   11 - 0xb
    "00011111", -- 1702 - 0x6a6  :   31 - 0x1f
    "00111001", -- 1703 - 0x6a7  :   57 - 0x39
    "01110000", -- 1704 - 0x6a8  :  112 - 0x70 -- Sprite 0xd5
    "01111000", -- 1705 - 0x6a9  :  120 - 0x78
    "00111111", -- 1706 - 0x6aa  :   63 - 0x3f
    "00111111", -- 1707 - 0x6ab  :   63 - 0x3f
    "00000011", -- 1708 - 0x6ac  :    3 - 0x3
    "00111000", -- 1709 - 0x6ad  :   56 - 0x38
    "00011100", -- 1710 - 0x6ae  :   28 - 0x1c
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "11000000", -- 1715 - 0x6b3  :  192 - 0xc0
    "11001000", -- 1716 - 0x6b4  :  200 - 0xc8
    "11111000", -- 1717 - 0x6b5  :  248 - 0xf8
    "11111100", -- 1718 - 0x6b6  :  252 - 0xfc
    "10011100", -- 1719 - 0x6b7  :  156 - 0x9c
    "00001100", -- 1720 - 0x6b8  :   12 - 0xc -- Sprite 0xd7
    "10011100", -- 1721 - 0x6b9  :  156 - 0x9c
    "11111000", -- 1722 - 0x6ba  :  248 - 0xf8
    "01111000", -- 1723 - 0x6bb  :  120 - 0x78
    "11100010", -- 1724 - 0x6bc  :  226 - 0xe2
    "00011110", -- 1725 - 0x6bd  :   30 - 0x1e
    "00001100", -- 1726 - 0x6be  :   12 - 0xc
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0xd8
    "00110000", -- 1729 - 0x6c1  :   48 - 0x30
    "00111100", -- 1730 - 0x6c2  :   60 - 0x3c
    "01111100", -- 1731 - 0x6c3  :  124 - 0x7c
    "01111100", -- 1732 - 0x6c4  :  124 - 0x7c
    "00111110", -- 1733 - 0x6c5  :   62 - 0x3e
    "00011100", -- 1734 - 0x6c6  :   28 - 0x1c
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- Sprite 0xd9
    "00001110", -- 1737 - 0x6c9  :   14 - 0xe
    "00111110", -- 1738 - 0x6ca  :   62 - 0x3e
    "01111110", -- 1739 - 0x6cb  :  126 - 0x7e
    "01111110", -- 1740 - 0x6cc  :  126 - 0x7e
    "00111100", -- 1741 - 0x6cd  :   60 - 0x3c
    "00001100", -- 1742 - 0x6ce  :   12 - 0xc
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0xda
    "00100000", -- 1745 - 0x6d1  :   32 - 0x20
    "01111110", -- 1746 - 0x6d2  :  126 - 0x7e
    "01111110", -- 1747 - 0x6d3  :  126 - 0x7e
    "01111110", -- 1748 - 0x6d4  :  126 - 0x7e
    "00111100", -- 1749 - 0x6d5  :   60 - 0x3c
    "00111000", -- 1750 - 0x6d6  :   56 - 0x38
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- Sprite 0xdb
    "00011100", -- 1753 - 0x6d9  :   28 - 0x1c
    "00111110", -- 1754 - 0x6da  :   62 - 0x3e
    "01111110", -- 1755 - 0x6db  :  126 - 0x7e
    "01111110", -- 1756 - 0x6dc  :  126 - 0x7e
    "00111100", -- 1757 - 0x6dd  :   60 - 0x3c
    "00010000", -- 1758 - 0x6de  :   16 - 0x10
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000001", -- 1763 - 0x6e3  :    1 - 0x1
    "00000011", -- 1764 - 0x6e4  :    3 - 0x3
    "00000001", -- 1765 - 0x6e5  :    1 - 0x1
    "00000001", -- 1766 - 0x6e6  :    1 - 0x1
    "00001111", -- 1767 - 0x6e7  :   15 - 0xf
    "00000111", -- 1768 - 0x6e8  :    7 - 0x7 -- Sprite 0xdd
    "00000111", -- 1769 - 0x6e9  :    7 - 0x7
    "00000111", -- 1770 - 0x6ea  :    7 - 0x7
    "00011111", -- 1771 - 0x6eb  :   31 - 0x1f
    "00001111", -- 1772 - 0x6ec  :   15 - 0xf
    "00000111", -- 1773 - 0x6ed  :    7 - 0x7
    "00000011", -- 1774 - 0x6ee  :    3 - 0x3
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0xde
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "10000000", -- 1780 - 0x6f4  :  128 - 0x80
    "10000000", -- 1781 - 0x6f5  :  128 - 0x80
    "10010000", -- 1782 - 0x6f6  :  144 - 0x90
    "11110000", -- 1783 - 0x6f7  :  240 - 0xf0
    "11100000", -- 1784 - 0x6f8  :  224 - 0xe0 -- Sprite 0xdf
    "11100000", -- 1785 - 0x6f9  :  224 - 0xe0
    "11110000", -- 1786 - 0x6fa  :  240 - 0xf0
    "11110000", -- 1787 - 0x6fb  :  240 - 0xf0
    "11100000", -- 1788 - 0x6fc  :  224 - 0xe0
    "11000000", -- 1789 - 0x6fd  :  192 - 0xc0
    "11000000", -- 1790 - 0x6fe  :  192 - 0xc0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00001111", -- 1792 - 0x700  :   15 - 0xf -- Sprite 0xe0
    "00011111", -- 1793 - 0x701  :   31 - 0x1f
    "00011111", -- 1794 - 0x702  :   31 - 0x1f
    "00111111", -- 1795 - 0x703  :   63 - 0x3f
    "01111111", -- 1796 - 0x704  :  127 - 0x7f
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "01111111", -- 1802 - 0x70a  :  127 - 0x7f
    "00111111", -- 1803 - 0x70b  :   63 - 0x3f
    "00111111", -- 1804 - 0x70c  :   63 - 0x3f
    "00011111", -- 1805 - 0x70d  :   31 - 0x1f
    "00001111", -- 1806 - 0x70e  :   15 - 0xf
    "00000111", -- 1807 - 0x70f  :    7 - 0x7
    "11111110", -- 1808 - 0x710  :  254 - 0xfe -- Sprite 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "00001111", -- 1811 - 0x713  :   15 - 0xf
    "10111111", -- 1812 - 0x714  :  191 - 0xbf
    "10100011", -- 1813 - 0x715  :  163 - 0xa3
    "11110111", -- 1814 - 0x716  :  247 - 0xf7
    "11110111", -- 1815 - 0x717  :  247 - 0xf7
    "11111111", -- 1816 - 0x718  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "00111111", -- 1818 - 0x71a  :   63 - 0x3f
    "00011111", -- 1819 - 0x71b  :   31 - 0x1f
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111100", -- 1821 - 0x71d  :  252 - 0xfc
    "11111000", -- 1822 - 0x71e  :  248 - 0xf8
    "11110000", -- 1823 - 0x71f  :  240 - 0xf0
    "00001111", -- 1824 - 0x720  :   15 - 0xf -- Sprite 0xe4
    "00011111", -- 1825 - 0x721  :   31 - 0x1f
    "00011111", -- 1826 - 0x722  :   31 - 0x1f
    "00111111", -- 1827 - 0x723  :   63 - 0x3f
    "01111111", -- 1828 - 0x724  :  127 - 0x7f
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "01111110", -- 1834 - 0x72a  :  126 - 0x7e
    "00111111", -- 1835 - 0x72b  :   63 - 0x3f
    "00111111", -- 1836 - 0x72c  :   63 - 0x3f
    "00011111", -- 1837 - 0x72d  :   31 - 0x1f
    "00001111", -- 1838 - 0x72e  :   15 - 0xf
    "00000111", -- 1839 - 0x72f  :    7 - 0x7
    "11111110", -- 1840 - 0x730  :  254 - 0xfe -- Sprite 0xe6
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11100011", -- 1843 - 0x733  :  227 - 0xe3
    "00010111", -- 1844 - 0x734  :   23 - 0x17
    "10110111", -- 1845 - 0x735  :  183 - 0xb7
    "10111111", -- 1846 - 0x736  :  191 - 0xbf
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "00111111", -- 1850 - 0x73a  :   63 - 0x3f
    "00001111", -- 1851 - 0x73b  :   15 - 0xf
    "00001110", -- 1852 - 0x73c  :   14 - 0xe
    "11111100", -- 1853 - 0x73d  :  252 - 0xfc
    "11111000", -- 1854 - 0x73e  :  248 - 0xf8
    "11110000", -- 1855 - 0x73f  :  240 - 0xf0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "00000101", -- 1857 - 0x741  :    5 - 0x5
    "00000111", -- 1858 - 0x742  :    7 - 0x7
    "00000011", -- 1859 - 0x743  :    3 - 0x3
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Sprite 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000011", -- 1872 - 0x750  :    3 - 0x3 -- Sprite 0xea
    "10011110", -- 1873 - 0x751  :  158 - 0x9e
    "00001110", -- 1874 - 0x752  :   14 - 0xe
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000100", -- 1892 - 0x764  :    4 - 0x4
    "00001110", -- 1893 - 0x765  :   14 - 0xe
    "00001111", -- 1894 - 0x766  :   15 - 0xf
    "00001011", -- 1895 - 0x767  :   11 - 0xb
    "00001111", -- 1896 - 0x768  :   15 - 0xf -- Sprite 0xed
    "00001100", -- 1897 - 0x769  :   12 - 0xc
    "00001111", -- 1898 - 0x76a  :   15 - 0xf
    "00001111", -- 1899 - 0x76b  :   15 - 0xf
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "01111111", -- 1901 - 0x76d  :  127 - 0x7f
    "11010101", -- 1902 - 0x76e  :  213 - 0xd5
    "01111111", -- 1903 - 0x76f  :  127 - 0x7f
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00100000", -- 1908 - 0x774  :   32 - 0x20
    "01110000", -- 1909 - 0x775  :  112 - 0x70
    "11110000", -- 1910 - 0x776  :  240 - 0xf0
    "11100000", -- 1911 - 0x777  :  224 - 0xe0
    "11110000", -- 1912 - 0x778  :  240 - 0xf0 -- Sprite 0xef
    "00110000", -- 1913 - 0x779  :   48 - 0x30
    "11110000", -- 1914 - 0x77a  :  240 - 0xf0
    "11110000", -- 1915 - 0x77b  :  240 - 0xf0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "11111110", -- 1917 - 0x77d  :  254 - 0xfe
    "01010101", -- 1918 - 0x77e  :   85 - 0x55
    "11111110", -- 1919 - 0x77f  :  254 - 0xfe
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000100", -- 1924 - 0x784  :    4 - 0x4
    "00001110", -- 1925 - 0x785  :   14 - 0xe
    "00001111", -- 1926 - 0x786  :   15 - 0xf
    "00001011", -- 1927 - 0x787  :   11 - 0xb
    "00001111", -- 1928 - 0x788  :   15 - 0xf -- Sprite 0xf1
    "00001100", -- 1929 - 0x789  :   12 - 0xc
    "00001111", -- 1930 - 0x78a  :   15 - 0xf
    "00001111", -- 1931 - 0x78b  :   15 - 0xf
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "01111111", -- 1933 - 0x78d  :  127 - 0x7f
    "10101010", -- 1934 - 0x78e  :  170 - 0xaa
    "01111111", -- 1935 - 0x78f  :  127 - 0x7f
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00100000", -- 1940 - 0x794  :   32 - 0x20
    "01110000", -- 1941 - 0x795  :  112 - 0x70
    "11110000", -- 1942 - 0x796  :  240 - 0xf0
    "11100000", -- 1943 - 0x797  :  224 - 0xe0
    "11110000", -- 1944 - 0x798  :  240 - 0xf0 -- Sprite 0xf3
    "00110000", -- 1945 - 0x799  :   48 - 0x30
    "11110000", -- 1946 - 0x79a  :  240 - 0xf0
    "11110000", -- 1947 - 0x79b  :  240 - 0xf0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "11111110", -- 1949 - 0x79d  :  254 - 0xfe
    "10101011", -- 1950 - 0x79e  :  171 - 0xab
    "11111110", -- 1951 - 0x79f  :  254 - 0xfe
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "00010101", -- 1953 - 0x7a1  :   21 - 0x15
    "00001010", -- 1954 - 0x7a2  :   10 - 0xa
    "00000101", -- 1955 - 0x7a3  :    5 - 0x5
    "00000010", -- 1956 - 0x7a4  :    2 - 0x2
    "00000101", -- 1957 - 0x7a5  :    5 - 0x5
    "00000111", -- 1958 - 0x7a6  :    7 - 0x7
    "00000111", -- 1959 - 0x7a7  :    7 - 0x7
    "00111100", -- 1960 - 0x7a8  :   60 - 0x3c -- Sprite 0xf5
    "01111011", -- 1961 - 0x7a9  :  123 - 0x7b
    "01111011", -- 1962 - 0x7aa  :  123 - 0x7b
    "01111111", -- 1963 - 0x7ab  :  127 - 0x7f
    "01111110", -- 1964 - 0x7ac  :  126 - 0x7e
    "01111111", -- 1965 - 0x7ad  :  127 - 0x7f
    "00111110", -- 1966 - 0x7ae  :   62 - 0x3e
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "01010000", -- 1969 - 0x7b1  :   80 - 0x50
    "10100000", -- 1970 - 0x7b2  :  160 - 0xa0
    "01000000", -- 1971 - 0x7b3  :   64 - 0x40
    "10100000", -- 1972 - 0x7b4  :  160 - 0xa0
    "01000000", -- 1973 - 0x7b5  :   64 - 0x40
    "11100000", -- 1974 - 0x7b6  :  224 - 0xe0
    "11100000", -- 1975 - 0x7b7  :  224 - 0xe0
    "01111000", -- 1976 - 0x7b8  :  120 - 0x78 -- Sprite 0xf7
    "10111100", -- 1977 - 0x7b9  :  188 - 0xbc
    "10111000", -- 1978 - 0x7ba  :  184 - 0xb8
    "10111110", -- 1979 - 0x7bb  :  190 - 0xbe
    "01111100", -- 1980 - 0x7bc  :  124 - 0x7c
    "11111110", -- 1981 - 0x7bd  :  254 - 0xfe
    "01111000", -- 1982 - 0x7be  :  120 - 0x78
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000011", -- 1984 - 0x7c0  :    3 - 0x3 -- Sprite 0xf8
    "00000011", -- 1985 - 0x7c1  :    3 - 0x3
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000011", -- 1987 - 0x7c3  :    3 - 0x3
    "00000111", -- 1988 - 0x7c4  :    7 - 0x7
    "00000110", -- 1989 - 0x7c5  :    6 - 0x6
    "00000111", -- 1990 - 0x7c6  :    7 - 0x7
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00011111", -- 1993 - 0x7c9  :   31 - 0x1f
    "00011111", -- 1994 - 0x7ca  :   31 - 0x1f
    "00001111", -- 1995 - 0x7cb  :   15 - 0xf
    "00000011", -- 1996 - 0x7cc  :    3 - 0x3
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "11100000", -- 2000 - 0x7d0  :  224 - 0xe0 -- Sprite 0xfa
    "11100000", -- 2001 - 0x7d1  :  224 - 0xe0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00110000", -- 2003 - 0x7d3  :   48 - 0x30
    "01110000", -- 2004 - 0x7d4  :  112 - 0x70
    "01100000", -- 2005 - 0x7d5  :   96 - 0x60
    "01110000", -- 2006 - 0x7d6  :  112 - 0x70
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "11111000", -- 2009 - 0x7d9  :  248 - 0xf8
    "11111000", -- 2010 - 0x7da  :  248 - 0xf8
    "11110000", -- 2011 - 0x7db  :  240 - 0xf0
    "11000000", -- 2012 - 0x7dc  :  192 - 0xc0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00111000", -- 2016 - 0x7e0  :   56 - 0x38 -- Sprite 0xfc
    "00111000", -- 2017 - 0x7e1  :   56 - 0x38
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "01111100", -- 2019 - 0x7e3  :  124 - 0x7c
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00111000", -- 2021 - 0x7e5  :   56 - 0x38
    "00111000", -- 2022 - 0x7e6  :   56 - 0x38
    "01111100", -- 2023 - 0x7e7  :  124 - 0x7c
    "01111100", -- 2024 - 0x7e8  :  124 - 0x7c -- Sprite 0xfd
    "01111100", -- 2025 - 0x7e9  :  124 - 0x7c
    "01111100", -- 2026 - 0x7ea  :  124 - 0x7c
    "00111000", -- 2027 - 0x7eb  :   56 - 0x38
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "01111100", -- 2029 - 0x7ed  :  124 - 0x7c
    "01111100", -- 2030 - 0x7ee  :  124 - 0x7c
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00010001", -- 2034 - 0x7f2  :   17 - 0x11
    "11010111", -- 2035 - 0x7f3  :  215 - 0xd7
    "11010111", -- 2036 - 0x7f4  :  215 - 0xd7
    "11010111", -- 2037 - 0x7f5  :  215 - 0xd7
    "00010001", -- 2038 - 0x7f6  :   17 - 0x11
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "11100110", -- 2042 - 0x7fa  :  230 - 0xe6
    "11110110", -- 2043 - 0x7fb  :  246 - 0xf6
    "11110110", -- 2044 - 0x7fc  :  246 - 0xf6
    "11110110", -- 2045 - 0x7fd  :  246 - 0xf6
    "11100110", -- 2046 - 0x7fe  :  230 - 0xe6
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
          -- Background pattern Table
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Background 0x0
    "01111111", -- 2049 - 0x801  :  127 - 0x7f
    "01111111", -- 2050 - 0x802  :  127 - 0x7f
    "01111111", -- 2051 - 0x803  :  127 - 0x7f
    "01111111", -- 2052 - 0x804  :  127 - 0x7f
    "01111111", -- 2053 - 0x805  :  127 - 0x7f
    "01101010", -- 2054 - 0x806  :  106 - 0x6a
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- Background 0x1
    "01111011", -- 2057 - 0x809  :  123 - 0x7b
    "01110011", -- 2058 - 0x80a  :  115 - 0x73
    "01111011", -- 2059 - 0x80b  :  123 - 0x7b
    "01110011", -- 2060 - 0x80c  :  115 - 0x73
    "01111011", -- 2061 - 0x80d  :  123 - 0x7b
    "01010011", -- 2062 - 0x80e  :   83 - 0x53
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "00000000", -- 2064 - 0x810  :    0 - 0x0 -- Background 0x2
    "11011110", -- 2065 - 0x811  :  222 - 0xde
    "10011110", -- 2066 - 0x812  :  158 - 0x9e
    "11011100", -- 2067 - 0x813  :  220 - 0xdc
    "10011110", -- 2068 - 0x814  :  158 - 0x9e
    "11011100", -- 2069 - 0x815  :  220 - 0xdc
    "10011010", -- 2070 - 0x816  :  154 - 0x9a
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- Background 0x3
    "11111110", -- 2073 - 0x819  :  254 - 0xfe
    "11111100", -- 2074 - 0x81a  :  252 - 0xfc
    "11111110", -- 2075 - 0x81b  :  254 - 0xfe
    "11111100", -- 2076 - 0x81c  :  252 - 0xfc
    "11111110", -- 2077 - 0x81d  :  254 - 0xfe
    "01010100", -- 2078 - 0x81e  :   84 - 0x54
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00000000", -- 2080 - 0x820  :    0 - 0x0 -- Background 0x4
    "01111111", -- 2081 - 0x821  :  127 - 0x7f
    "01011111", -- 2082 - 0x822  :   95 - 0x5f
    "01111001", -- 2083 - 0x823  :  121 - 0x79
    "01111001", -- 2084 - 0x824  :  121 - 0x79
    "01001001", -- 2085 - 0x825  :   73 - 0x49
    "01001111", -- 2086 - 0x826  :   79 - 0x4f
    "01001110", -- 2087 - 0x827  :   78 - 0x4e
    "01111000", -- 2088 - 0x828  :  120 - 0x78 -- Background 0x5
    "01110000", -- 2089 - 0x829  :  112 - 0x70
    "01100000", -- 2090 - 0x82a  :   96 - 0x60
    "01100000", -- 2091 - 0x82b  :   96 - 0x60
    "01110001", -- 2092 - 0x82c  :  113 - 0x71
    "01011111", -- 2093 - 0x82d  :   95 - 0x5f
    "01111111", -- 2094 - 0x82e  :  127 - 0x7f
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00000000", -- 2096 - 0x830  :    0 - 0x0 -- Background 0x6
    "11111110", -- 2097 - 0x831  :  254 - 0xfe
    "11111010", -- 2098 - 0x832  :  250 - 0xfa
    "10011110", -- 2099 - 0x833  :  158 - 0x9e
    "10011110", -- 2100 - 0x834  :  158 - 0x9e
    "10010010", -- 2101 - 0x835  :  146 - 0x92
    "11110010", -- 2102 - 0x836  :  242 - 0xf2
    "01110010", -- 2103 - 0x837  :  114 - 0x72
    "00011110", -- 2104 - 0x838  :   30 - 0x1e -- Background 0x7
    "00001110", -- 2105 - 0x839  :   14 - 0xe
    "00000110", -- 2106 - 0x83a  :    6 - 0x6
    "00000110", -- 2107 - 0x83b  :    6 - 0x6
    "10001110", -- 2108 - 0x83c  :  142 - 0x8e
    "11111010", -- 2109 - 0x83d  :  250 - 0xfa
    "11111110", -- 2110 - 0x83e  :  254 - 0xfe
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0 -- Background 0x8
    "01111111", -- 2113 - 0x841  :  127 - 0x7f
    "01011111", -- 2114 - 0x842  :   95 - 0x5f
    "01111111", -- 2115 - 0x843  :  127 - 0x7f
    "01111111", -- 2116 - 0x844  :  127 - 0x7f
    "01111111", -- 2117 - 0x845  :  127 - 0x7f
    "01111111", -- 2118 - 0x846  :  127 - 0x7f
    "01111111", -- 2119 - 0x847  :  127 - 0x7f
    "01111111", -- 2120 - 0x848  :  127 - 0x7f -- Background 0x9
    "01111111", -- 2121 - 0x849  :  127 - 0x7f
    "01111111", -- 2122 - 0x84a  :  127 - 0x7f
    "01111111", -- 2123 - 0x84b  :  127 - 0x7f
    "01111111", -- 2124 - 0x84c  :  127 - 0x7f
    "01011111", -- 2125 - 0x84d  :   95 - 0x5f
    "01111111", -- 2126 - 0x84e  :  127 - 0x7f
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00000000", -- 2128 - 0x850  :    0 - 0x0 -- Background 0xa
    "11111110", -- 2129 - 0x851  :  254 - 0xfe
    "11111010", -- 2130 - 0x852  :  250 - 0xfa
    "11111110", -- 2131 - 0x853  :  254 - 0xfe
    "11111110", -- 2132 - 0x854  :  254 - 0xfe
    "11111110", -- 2133 - 0x855  :  254 - 0xfe
    "11111110", -- 2134 - 0x856  :  254 - 0xfe
    "11111110", -- 2135 - 0x857  :  254 - 0xfe
    "11111110", -- 2136 - 0x858  :  254 - 0xfe -- Background 0xb
    "11111110", -- 2137 - 0x859  :  254 - 0xfe
    "11111110", -- 2138 - 0x85a  :  254 - 0xfe
    "11111110", -- 2139 - 0x85b  :  254 - 0xfe
    "11111110", -- 2140 - 0x85c  :  254 - 0xfe
    "11111010", -- 2141 - 0x85d  :  250 - 0xfa
    "11111110", -- 2142 - 0x85e  :  254 - 0xfe
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Background 0xc
    "00111111", -- 2145 - 0x861  :   63 - 0x3f
    "01011111", -- 2146 - 0x862  :   95 - 0x5f
    "01101111", -- 2147 - 0x863  :  111 - 0x6f
    "01110000", -- 2148 - 0x864  :  112 - 0x70
    "01110111", -- 2149 - 0x865  :  119 - 0x77
    "01110111", -- 2150 - 0x866  :  119 - 0x77
    "01110111", -- 2151 - 0x867  :  119 - 0x77
    "01110111", -- 2152 - 0x868  :  119 - 0x77 -- Background 0xd
    "01110111", -- 2153 - 0x869  :  119 - 0x77
    "01110111", -- 2154 - 0x86a  :  119 - 0x77
    "01110000", -- 2155 - 0x86b  :  112 - 0x70
    "01101111", -- 2156 - 0x86c  :  111 - 0x6f
    "01011111", -- 2157 - 0x86d  :   95 - 0x5f
    "00010101", -- 2158 - 0x86e  :   21 - 0x15
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0 -- Background 0xe
    "11111100", -- 2161 - 0x871  :  252 - 0xfc
    "11111000", -- 2162 - 0x872  :  248 - 0xf8
    "11110110", -- 2163 - 0x873  :  246 - 0xf6
    "00001100", -- 2164 - 0x874  :   12 - 0xc
    "11101110", -- 2165 - 0x875  :  238 - 0xee
    "11101100", -- 2166 - 0x876  :  236 - 0xec
    "11101110", -- 2167 - 0x877  :  238 - 0xee
    "11101100", -- 2168 - 0x878  :  236 - 0xec -- Background 0xf
    "11101110", -- 2169 - 0x879  :  238 - 0xee
    "11101100", -- 2170 - 0x87a  :  236 - 0xec
    "00001110", -- 2171 - 0x87b  :   14 - 0xe
    "11110100", -- 2172 - 0x87c  :  244 - 0xf4
    "11111010", -- 2173 - 0x87d  :  250 - 0xfa
    "01010100", -- 2174 - 0x87e  :   84 - 0x54
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "01100000", -- 2176 - 0x880  :   96 - 0x60 -- Background 0x10
    "01100000", -- 2177 - 0x881  :   96 - 0x60
    "01100000", -- 2178 - 0x882  :   96 - 0x60
    "01101111", -- 2179 - 0x883  :  111 - 0x6f
    "01101010", -- 2180 - 0x884  :  106 - 0x6a
    "01100000", -- 2181 - 0x885  :   96 - 0x60
    "01100000", -- 2182 - 0x886  :   96 - 0x60
    "01100000", -- 2183 - 0x887  :   96 - 0x60
    "00000110", -- 2184 - 0x888  :    6 - 0x6 -- Background 0x11
    "00000100", -- 2185 - 0x889  :    4 - 0x4
    "00000110", -- 2186 - 0x88a  :    6 - 0x6
    "11110100", -- 2187 - 0x88b  :  244 - 0xf4
    "10100110", -- 2188 - 0x88c  :  166 - 0xa6
    "00000100", -- 2189 - 0x88d  :    4 - 0x4
    "00000110", -- 2190 - 0x88e  :    6 - 0x6
    "00000100", -- 2191 - 0x88f  :    4 - 0x4
    "00000000", -- 2192 - 0x890  :    0 - 0x0 -- Background 0x12
    "00001000", -- 2193 - 0x891  :    8 - 0x8
    "00001000", -- 2194 - 0x892  :    8 - 0x8
    "00011100", -- 2195 - 0x893  :   28 - 0x1c
    "00011100", -- 2196 - 0x894  :   28 - 0x1c
    "00111100", -- 2197 - 0x895  :   60 - 0x3c
    "00111100", -- 2198 - 0x896  :   60 - 0x3c
    "00111100", -- 2199 - 0x897  :   60 - 0x3c
    "00111100", -- 2200 - 0x898  :   60 - 0x3c -- Background 0x13
    "01111110", -- 2201 - 0x899  :  126 - 0x7e
    "01111110", -- 2202 - 0x89a  :  126 - 0x7e
    "01111110", -- 2203 - 0x89b  :  126 - 0x7e
    "01111110", -- 2204 - 0x89c  :  126 - 0x7e
    "01111110", -- 2205 - 0x89d  :  126 - 0x7e
    "01111110", -- 2206 - 0x89e  :  126 - 0x7e
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x14
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000101", -- 2210 - 0x8a2  :    5 - 0x5
    "00000011", -- 2211 - 0x8a3  :    3 - 0x3
    "00000000", -- 2212 - 0x8a4  :    0 - 0x0
    "00000000", -- 2213 - 0x8a5  :    0 - 0x0
    "00000010", -- 2214 - 0x8a6  :    2 - 0x2
    "00001111", -- 2215 - 0x8a7  :   15 - 0xf
    "00011100", -- 2216 - 0x8a8  :   28 - 0x1c -- Background 0x15
    "00111010", -- 2217 - 0x8a9  :   58 - 0x3a
    "00111100", -- 2218 - 0x8aa  :   60 - 0x3c
    "00111111", -- 2219 - 0x8ab  :   63 - 0x3f
    "00111000", -- 2220 - 0x8ac  :   56 - 0x38
    "00011110", -- 2221 - 0x8ad  :   30 - 0x1e
    "00001111", -- 2222 - 0x8ae  :   15 - 0xf
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "00000000", -- 2224 - 0x8b0  :    0 - 0x0 -- Background 0x16
    "00000000", -- 2225 - 0x8b1  :    0 - 0x0
    "01000000", -- 2226 - 0x8b2  :   64 - 0x40
    "11000000", -- 2227 - 0x8b3  :  192 - 0xc0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "10000000", -- 2229 - 0x8b5  :  128 - 0x80
    "11000000", -- 2230 - 0x8b6  :  192 - 0xc0
    "01110000", -- 2231 - 0x8b7  :  112 - 0x70
    "00011000", -- 2232 - 0x8b8  :   24 - 0x18 -- Background 0x17
    "11111100", -- 2233 - 0x8b9  :  252 - 0xfc
    "00111100", -- 2234 - 0x8ba  :   60 - 0x3c
    "01011100", -- 2235 - 0x8bb  :   92 - 0x5c
    "00111100", -- 2236 - 0x8bc  :   60 - 0x3c
    "11111000", -- 2237 - 0x8bd  :  248 - 0xf8
    "11110000", -- 2238 - 0x8be  :  240 - 0xf0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Background 0x18
    "00111111", -- 2241 - 0x8c1  :   63 - 0x3f
    "00111111", -- 2242 - 0x8c2  :   63 - 0x3f
    "01111111", -- 2243 - 0x8c3  :  127 - 0x7f
    "01111111", -- 2244 - 0x8c4  :  127 - 0x7f
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "00000000", -- 2246 - 0x8c6  :    0 - 0x0
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- Background 0x19
    "11111100", -- 2249 - 0x8c9  :  252 - 0xfc
    "11111100", -- 2250 - 0x8ca  :  252 - 0xfc
    "11111110", -- 2251 - 0x8cb  :  254 - 0xfe
    "11111110", -- 2252 - 0x8cc  :  254 - 0xfe
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "00000000", -- 2256 - 0x8d0  :    0 - 0x0 -- Background 0x1a
    "00000000", -- 2257 - 0x8d1  :    0 - 0x0
    "00000000", -- 2258 - 0x8d2  :    0 - 0x0
    "00111111", -- 2259 - 0x8d3  :   63 - 0x3f
    "00111111", -- 2260 - 0x8d4  :   63 - 0x3f
    "01111111", -- 2261 - 0x8d5  :  127 - 0x7f
    "01111111", -- 2262 - 0x8d6  :  127 - 0x7f
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- Background 0x1b
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "11111100", -- 2267 - 0x8db  :  252 - 0xfc
    "11111100", -- 2268 - 0x8dc  :  252 - 0xfc
    "11111110", -- 2269 - 0x8dd  :  254 - 0xfe
    "11111110", -- 2270 - 0x8de  :  254 - 0xfe
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Background 0x1c
    "01111111", -- 2273 - 0x8e1  :  127 - 0x7f
    "01111111", -- 2274 - 0x8e2  :  127 - 0x7f
    "01111111", -- 2275 - 0x8e3  :  127 - 0x7f
    "01100100", -- 2276 - 0x8e4  :  100 - 0x64
    "01011011", -- 2277 - 0x8e5  :   91 - 0x5b
    "01011001", -- 2278 - 0x8e6  :   89 - 0x59
    "01111111", -- 2279 - 0x8e7  :  127 - 0x7f
    "01111111", -- 2280 - 0x8e8  :  127 - 0x7f -- Background 0x1d
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000001", -- 2282 - 0x8ea  :    1 - 0x1
    "00000001", -- 2283 - 0x8eb  :    1 - 0x1
    "00000001", -- 2284 - 0x8ec  :    1 - 0x1
    "00000001", -- 2285 - 0x8ed  :    1 - 0x1
    "00000001", -- 2286 - 0x8ee  :    1 - 0x1
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "00000000", -- 2288 - 0x8f0  :    0 - 0x0 -- Background 0x1e
    "11111110", -- 2289 - 0x8f1  :  254 - 0xfe
    "11111110", -- 2290 - 0x8f2  :  254 - 0xfe
    "11111110", -- 2291 - 0x8f3  :  254 - 0xfe
    "10111110", -- 2292 - 0x8f4  :  190 - 0xbe
    "00001010", -- 2293 - 0x8f5  :   10 - 0xa
    "11100010", -- 2294 - 0x8f6  :  226 - 0xe2
    "11111110", -- 2295 - 0x8f7  :  254 - 0xfe
    "11111110", -- 2296 - 0x8f8  :  254 - 0xfe -- Background 0x1f
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "10000000", -- 2298 - 0x8fa  :  128 - 0x80
    "10000000", -- 2299 - 0x8fb  :  128 - 0x80
    "10000000", -- 2300 - 0x8fc  :  128 - 0x80
    "10000000", -- 2301 - 0x8fd  :  128 - 0x80
    "10000000", -- 2302 - 0x8fe  :  128 - 0x80
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x20
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000000", -- 2308 - 0x904  :    0 - 0x0
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "00000000", -- 2310 - 0x906  :    0 - 0x0
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- Background 0x21
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00000000", -- 2316 - 0x90c  :    0 - 0x0
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "00000000", -- 2318 - 0x90e  :    0 - 0x0
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "00000000", -- 2320 - 0x910  :    0 - 0x0 -- Background 0x22
    "00000000", -- 2321 - 0x911  :    0 - 0x0
    "00011000", -- 2322 - 0x912  :   24 - 0x18
    "00010000", -- 2323 - 0x913  :   16 - 0x10
    "00011010", -- 2324 - 0x914  :   26 - 0x1a
    "00010001", -- 2325 - 0x915  :   17 - 0x11
    "00011010", -- 2326 - 0x916  :   26 - 0x1a
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "00000000", -- 2328 - 0x918  :    0 - 0x0 -- Background 0x23
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00101000", -- 2331 - 0x91b  :   40 - 0x28
    "10001100", -- 2332 - 0x91c  :  140 - 0x8c
    "00101000", -- 2333 - 0x91d  :   40 - 0x28
    "10101100", -- 2334 - 0x91e  :  172 - 0xac
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Background 0x24
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00011100", -- 2344 - 0x928  :   28 - 0x1c -- Background 0x25
    "00111001", -- 2345 - 0x929  :   57 - 0x39
    "00111111", -- 2346 - 0x92a  :   63 - 0x3f
    "00111110", -- 2347 - 0x92b  :   62 - 0x3e
    "00111111", -- 2348 - 0x92c  :   63 - 0x3f
    "00011110", -- 2349 - 0x92d  :   30 - 0x1e
    "00001111", -- 2350 - 0x92e  :   15 - 0xf
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "00000000", -- 2353 - 0x931  :    0 - 0x0
    "01000000", -- 2354 - 0x932  :   64 - 0x40
    "11000000", -- 2355 - 0x933  :  192 - 0xc0
    "00000000", -- 2356 - 0x934  :    0 - 0x0
    "10000000", -- 2357 - 0x935  :  128 - 0x80
    "11000000", -- 2358 - 0x936  :  192 - 0xc0
    "11110000", -- 2359 - 0x937  :  240 - 0xf0
    "00111000", -- 2360 - 0x938  :   56 - 0x38 -- Background 0x27
    "10011100", -- 2361 - 0x939  :  156 - 0x9c
    "10011100", -- 2362 - 0x93a  :  156 - 0x9c
    "00111100", -- 2363 - 0x93b  :   60 - 0x3c
    "11111100", -- 2364 - 0x93c  :  252 - 0xfc
    "01111000", -- 2365 - 0x93d  :  120 - 0x78
    "11110000", -- 2366 - 0x93e  :  240 - 0xf0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "00111110", -- 2369 - 0x941  :   62 - 0x3e
    "01011101", -- 2370 - 0x942  :   93 - 0x5d
    "01101011", -- 2371 - 0x943  :  107 - 0x6b
    "01110101", -- 2372 - 0x944  :  117 - 0x75
    "01110001", -- 2373 - 0x945  :  113 - 0x71
    "01110101", -- 2374 - 0x946  :  117 - 0x75
    "01110100", -- 2375 - 0x947  :  116 - 0x74
    "01110000", -- 2376 - 0x948  :  112 - 0x70 -- Background 0x29
    "01110111", -- 2377 - 0x949  :  119 - 0x77
    "01110111", -- 2378 - 0x94a  :  119 - 0x77
    "01110000", -- 2379 - 0x94b  :  112 - 0x70
    "01101111", -- 2380 - 0x94c  :  111 - 0x6f
    "01011111", -- 2381 - 0x94d  :   95 - 0x5f
    "00010101", -- 2382 - 0x94e  :   21 - 0x15
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00000000", -- 2384 - 0x950  :    0 - 0x0 -- Background 0x2a
    "01111100", -- 2385 - 0x951  :  124 - 0x7c
    "10111000", -- 2386 - 0x952  :  184 - 0xb8
    "11010110", -- 2387 - 0x953  :  214 - 0xd6
    "10101100", -- 2388 - 0x954  :  172 - 0xac
    "10001110", -- 2389 - 0x955  :  142 - 0x8e
    "10101100", -- 2390 - 0x956  :  172 - 0xac
    "00101110", -- 2391 - 0x957  :   46 - 0x2e
    "00001100", -- 2392 - 0x958  :   12 - 0xc -- Background 0x2b
    "11101110", -- 2393 - 0x959  :  238 - 0xee
    "11101100", -- 2394 - 0x95a  :  236 - 0xec
    "00001110", -- 2395 - 0x95b  :   14 - 0xe
    "11110100", -- 2396 - 0x95c  :  244 - 0xf4
    "11111010", -- 2397 - 0x95d  :  250 - 0xfa
    "01010100", -- 2398 - 0x95e  :   84 - 0x54
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00011110", -- 2408 - 0x968  :   30 - 0x1e -- Background 0x2d
    "00111110", -- 2409 - 0x969  :   62 - 0x3e
    "00111110", -- 2410 - 0x96a  :   62 - 0x3e
    "00111110", -- 2411 - 0x96b  :   62 - 0x3e
    "00111111", -- 2412 - 0x96c  :   63 - 0x3f
    "00011110", -- 2413 - 0x96d  :   30 - 0x1e
    "00001111", -- 2414 - 0x96e  :   15 - 0xf
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "01111000", -- 2424 - 0x978  :  120 - 0x78 -- Background 0x2f
    "01111100", -- 2425 - 0x979  :  124 - 0x7c
    "01111100", -- 2426 - 0x97a  :  124 - 0x7c
    "01111100", -- 2427 - 0x97b  :  124 - 0x7c
    "11111100", -- 2428 - 0x97c  :  252 - 0xfc
    "01111000", -- 2429 - 0x97d  :  120 - 0x78
    "11110000", -- 2430 - 0x97e  :  240 - 0xf0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Background 0x30
    "00011000", -- 2433 - 0x981  :   24 - 0x18
    "00111100", -- 2434 - 0x982  :   60 - 0x3c
    "01011010", -- 2435 - 0x983  :   90 - 0x5a
    "00011000", -- 2436 - 0x984  :   24 - 0x18
    "00011000", -- 2437 - 0x985  :   24 - 0x18
    "00011000", -- 2438 - 0x986  :   24 - 0x18
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- Background 0x31
    "00011000", -- 2441 - 0x989  :   24 - 0x18
    "00011000", -- 2442 - 0x98a  :   24 - 0x18
    "00011000", -- 2443 - 0x98b  :   24 - 0x18
    "01011010", -- 2444 - 0x98c  :   90 - 0x5a
    "00111100", -- 2445 - 0x98d  :   60 - 0x3c
    "00011000", -- 2446 - 0x98e  :   24 - 0x18
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000001", -- 2448 - 0x990  :    1 - 0x1 -- Background 0x32
    "00000001", -- 2449 - 0x991  :    1 - 0x1
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000001", -- 2451 - 0x993  :    1 - 0x1
    "00000001", -- 2452 - 0x994  :    1 - 0x1
    "00000001", -- 2453 - 0x995  :    1 - 0x1
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000001", -- 2455 - 0x997  :    1 - 0x1
    "10000000", -- 2456 - 0x998  :  128 - 0x80 -- Background 0x33
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "10000000", -- 2458 - 0x99a  :  128 - 0x80
    "10000000", -- 2459 - 0x99b  :  128 - 0x80
    "10000000", -- 2460 - 0x99c  :  128 - 0x80
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "10000000", -- 2462 - 0x99e  :  128 - 0x80
    "10000000", -- 2463 - 0x99f  :  128 - 0x80
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Background 0x34
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00011000", -- 2466 - 0x9a2  :   24 - 0x18
    "00111100", -- 2467 - 0x9a3  :   60 - 0x3c
    "00111110", -- 2468 - 0x9a4  :   62 - 0x3e
    "01111111", -- 2469 - 0x9a5  :  127 - 0x7f
    "01111111", -- 2470 - 0x9a6  :  127 - 0x7f
    "01111111", -- 2471 - 0x9a7  :  127 - 0x7f
    "00111111", -- 2472 - 0x9a8  :   63 - 0x3f -- Background 0x35
    "00111111", -- 2473 - 0x9a9  :   63 - 0x3f
    "00011111", -- 2474 - 0x9aa  :   31 - 0x1f
    "00001111", -- 2475 - 0x9ab  :   15 - 0xf
    "00000111", -- 2476 - 0x9ac  :    7 - 0x7
    "00000011", -- 2477 - 0x9ad  :    3 - 0x3
    "00000001", -- 2478 - 0x9ae  :    1 - 0x1
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0 -- Background 0x36
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00011000", -- 2482 - 0x9b2  :   24 - 0x18
    "00111100", -- 2483 - 0x9b3  :   60 - 0x3c
    "01111100", -- 2484 - 0x9b4  :  124 - 0x7c
    "11111110", -- 2485 - 0x9b5  :  254 - 0xfe
    "11111110", -- 2486 - 0x9b6  :  254 - 0xfe
    "11111110", -- 2487 - 0x9b7  :  254 - 0xfe
    "11111100", -- 2488 - 0x9b8  :  252 - 0xfc -- Background 0x37
    "11111100", -- 2489 - 0x9b9  :  252 - 0xfc
    "11111000", -- 2490 - 0x9ba  :  248 - 0xf8
    "11110000", -- 2491 - 0x9bb  :  240 - 0xf0
    "11100000", -- 2492 - 0x9bc  :  224 - 0xe0
    "11000000", -- 2493 - 0x9bd  :  192 - 0xc0
    "10000000", -- 2494 - 0x9be  :  128 - 0x80
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000110", -- 2498 - 0x9c2  :    6 - 0x6
    "00000111", -- 2499 - 0x9c3  :    7 - 0x7
    "00000111", -- 2500 - 0x9c4  :    7 - 0x7
    "00000011", -- 2501 - 0x9c5  :    3 - 0x3
    "00000001", -- 2502 - 0x9c6  :    1 - 0x1
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "01100000", -- 2514 - 0x9d2  :   96 - 0x60
    "11100000", -- 2515 - 0x9d3  :  224 - 0xe0
    "11100000", -- 2516 - 0x9d4  :  224 - 0xe0
    "11000000", -- 2517 - 0x9d5  :  192 - 0xc0
    "10000000", -- 2518 - 0x9d6  :  128 - 0x80
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00101010", -- 2521 - 0x9d9  :   42 - 0x2a
    "01000000", -- 2522 - 0x9da  :   64 - 0x40
    "00000010", -- 2523 - 0x9db  :    2 - 0x2
    "01000000", -- 2524 - 0x9dc  :   64 - 0x40
    "00000010", -- 2525 - 0x9dd  :    2 - 0x2
    "01010100", -- 2526 - 0x9de  :   84 - 0x54
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "11111111", -- 2536 - 0x9e8  :  255 - 0xff -- Background 0x3d
    "11111111", -- 2537 - 0x9e9  :  255 - 0xff
    "11111111", -- 2538 - 0x9ea  :  255 - 0xff
    "11111111", -- 2539 - 0x9eb  :  255 - 0xff
    "11111111", -- 2540 - 0x9ec  :  255 - 0xff
    "11111111", -- 2541 - 0x9ed  :  255 - 0xff
    "11111111", -- 2542 - 0x9ee  :  255 - 0xff
    "11111111", -- 2543 - 0x9ef  :  255 - 0xff
    "11111111", -- 2544 - 0x9f0  :  255 - 0xff -- Background 0x3e
    "11111111", -- 2545 - 0x9f1  :  255 - 0xff
    "11111111", -- 2546 - 0x9f2  :  255 - 0xff
    "11111111", -- 2547 - 0x9f3  :  255 - 0xff
    "11111111", -- 2548 - 0x9f4  :  255 - 0xff
    "11111111", -- 2549 - 0x9f5  :  255 - 0xff
    "11111111", -- 2550 - 0x9f6  :  255 - 0xff
    "11111111", -- 2551 - 0x9f7  :  255 - 0xff
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Background 0x40
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- Background 0x41
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Background 0x42
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "00000000", -- 2580 - 0xa14  :    0 - 0x0
    "00000000", -- 2581 - 0xa15  :    0 - 0x0
    "00000000", -- 2582 - 0xa16  :    0 - 0x0
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00000000", -- 2584 - 0xa18  :    0 - 0x0 -- Background 0x43
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Background 0x44
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "00000000", -- 2594 - 0xa22  :    0 - 0x0
    "00000000", -- 2595 - 0xa23  :    0 - 0x0
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "00000000", -- 2598 - 0xa26  :    0 - 0x0
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- Background 0x45
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00000000", -- 2608 - 0xa30  :    0 - 0x0 -- Background 0x46
    "00000000", -- 2609 - 0xa31  :    0 - 0x0
    "00000000", -- 2610 - 0xa32  :    0 - 0x0
    "00000000", -- 2611 - 0xa33  :    0 - 0x0
    "00000000", -- 2612 - 0xa34  :    0 - 0x0
    "00000000", -- 2613 - 0xa35  :    0 - 0x0
    "00000000", -- 2614 - 0xa36  :    0 - 0x0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- Background 0x47
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0x48
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- Background 0x49
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "00000000", -- 2648 - 0xa58  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00000000", -- 2658 - 0xa62  :    0 - 0x0
    "00000000", -- 2659 - 0xa63  :    0 - 0x0
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0 -- Background 0x4e
    "00000000", -- 2673 - 0xa71  :    0 - 0x0
    "00000000", -- 2674 - 0xa72  :    0 - 0x0
    "00000000", -- 2675 - 0xa73  :    0 - 0x0
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "00000000", -- 2677 - 0xa75  :    0 - 0x0
    "00000000", -- 2678 - 0xa76  :    0 - 0x0
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00000000", -- 2680 - 0xa78  :    0 - 0x0 -- Background 0x4f
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000000", -- 2685 - 0xa7d  :    0 - 0x0
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Background 0x50
    "00111111", -- 2689 - 0xa81  :   63 - 0x3f
    "01111111", -- 2690 - 0xa82  :  127 - 0x7f
    "01111111", -- 2691 - 0xa83  :  127 - 0x7f
    "01111111", -- 2692 - 0xa84  :  127 - 0x7f
    "00111100", -- 2693 - 0xa85  :   60 - 0x3c
    "00000000", -- 2694 - 0xa86  :    0 - 0x0
    "01000000", -- 2695 - 0xa87  :   64 - 0x40
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- Background 0x51
    "11111100", -- 2697 - 0xa89  :  252 - 0xfc
    "11111110", -- 2698 - 0xa8a  :  254 - 0xfe
    "11111110", -- 2699 - 0xa8b  :  254 - 0xfe
    "11111110", -- 2700 - 0xa8c  :  254 - 0xfe
    "00111100", -- 2701 - 0xa8d  :   60 - 0x3c
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000010", -- 2703 - 0xa8f  :    2 - 0x2
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00000011", -- 2706 - 0xa92  :    3 - 0x3
    "00000111", -- 2707 - 0xa93  :    7 - 0x7
    "00001111", -- 2708 - 0xa94  :   15 - 0xf
    "00011111", -- 2709 - 0xa95  :   31 - 0x1f
    "00111111", -- 2710 - 0xa96  :   63 - 0x3f
    "00110000", -- 2711 - 0xa97  :   48 - 0x30
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- Background 0x53
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "10100000", -- 2714 - 0xa9a  :  160 - 0xa0
    "10110000", -- 2715 - 0xa9b  :  176 - 0xb0
    "10110000", -- 2716 - 0xa9c  :  176 - 0xb0
    "10111000", -- 2717 - 0xa9d  :  184 - 0xb8
    "01111100", -- 2718 - 0xa9e  :  124 - 0x7c
    "01111100", -- 2719 - 0xa9f  :  124 - 0x7c
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Background 0x54
    "00100001", -- 2721 - 0xaa1  :   33 - 0x21
    "01110001", -- 2722 - 0xaa2  :  113 - 0x71
    "00111010", -- 2723 - 0xaa3  :   58 - 0x3a
    "01101101", -- 2724 - 0xaa4  :  109 - 0x6d
    "00111000", -- 2725 - 0xaa5  :   56 - 0x38
    "00011101", -- 2726 - 0xaa6  :   29 - 0x1d
    "00101111", -- 2727 - 0xaa7  :   47 - 0x2f
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- Background 0x55
    "00100001", -- 2729 - 0xaa9  :   33 - 0x21
    "01110001", -- 2730 - 0xaaa  :  113 - 0x71
    "00111010", -- 2731 - 0xaab  :   58 - 0x3a
    "01101101", -- 2732 - 0xaac  :  109 - 0x6d
    "10111000", -- 2733 - 0xaad  :  184 - 0xb8
    "00011101", -- 2734 - 0xaae  :   29 - 0x1d
    "10101111", -- 2735 - 0xaaf  :  175 - 0xaf
    "00000000", -- 2736 - 0xab0  :    0 - 0x0 -- Background 0x56
    "00100000", -- 2737 - 0xab1  :   32 - 0x20
    "01110000", -- 2738 - 0xab2  :  112 - 0x70
    "00111010", -- 2739 - 0xab3  :   58 - 0x3a
    "01101100", -- 2740 - 0xab4  :  108 - 0x6c
    "10111000", -- 2741 - 0xab5  :  184 - 0xb8
    "00011100", -- 2742 - 0xab6  :   28 - 0x1c
    "10101110", -- 2743 - 0xab7  :  174 - 0xae
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- Background 0x57
    "01111111", -- 2745 - 0xab9  :  127 - 0x7f
    "01001100", -- 2746 - 0xaba  :   76 - 0x4c
    "00110011", -- 2747 - 0xabb  :   51 - 0x33
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Background 0x58
    "11111111", -- 2753 - 0xac1  :  255 - 0xff
    "11001100", -- 2754 - 0xac2  :  204 - 0xcc
    "00110011", -- 2755 - 0xac3  :   51 - 0x33
    "11001100", -- 2756 - 0xac4  :  204 - 0xcc
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- Background 0x59
    "11111110", -- 2761 - 0xac9  :  254 - 0xfe
    "11001100", -- 2762 - 0xaca  :  204 - 0xcc
    "00110000", -- 2763 - 0xacb  :   48 - 0x30
    "11000000", -- 2764 - 0xacc  :  192 - 0xc0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "00000000", -- 2771 - 0xad3  :    0 - 0x0
    "00000000", -- 2772 - 0xad4  :    0 - 0x0
    "00000000", -- 2773 - 0xad5  :    0 - 0x0
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000001", -- 2780 - 0xadc  :    1 - 0x1
    "00000001", -- 2781 - 0xadd  :    1 - 0x1
    "00000011", -- 2782 - 0xade  :    3 - 0x3
    "00000011", -- 2783 - 0xadf  :    3 - 0x3
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000001", -- 2786 - 0xae2  :    1 - 0x1
    "01111110", -- 2787 - 0xae3  :  126 - 0x7e
    "11111111", -- 2788 - 0xae4  :  255 - 0xff
    "11111111", -- 2789 - 0xae5  :  255 - 0xff
    "11111111", -- 2790 - 0xae6  :  255 - 0xff
    "11111111", -- 2791 - 0xae7  :  255 - 0xff
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- Background 0x5d
    "11111111", -- 2793 - 0xae9  :  255 - 0xff
    "11111111", -- 2794 - 0xaea  :  255 - 0xff
    "11111111", -- 2795 - 0xaeb  :  255 - 0xff
    "01111111", -- 2796 - 0xaec  :  127 - 0x7f
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "11111111", -- 2798 - 0xaee  :  255 - 0xff
    "11111111", -- 2799 - 0xaef  :  255 - 0xff
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0x5e
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "10000000", -- 2802 - 0xaf2  :  128 - 0x80
    "01111110", -- 2803 - 0xaf3  :  126 - 0x7e
    "10111111", -- 2804 - 0xaf4  :  191 - 0xbf
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111111", -- 2806 - 0xaf6  :  255 - 0xff
    "11111111", -- 2807 - 0xaf7  :  255 - 0xff
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "10000000", -- 2812 - 0xafc  :  128 - 0x80
    "10000000", -- 2813 - 0xafd  :  128 - 0x80
    "11000000", -- 2814 - 0xafe  :  192 - 0xc0
    "11000000", -- 2815 - 0xaff  :  192 - 0xc0
    "01111111", -- 2816 - 0xb00  :  127 - 0x7f -- Background 0x60
    "01111111", -- 2817 - 0xb01  :  127 - 0x7f
    "01111101", -- 2818 - 0xb02  :  125 - 0x7d
    "01111111", -- 2819 - 0xb03  :  127 - 0x7f
    "00111111", -- 2820 - 0xb04  :   63 - 0x3f
    "01111111", -- 2821 - 0xb05  :  127 - 0x7f
    "01111111", -- 2822 - 0xb06  :  127 - 0x7f
    "01110111", -- 2823 - 0xb07  :  119 - 0x77
    "11111110", -- 2824 - 0xb08  :  254 - 0xfe -- Background 0x61
    "11111110", -- 2825 - 0xb09  :  254 - 0xfe
    "11111100", -- 2826 - 0xb0a  :  252 - 0xfc
    "11111110", -- 2827 - 0xb0b  :  254 - 0xfe
    "10111110", -- 2828 - 0xb0c  :  190 - 0xbe
    "11111110", -- 2829 - 0xb0d  :  254 - 0xfe
    "11111110", -- 2830 - 0xb0e  :  254 - 0xfe
    "11110110", -- 2831 - 0xb0f  :  246 - 0xf6
    "00000111", -- 2832 - 0xb10  :    7 - 0x7 -- Background 0x62
    "00011111", -- 2833 - 0xb11  :   31 - 0x1f
    "00111111", -- 2834 - 0xb12  :   63 - 0x3f
    "00111111", -- 2835 - 0xb13  :   63 - 0x3f
    "00111111", -- 2836 - 0xb14  :   63 - 0x3f
    "00011111", -- 2837 - 0xb15  :   31 - 0x1f
    "00001111", -- 2838 - 0xb16  :   15 - 0xf
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "01111110", -- 2840 - 0xb18  :  126 - 0x7e -- Background 0x63
    "01111100", -- 2841 - 0xb19  :  124 - 0x7c
    "00111110", -- 2842 - 0xb1a  :   62 - 0x3e
    "10111100", -- 2843 - 0xb1b  :  188 - 0xbc
    "10111110", -- 2844 - 0xb1c  :  190 - 0xbe
    "10011100", -- 2845 - 0xb1d  :  156 - 0x9c
    "11011000", -- 2846 - 0xb1e  :  216 - 0xd8
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "01000110", -- 2848 - 0xb20  :   70 - 0x46 -- Background 0x64
    "01101011", -- 2849 - 0xb21  :  107 - 0x6b
    "01110001", -- 2850 - 0xb22  :  113 - 0x71
    "00111010", -- 2851 - 0xb23  :   58 - 0x3a
    "01101101", -- 2852 - 0xb24  :  109 - 0x6d
    "00111000", -- 2853 - 0xb25  :   56 - 0x38
    "00011101", -- 2854 - 0xb26  :   29 - 0x1d
    "00101111", -- 2855 - 0xb27  :   47 - 0x2f
    "01000110", -- 2856 - 0xb28  :   70 - 0x46 -- Background 0x65
    "11101011", -- 2857 - 0xb29  :  235 - 0xeb
    "01110001", -- 2858 - 0xb2a  :  113 - 0x71
    "00111010", -- 2859 - 0xb2b  :   58 - 0x3a
    "01101101", -- 2860 - 0xb2c  :  109 - 0x6d
    "10111000", -- 2861 - 0xb2d  :  184 - 0xb8
    "00011101", -- 2862 - 0xb2e  :   29 - 0x1d
    "10101111", -- 2863 - 0xb2f  :  175 - 0xaf
    "01000110", -- 2864 - 0xb30  :   70 - 0x46 -- Background 0x66
    "11101010", -- 2865 - 0xb31  :  234 - 0xea
    "01110000", -- 2866 - 0xb32  :  112 - 0x70
    "00111010", -- 2867 - 0xb33  :   58 - 0x3a
    "01101100", -- 2868 - 0xb34  :  108 - 0x6c
    "10111000", -- 2869 - 0xb35  :  184 - 0xb8
    "00011100", -- 2870 - 0xb36  :   28 - 0x1c
    "10101110", -- 2871 - 0xb37  :  174 - 0xae
    "00000000", -- 2872 - 0xb38  :    0 - 0x0 -- Background 0x67
    "01111111", -- 2873 - 0xb39  :  127 - 0x7f
    "01111111", -- 2874 - 0xb3a  :  127 - 0x7f
    "00110011", -- 2875 - 0xb3b  :   51 - 0x33
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Background 0x68
    "11111111", -- 2881 - 0xb41  :  255 - 0xff
    "11111111", -- 2882 - 0xb42  :  255 - 0xff
    "11111111", -- 2883 - 0xb43  :  255 - 0xff
    "11001100", -- 2884 - 0xb44  :  204 - 0xcc
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- Background 0x69
    "11111110", -- 2889 - 0xb49  :  254 - 0xfe
    "11111110", -- 2890 - 0xb4a  :  254 - 0xfe
    "11110000", -- 2891 - 0xb4b  :  240 - 0xf0
    "11000000", -- 2892 - 0xb4c  :  192 - 0xc0
    "00000000", -- 2893 - 0xb4d  :    0 - 0x0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00111101", -- 2904 - 0xb58  :   61 - 0x3d -- Background 0x6b
    "01111111", -- 2905 - 0xb59  :  127 - 0x7f
    "01111111", -- 2906 - 0xb5a  :  127 - 0x7f
    "01111111", -- 2907 - 0xb5b  :  127 - 0x7f
    "00111111", -- 2908 - 0xb5c  :   63 - 0x3f
    "00001111", -- 2909 - 0xb5d  :   15 - 0xf
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Background 0x6c
    "11111111", -- 2913 - 0xb61  :  255 - 0xff
    "11111111", -- 2914 - 0xb62  :  255 - 0xff
    "11111111", -- 2915 - 0xb63  :  255 - 0xff
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11111111", -- 2917 - 0xb65  :  255 - 0xff
    "11111110", -- 2918 - 0xb66  :  254 - 0xfe
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "10111000", -- 2936 - 0xb78  :  184 - 0xb8 -- Background 0x6f
    "11111100", -- 2937 - 0xb79  :  252 - 0xfc
    "11111110", -- 2938 - 0xb7a  :  254 - 0xfe
    "11111110", -- 2939 - 0xb7b  :  254 - 0xfe
    "11111100", -- 2940 - 0xb7c  :  252 - 0xfc
    "11110000", -- 2941 - 0xb7d  :  240 - 0xf0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0x70
    "00111111", -- 2945 - 0xb81  :   63 - 0x3f
    "01111111", -- 2946 - 0xb82  :  127 - 0x7f
    "01111111", -- 2947 - 0xb83  :  127 - 0x7f
    "00011100", -- 2948 - 0xb84  :   28 - 0x1c
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- Background 0x71
    "11111111", -- 2953 - 0xb89  :  255 - 0xff
    "11111111", -- 2954 - 0xb8a  :  255 - 0xff
    "11111111", -- 2955 - 0xb8b  :  255 - 0xff
    "11111111", -- 2956 - 0xb8c  :  255 - 0xff
    "00111100", -- 2957 - 0xb8d  :   60 - 0x3c
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Background 0x72
    "11111100", -- 2961 - 0xb91  :  252 - 0xfc
    "11111110", -- 2962 - 0xb92  :  254 - 0xfe
    "11111110", -- 2963 - 0xb93  :  254 - 0xfe
    "00111000", -- 2964 - 0xb94  :   56 - 0x38
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "11111111", -- 2968 - 0xb98  :  255 - 0xff -- Background 0x73
    "11111111", -- 2969 - 0xb99  :  255 - 0xff
    "11111101", -- 2970 - 0xb9a  :  253 - 0xfd
    "11111111", -- 2971 - 0xb9b  :  255 - 0xff
    "10111111", -- 2972 - 0xb9c  :  191 - 0xbf
    "11111111", -- 2973 - 0xb9d  :  255 - 0xff
    "11111111", -- 2974 - 0xb9e  :  255 - 0xff
    "11110111", -- 2975 - 0xb9f  :  247 - 0xf7
    "01000110", -- 2976 - 0xba0  :   70 - 0x46 -- Background 0x74
    "01101011", -- 2977 - 0xba1  :  107 - 0x6b
    "01110001", -- 2978 - 0xba2  :  113 - 0x71
    "00111010", -- 2979 - 0xba3  :   58 - 0x3a
    "01101101", -- 2980 - 0xba4  :  109 - 0x6d
    "00111000", -- 2981 - 0xba5  :   56 - 0x38
    "00011101", -- 2982 - 0xba6  :   29 - 0x1d
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "01000110", -- 2984 - 0xba8  :   70 - 0x46 -- Background 0x75
    "11101011", -- 2985 - 0xba9  :  235 - 0xeb
    "01110001", -- 2986 - 0xbaa  :  113 - 0x71
    "00111010", -- 2987 - 0xbab  :   58 - 0x3a
    "01101101", -- 2988 - 0xbac  :  109 - 0x6d
    "10111000", -- 2989 - 0xbad  :  184 - 0xb8
    "00011101", -- 2990 - 0xbae  :   29 - 0x1d
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "01000110", -- 2992 - 0xbb0  :   70 - 0x46 -- Background 0x76
    "11101010", -- 2993 - 0xbb1  :  234 - 0xea
    "01110000", -- 2994 - 0xbb2  :  112 - 0x70
    "00111010", -- 2995 - 0xbb3  :   58 - 0x3a
    "01101100", -- 2996 - 0xbb4  :  108 - 0x6c
    "10111000", -- 2997 - 0xbb5  :  184 - 0xb8
    "00011100", -- 2998 - 0xbb6  :   28 - 0x1c
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "10000001", -- 3000 - 0xbb8  :  129 - 0x81 -- Background 0x77
    "11111111", -- 3001 - 0xbb9  :  255 - 0xff
    "11111101", -- 3002 - 0xbba  :  253 - 0xfd
    "11111111", -- 3003 - 0xbbb  :  255 - 0xff
    "10111111", -- 3004 - 0xbbc  :  191 - 0xbf
    "11111111", -- 3005 - 0xbbd  :  255 - 0xff
    "11111111", -- 3006 - 0xbbe  :  255 - 0xff
    "11110111", -- 3007 - 0xbbf  :  247 - 0xf7
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- Background 0x79
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Background 0x7c
    "00100010", -- 3041 - 0xbe1  :   34 - 0x22
    "01110111", -- 3042 - 0xbe2  :  119 - 0x77
    "11111111", -- 3043 - 0xbe3  :  255 - 0xff
    "11111011", -- 3044 - 0xbe4  :  251 - 0xfb
    "11110101", -- 3045 - 0xbe5  :  245 - 0xf5
    "11101111", -- 3046 - 0xbe6  :  239 - 0xef
    "11111111", -- 3047 - 0xbe7  :  255 - 0xff
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- Background 0x7d
    "01110011", -- 3049 - 0xbe9  :  115 - 0x73
    "11111111", -- 3050 - 0xbea  :  255 - 0xff
    "11111111", -- 3051 - 0xbeb  :  255 - 0xff
    "11111011", -- 3052 - 0xbec  :  251 - 0xfb
    "11111101", -- 3053 - 0xbed  :  253 - 0xfd
    "11101111", -- 3054 - 0xbee  :  239 - 0xef
    "11111111", -- 3055 - 0xbef  :  255 - 0xff
    "11011111", -- 3056 - 0xbf0  :  223 - 0xdf -- Background 0x7e
    "10101111", -- 3057 - 0xbf1  :  175 - 0xaf
    "01111111", -- 3058 - 0xbf2  :  127 - 0x7f
    "11111111", -- 3059 - 0xbf3  :  255 - 0xff
    "11111011", -- 3060 - 0xbf4  :  251 - 0xfb
    "11110101", -- 3061 - 0xbf5  :  245 - 0xf5
    "11101111", -- 3062 - 0xbf6  :  239 - 0xef
    "11111111", -- 3063 - 0xbf7  :  255 - 0xff
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- Background 0x7f
    "10101111", -- 3065 - 0xbf9  :  175 - 0xaf
    "01111111", -- 3066 - 0xbfa  :  127 - 0x7f
    "11111111", -- 3067 - 0xbfb  :  255 - 0xff
    "11111011", -- 3068 - 0xbfc  :  251 - 0xfb
    "11110101", -- 3069 - 0xbfd  :  245 - 0xf5
    "11101111", -- 3070 - 0xbfe  :  239 - 0xef
    "11111111", -- 3071 - 0xbff  :  255 - 0xff
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0x80
    "01111111", -- 3073 - 0xc01  :  127 - 0x7f
    "00110000", -- 3074 - 0xc02  :   48 - 0x30
    "00110000", -- 3075 - 0xc03  :   48 - 0x30
    "00110000", -- 3076 - 0xc04  :   48 - 0x30
    "01111111", -- 3077 - 0xc05  :  127 - 0x7f
    "00110000", -- 3078 - 0xc06  :   48 - 0x30
    "00110000", -- 3079 - 0xc07  :   48 - 0x30
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- Background 0x81
    "01111111", -- 3081 - 0xc09  :  127 - 0x7f
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "01111111", -- 3083 - 0xc0b  :  127 - 0x7f
    "01111111", -- 3084 - 0xc0c  :  127 - 0x7f
    "00100000", -- 3085 - 0xc0d  :   32 - 0x20
    "01000000", -- 3086 - 0xc0e  :   64 - 0x40
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Background 0x82
    "11111110", -- 3089 - 0xc11  :  254 - 0xfe
    "00001100", -- 3090 - 0xc12  :   12 - 0xc
    "00001100", -- 3091 - 0xc13  :   12 - 0xc
    "00001100", -- 3092 - 0xc14  :   12 - 0xc
    "11111110", -- 3093 - 0xc15  :  254 - 0xfe
    "00001100", -- 3094 - 0xc16  :   12 - 0xc
    "00001100", -- 3095 - 0xc17  :   12 - 0xc
    "00000000", -- 3096 - 0xc18  :    0 - 0x0 -- Background 0x83
    "11111111", -- 3097 - 0xc19  :  255 - 0xff
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "11111111", -- 3099 - 0xc1b  :  255 - 0xff
    "11111111", -- 3100 - 0xc1c  :  255 - 0xff
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0x84
    "11111111", -- 3105 - 0xc21  :  255 - 0xff
    "11111111", -- 3106 - 0xc22  :  255 - 0xff
    "11111111", -- 3107 - 0xc23  :  255 - 0xff
    "11111111", -- 3108 - 0xc24  :  255 - 0xff
    "11101111", -- 3109 - 0xc25  :  239 - 0xef
    "10111011", -- 3110 - 0xc26  :  187 - 0xbb
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- Background 0x85
    "11111110", -- 3113 - 0xc29  :  254 - 0xfe
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "11111110", -- 3115 - 0xc2b  :  254 - 0xfe
    "11111110", -- 3116 - 0xc2c  :  254 - 0xfe
    "00001100", -- 3117 - 0xc2d  :   12 - 0xc
    "00000010", -- 3118 - 0xc2e  :    2 - 0x2
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0x86
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "00000000", -- 3126 - 0xc36  :    0 - 0x0
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- Background 0x87
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0x88
    "00000111", -- 3137 - 0xc41  :    7 - 0x7
    "00011111", -- 3138 - 0xc42  :   31 - 0x1f
    "00111100", -- 3139 - 0xc43  :   60 - 0x3c
    "00110001", -- 3140 - 0xc44  :   49 - 0x31
    "01110100", -- 3141 - 0xc45  :  116 - 0x74
    "01100101", -- 3142 - 0xc46  :  101 - 0x65
    "01101010", -- 3143 - 0xc47  :  106 - 0x6a
    "01100100", -- 3144 - 0xc48  :  100 - 0x64 -- Background 0x89
    "01101101", -- 3145 - 0xc49  :  109 - 0x6d
    "01110010", -- 3146 - 0xc4a  :  114 - 0x72
    "00110000", -- 3147 - 0xc4b  :   48 - 0x30
    "00111100", -- 3148 - 0xc4c  :   60 - 0x3c
    "00011111", -- 3149 - 0xc4d  :   31 - 0x1f
    "00000111", -- 3150 - 0xc4e  :    7 - 0x7
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0x8a
    "11100000", -- 3153 - 0xc51  :  224 - 0xe0
    "11111000", -- 3154 - 0xc52  :  248 - 0xf8
    "00111100", -- 3155 - 0xc53  :   60 - 0x3c
    "01001100", -- 3156 - 0xc54  :   76 - 0x4c
    "01101110", -- 3157 - 0xc55  :  110 - 0x6e
    "00100110", -- 3158 - 0xc56  :   38 - 0x26
    "01000110", -- 3159 - 0xc57  :   70 - 0x46
    "10010110", -- 3160 - 0xc58  :  150 - 0x96 -- Background 0x8b
    "01100110", -- 3161 - 0xc59  :  102 - 0x66
    "10101110", -- 3162 - 0xc5a  :  174 - 0xae
    "01001100", -- 3163 - 0xc5b  :   76 - 0x4c
    "00111100", -- 3164 - 0xc5c  :   60 - 0x3c
    "11111000", -- 3165 - 0xc5d  :  248 - 0xf8
    "11100000", -- 3166 - 0xc5e  :  224 - 0xe0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Background 0x8c
    "00000111", -- 3169 - 0xc61  :    7 - 0x7
    "00011111", -- 3170 - 0xc62  :   31 - 0x1f
    "00111111", -- 3171 - 0xc63  :   63 - 0x3f
    "00111111", -- 3172 - 0xc64  :   63 - 0x3f
    "01111111", -- 3173 - 0xc65  :  127 - 0x7f
    "01111111", -- 3174 - 0xc66  :  127 - 0x7f
    "01111111", -- 3175 - 0xc67  :  127 - 0x7f
    "01111111", -- 3176 - 0xc68  :  127 - 0x7f -- Background 0x8d
    "01111111", -- 3177 - 0xc69  :  127 - 0x7f
    "01111111", -- 3178 - 0xc6a  :  127 - 0x7f
    "00111111", -- 3179 - 0xc6b  :   63 - 0x3f
    "00111111", -- 3180 - 0xc6c  :   63 - 0x3f
    "00011111", -- 3181 - 0xc6d  :   31 - 0x1f
    "00000111", -- 3182 - 0xc6e  :    7 - 0x7
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000000", -- 3184 - 0xc70  :    0 - 0x0 -- Background 0x8e
    "11100000", -- 3185 - 0xc71  :  224 - 0xe0
    "11111000", -- 3186 - 0xc72  :  248 - 0xf8
    "11111100", -- 3187 - 0xc73  :  252 - 0xfc
    "11111100", -- 3188 - 0xc74  :  252 - 0xfc
    "11111110", -- 3189 - 0xc75  :  254 - 0xfe
    "11111110", -- 3190 - 0xc76  :  254 - 0xfe
    "11111110", -- 3191 - 0xc77  :  254 - 0xfe
    "11111110", -- 3192 - 0xc78  :  254 - 0xfe -- Background 0x8f
    "11111110", -- 3193 - 0xc79  :  254 - 0xfe
    "11111110", -- 3194 - 0xc7a  :  254 - 0xfe
    "11111100", -- 3195 - 0xc7b  :  252 - 0xfc
    "11111100", -- 3196 - 0xc7c  :  252 - 0xfc
    "11111000", -- 3197 - 0xc7d  :  248 - 0xf8
    "11100000", -- 3198 - 0xc7e  :  224 - 0xe0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00010000", -- 3204 - 0xc84  :   16 - 0x10
    "00011100", -- 3205 - 0xc85  :   28 - 0x1c
    "00001110", -- 3206 - 0xc86  :   14 - 0xe
    "00000111", -- 3207 - 0xc87  :    7 - 0x7
    "00000011", -- 3208 - 0xc88  :    3 - 0x3 -- Background 0x91
    "00000001", -- 3209 - 0xc89  :    1 - 0x1
    "00110000", -- 3210 - 0xc8a  :   48 - 0x30
    "00001111", -- 3211 - 0xc8b  :   15 - 0xf
    "00000011", -- 3212 - 0xc8c  :    3 - 0x3
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "01111111", -- 3214 - 0xc8e  :  127 - 0x7f
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00000000", -- 3216 - 0xc90  :    0 - 0x0 -- Background 0x92
    "01000010", -- 3217 - 0xc91  :   66 - 0x42
    "01000010", -- 3218 - 0xc92  :   66 - 0x42
    "01100110", -- 3219 - 0xc93  :  102 - 0x66
    "01100110", -- 3220 - 0xc94  :  102 - 0x66
    "01100110", -- 3221 - 0xc95  :  102 - 0x66
    "11111110", -- 3222 - 0xc96  :  254 - 0xfe
    "11111111", -- 3223 - 0xc97  :  255 - 0xff
    "01111110", -- 3224 - 0xc98  :  126 - 0x7e -- Background 0x93
    "01111110", -- 3225 - 0xc99  :  126 - 0x7e
    "01111110", -- 3226 - 0xc9a  :  126 - 0x7e
    "01111110", -- 3227 - 0xc9b  :  126 - 0x7e
    "01111110", -- 3228 - 0xc9c  :  126 - 0x7e
    "01111110", -- 3229 - 0xc9d  :  126 - 0x7e
    "01111110", -- 3230 - 0xc9e  :  126 - 0x7e
    "01111110", -- 3231 - 0xc9f  :  126 - 0x7e
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00000000", -- 3235 - 0xca3  :    0 - 0x0
    "00001000", -- 3236 - 0xca4  :    8 - 0x8
    "00111000", -- 3237 - 0xca5  :   56 - 0x38
    "01110000", -- 3238 - 0xca6  :  112 - 0x70
    "11100000", -- 3239 - 0xca7  :  224 - 0xe0
    "11000000", -- 3240 - 0xca8  :  192 - 0xc0 -- Background 0x95
    "10000000", -- 3241 - 0xca9  :  128 - 0x80
    "00001100", -- 3242 - 0xcaa  :   12 - 0xc
    "11110000", -- 3243 - 0xcab  :  240 - 0xf0
    "11000000", -- 3244 - 0xcac  :  192 - 0xc0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "11111110", -- 3246 - 0xcae  :  254 - 0xfe
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Background 0x96
    "00111111", -- 3249 - 0xcb1  :   63 - 0x3f
    "01111111", -- 3250 - 0xcb2  :  127 - 0x7f
    "01111111", -- 3251 - 0xcb3  :  127 - 0x7f
    "01111111", -- 3252 - 0xcb4  :  127 - 0x7f
    "01111111", -- 3253 - 0xcb5  :  127 - 0x7f
    "01111111", -- 3254 - 0xcb6  :  127 - 0x7f
    "01111111", -- 3255 - 0xcb7  :  127 - 0x7f
    "01111111", -- 3256 - 0xcb8  :  127 - 0x7f -- Background 0x97
    "01111111", -- 3257 - 0xcb9  :  127 - 0x7f
    "00111111", -- 3258 - 0xcba  :   63 - 0x3f
    "01111111", -- 3259 - 0xcbb  :  127 - 0x7f
    "01111111", -- 3260 - 0xcbc  :  127 - 0x7f
    "01111111", -- 3261 - 0xcbd  :  127 - 0x7f
    "01111111", -- 3262 - 0xcbe  :  127 - 0x7f
    "01111111", -- 3263 - 0xcbf  :  127 - 0x7f
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Background 0x98
    "11011111", -- 3265 - 0xcc1  :  223 - 0xdf
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111111", -- 3267 - 0xcc3  :  255 - 0xff
    "11111111", -- 3268 - 0xcc4  :  255 - 0xff
    "11111111", -- 3269 - 0xcc5  :  255 - 0xff
    "11111111", -- 3270 - 0xcc6  :  255 - 0xff
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "11111111", -- 3272 - 0xcc8  :  255 - 0xff -- Background 0x99
    "11111111", -- 3273 - 0xcc9  :  255 - 0xff
    "10111111", -- 3274 - 0xcca  :  191 - 0xbf
    "11111111", -- 3275 - 0xccb  :  255 - 0xff
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "11111111", -- 3277 - 0xccd  :  255 - 0xff
    "11111111", -- 3278 - 0xcce  :  255 - 0xff
    "11111111", -- 3279 - 0xccf  :  255 - 0xff
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0x9a
    "10111100", -- 3281 - 0xcd1  :  188 - 0xbc
    "11111110", -- 3282 - 0xcd2  :  254 - 0xfe
    "11111110", -- 3283 - 0xcd3  :  254 - 0xfe
    "11111110", -- 3284 - 0xcd4  :  254 - 0xfe
    "11111110", -- 3285 - 0xcd5  :  254 - 0xfe
    "11111110", -- 3286 - 0xcd6  :  254 - 0xfe
    "11111110", -- 3287 - 0xcd7  :  254 - 0xfe
    "11111110", -- 3288 - 0xcd8  :  254 - 0xfe -- Background 0x9b
    "11111110", -- 3289 - 0xcd9  :  254 - 0xfe
    "10111110", -- 3290 - 0xcda  :  190 - 0xbe
    "11111110", -- 3291 - 0xcdb  :  254 - 0xfe
    "11111110", -- 3292 - 0xcdc  :  254 - 0xfe
    "11111110", -- 3293 - 0xcdd  :  254 - 0xfe
    "11111110", -- 3294 - 0xcde  :  254 - 0xfe
    "11111110", -- 3295 - 0xcdf  :  254 - 0xfe
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0x9c
    "00111111", -- 3297 - 0xce1  :   63 - 0x3f
    "01011111", -- 3298 - 0xce2  :   95 - 0x5f
    "01101111", -- 3299 - 0xce3  :  111 - 0x6f
    "01110111", -- 3300 - 0xce4  :  119 - 0x77
    "01111011", -- 3301 - 0xce5  :  123 - 0x7b
    "00010101", -- 3302 - 0xce6  :   21 - 0x15
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- Background 0x9d
    "10111110", -- 3305 - 0xce9  :  190 - 0xbe
    "11011110", -- 3306 - 0xcea  :  222 - 0xde
    "11101110", -- 3307 - 0xceb  :  238 - 0xee
    "11110110", -- 3308 - 0xcec  :  246 - 0xf6
    "11111010", -- 3309 - 0xced  :  250 - 0xfa
    "01010100", -- 3310 - 0xcee  :   84 - 0x54
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Background 0x9e
    "10111111", -- 3313 - 0xcf1  :  191 - 0xbf
    "11011111", -- 3314 - 0xcf2  :  223 - 0xdf
    "11101111", -- 3315 - 0xcf3  :  239 - 0xef
    "11110111", -- 3316 - 0xcf4  :  247 - 0xf7
    "11111011", -- 3317 - 0xcf5  :  251 - 0xfb
    "01010101", -- 3318 - 0xcf6  :   85 - 0x55
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Background 0xa0
    "01111111", -- 3329 - 0xd01  :  127 - 0x7f
    "00000000", -- 3330 - 0xd02  :    0 - 0x0
    "00000001", -- 3331 - 0xd03  :    1 - 0x1
    "00000001", -- 3332 - 0xd04  :    1 - 0x1
    "00000001", -- 3333 - 0xd05  :    1 - 0x1
    "00000001", -- 3334 - 0xd06  :    1 - 0x1
    "00000001", -- 3335 - 0xd07  :    1 - 0x1
    "00000001", -- 3336 - 0xd08  :    1 - 0x1 -- Background 0xa1
    "00000001", -- 3337 - 0xd09  :    1 - 0x1
    "00000001", -- 3338 - 0xd0a  :    1 - 0x1
    "00000001", -- 3339 - 0xd0b  :    1 - 0x1
    "00000001", -- 3340 - 0xd0c  :    1 - 0x1
    "00000001", -- 3341 - 0xd0d  :    1 - 0x1
    "00000001", -- 3342 - 0xd0e  :    1 - 0x1
    "00000001", -- 3343 - 0xd0f  :    1 - 0x1
    "00000000", -- 3344 - 0xd10  :    0 - 0x0 -- Background 0xa2
    "11111110", -- 3345 - 0xd11  :  254 - 0xfe
    "00000000", -- 3346 - 0xd12  :    0 - 0x0
    "10000000", -- 3347 - 0xd13  :  128 - 0x80
    "10000000", -- 3348 - 0xd14  :  128 - 0x80
    "10000000", -- 3349 - 0xd15  :  128 - 0x80
    "10000000", -- 3350 - 0xd16  :  128 - 0x80
    "10000000", -- 3351 - 0xd17  :  128 - 0x80
    "10000000", -- 3352 - 0xd18  :  128 - 0x80 -- Background 0xa3
    "10000000", -- 3353 - 0xd19  :  128 - 0x80
    "10000000", -- 3354 - 0xd1a  :  128 - 0x80
    "10000000", -- 3355 - 0xd1b  :  128 - 0x80
    "10000000", -- 3356 - 0xd1c  :  128 - 0x80
    "10000000", -- 3357 - 0xd1d  :  128 - 0x80
    "10000000", -- 3358 - 0xd1e  :  128 - 0x80
    "10000000", -- 3359 - 0xd1f  :  128 - 0x80
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xa4
    "00110000", -- 3361 - 0xd21  :   48 - 0x30
    "00111000", -- 3362 - 0xd22  :   56 - 0x38
    "01111000", -- 3363 - 0xd23  :  120 - 0x78
    "01111100", -- 3364 - 0xd24  :  124 - 0x7c
    "01111101", -- 3365 - 0xd25  :  125 - 0x7d
    "00011101", -- 3366 - 0xd26  :   29 - 0x1d
    "00001101", -- 3367 - 0xd27  :   13 - 0xd
    "00001101", -- 3368 - 0xd28  :   13 - 0xd -- Background 0xa5
    "00011101", -- 3369 - 0xd29  :   29 - 0x1d
    "00111101", -- 3370 - 0xd2a  :   61 - 0x3d
    "00111111", -- 3371 - 0xd2b  :   63 - 0x3f
    "00111111", -- 3372 - 0xd2c  :   63 - 0x3f
    "00011111", -- 3373 - 0xd2d  :   31 - 0x1f
    "00000001", -- 3374 - 0xd2e  :    1 - 0x1
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00000000", -- 3376 - 0xd30  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "11100000", -- 3378 - 0xd32  :  224 - 0xe0
    "11111000", -- 3379 - 0xd33  :  248 - 0xf8
    "11111000", -- 3380 - 0xd34  :  248 - 0xf8
    "11110000", -- 3381 - 0xd35  :  240 - 0xf0
    "11000000", -- 3382 - 0xd36  :  192 - 0xc0
    "11000000", -- 3383 - 0xd37  :  192 - 0xc0
    "11000000", -- 3384 - 0xd38  :  192 - 0xc0 -- Background 0xa7
    "11110000", -- 3385 - 0xd39  :  240 - 0xf0
    "11110000", -- 3386 - 0xd3a  :  240 - 0xf0
    "11000000", -- 3387 - 0xd3b  :  192 - 0xc0
    "11000000", -- 3388 - 0xd3c  :  192 - 0xc0
    "11000000", -- 3389 - 0xd3d  :  192 - 0xc0
    "11000000", -- 3390 - 0xd3e  :  192 - 0xc0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xa8
    "01100000", -- 3393 - 0xd41  :   96 - 0x60
    "01100000", -- 3394 - 0xd42  :   96 - 0x60
    "01100000", -- 3395 - 0xd43  :   96 - 0x60
    "01100000", -- 3396 - 0xd44  :   96 - 0x60
    "01100000", -- 3397 - 0xd45  :   96 - 0x60
    "01100000", -- 3398 - 0xd46  :   96 - 0x60
    "01100000", -- 3399 - 0xd47  :   96 - 0x60
    "01100000", -- 3400 - 0xd48  :   96 - 0x60 -- Background 0xa9
    "01100000", -- 3401 - 0xd49  :   96 - 0x60
    "01100000", -- 3402 - 0xd4a  :   96 - 0x60
    "01100000", -- 3403 - 0xd4b  :   96 - 0x60
    "01100000", -- 3404 - 0xd4c  :   96 - 0x60
    "01100000", -- 3405 - 0xd4d  :   96 - 0x60
    "01100000", -- 3406 - 0xd4e  :   96 - 0x60
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Background 0xaa
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- Background 0xab
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000000", -- 3419 - 0xd5b  :    0 - 0x0
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00000000", -- 3422 - 0xd5e  :    0 - 0x0
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xac
    "00000110", -- 3425 - 0xd61  :    6 - 0x6
    "00000110", -- 3426 - 0xd62  :    6 - 0x6
    "00000110", -- 3427 - 0xd63  :    6 - 0x6
    "00000110", -- 3428 - 0xd64  :    6 - 0x6
    "00000110", -- 3429 - 0xd65  :    6 - 0x6
    "00000110", -- 3430 - 0xd66  :    6 - 0x6
    "00000110", -- 3431 - 0xd67  :    6 - 0x6
    "00000110", -- 3432 - 0xd68  :    6 - 0x6 -- Background 0xad
    "00000110", -- 3433 - 0xd69  :    6 - 0x6
    "00000110", -- 3434 - 0xd6a  :    6 - 0x6
    "00000110", -- 3435 - 0xd6b  :    6 - 0x6
    "00000110", -- 3436 - 0xd6c  :    6 - 0x6
    "00000110", -- 3437 - 0xd6d  :    6 - 0x6
    "00000110", -- 3438 - 0xd6e  :    6 - 0x6
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "00000000", -- 3440 - 0xd70  :    0 - 0x0 -- Background 0xae
    "00000001", -- 3441 - 0xd71  :    1 - 0x1
    "00000011", -- 3442 - 0xd72  :    3 - 0x3
    "00000010", -- 3443 - 0xd73  :    2 - 0x2
    "00000010", -- 3444 - 0xd74  :    2 - 0x2
    "00000000", -- 3445 - 0xd75  :    0 - 0x0
    "00000011", -- 3446 - 0xd76  :    3 - 0x3
    "00000010", -- 3447 - 0xd77  :    2 - 0x2
    "00000001", -- 3448 - 0xd78  :    1 - 0x1 -- Background 0xaf
    "00000011", -- 3449 - 0xd79  :    3 - 0x3
    "00000101", -- 3450 - 0xd7a  :    5 - 0x5
    "00000100", -- 3451 - 0xd7b  :    4 - 0x4
    "00000101", -- 3452 - 0xd7c  :    5 - 0x5
    "00001101", -- 3453 - 0xd7d  :   13 - 0xd
    "00001100", -- 3454 - 0xd7e  :   12 - 0xc
    "00000001", -- 3455 - 0xd7f  :    1 - 0x1
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xb0
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "01000000", -- 3458 - 0xd82  :   64 - 0x40
    "11110000", -- 3459 - 0xd83  :  240 - 0xf0
    "11101000", -- 3460 - 0xd84  :  232 - 0xe8
    "10010000", -- 3461 - 0xd85  :  144 - 0x90
    "01010000", -- 3462 - 0xd86  :   80 - 0x50
    "11010000", -- 3463 - 0xd87  :  208 - 0xd0
    "11111000", -- 3464 - 0xd88  :  248 - 0xf8 -- Background 0xb1
    "11000000", -- 3465 - 0xd89  :  192 - 0xc0
    "11100000", -- 3466 - 0xd8a  :  224 - 0xe0
    "01000000", -- 3467 - 0xd8b  :   64 - 0x40
    "10000000", -- 3468 - 0xd8c  :  128 - 0x80
    "11000000", -- 3469 - 0xd8d  :  192 - 0xc0
    "11100000", -- 3470 - 0xd8e  :  224 - 0xe0
    "01110000", -- 3471 - 0xd8f  :  112 - 0x70
    "00000001", -- 3472 - 0xd90  :    1 - 0x1 -- Background 0xb2
    "00001101", -- 3473 - 0xd91  :   13 - 0xd
    "00001101", -- 3474 - 0xd92  :   13 - 0xd
    "00000011", -- 3475 - 0xd93  :    3 - 0x3
    "00000011", -- 3476 - 0xd94  :    3 - 0x3
    "00000111", -- 3477 - 0xd95  :    7 - 0x7
    "00000111", -- 3478 - 0xd96  :    7 - 0x7
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "00111111", -- 3480 - 0xd98  :   63 - 0x3f -- Background 0xb3
    "00111111", -- 3481 - 0xd99  :   63 - 0x3f
    "00111111", -- 3482 - 0xd9a  :   63 - 0x3f
    "00111111", -- 3483 - 0xd9b  :   63 - 0x3f
    "00111111", -- 3484 - 0xd9c  :   63 - 0x3f
    "00111111", -- 3485 - 0xd9d  :   63 - 0x3f
    "00110101", -- 3486 - 0xd9e  :   53 - 0x35
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "10110000", -- 3488 - 0xda0  :  176 - 0xb0 -- Background 0xb4
    "11000000", -- 3489 - 0xda1  :  192 - 0xc0
    "11100000", -- 3490 - 0xda2  :  224 - 0xe0
    "11100000", -- 3491 - 0xda3  :  224 - 0xe0
    "11110000", -- 3492 - 0xda4  :  240 - 0xf0
    "11110000", -- 3493 - 0xda5  :  240 - 0xf0
    "11110000", -- 3494 - 0xda6  :  240 - 0xf0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "11111100", -- 3496 - 0xda8  :  252 - 0xfc -- Background 0xb5
    "11111000", -- 3497 - 0xda9  :  248 - 0xf8
    "11111100", -- 3498 - 0xdaa  :  252 - 0xfc
    "11111000", -- 3499 - 0xdab  :  248 - 0xf8
    "11111100", -- 3500 - 0xdac  :  252 - 0xfc
    "11111000", -- 3501 - 0xdad  :  248 - 0xf8
    "01010100", -- 3502 - 0xdae  :   84 - 0x54
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Background 0xb6
    "01111111", -- 3505 - 0xdb1  :  127 - 0x7f
    "01111111", -- 3506 - 0xdb2  :  127 - 0x7f
    "01111111", -- 3507 - 0xdb3  :  127 - 0x7f
    "01111111", -- 3508 - 0xdb4  :  127 - 0x7f
    "01111111", -- 3509 - 0xdb5  :  127 - 0x7f
    "01101010", -- 3510 - 0xdb6  :  106 - 0x6a
    "00000000", -- 3511 - 0xdb7  :    0 - 0x0
    "00000000", -- 3512 - 0xdb8  :    0 - 0x0 -- Background 0xb7
    "01111011", -- 3513 - 0xdb9  :  123 - 0x7b
    "01110011", -- 3514 - 0xdba  :  115 - 0x73
    "01111011", -- 3515 - 0xdbb  :  123 - 0x7b
    "01110011", -- 3516 - 0xdbc  :  115 - 0x73
    "01111011", -- 3517 - 0xdbd  :  123 - 0x7b
    "01010011", -- 3518 - 0xdbe  :   83 - 0x53
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xb8
    "11011110", -- 3521 - 0xdc1  :  222 - 0xde
    "10011110", -- 3522 - 0xdc2  :  158 - 0x9e
    "11011100", -- 3523 - 0xdc3  :  220 - 0xdc
    "10011110", -- 3524 - 0xdc4  :  158 - 0x9e
    "11011100", -- 3525 - 0xdc5  :  220 - 0xdc
    "10011010", -- 3526 - 0xdc6  :  154 - 0x9a
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0 -- Background 0xb9
    "11111110", -- 3529 - 0xdc9  :  254 - 0xfe
    "11111100", -- 3530 - 0xdca  :  252 - 0xfc
    "11111110", -- 3531 - 0xdcb  :  254 - 0xfe
    "11111100", -- 3532 - 0xdcc  :  252 - 0xfc
    "11111110", -- 3533 - 0xdcd  :  254 - 0xfe
    "01010100", -- 3534 - 0xdce  :   84 - 0x54
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Background 0xba
    "01111111", -- 3537 - 0xdd1  :  127 - 0x7f
    "01111111", -- 3538 - 0xdd2  :  127 - 0x7f
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "01111111", -- 3540 - 0xdd4  :  127 - 0x7f
    "01111111", -- 3541 - 0xdd5  :  127 - 0x7f
    "01101010", -- 3542 - 0xdd6  :  106 - 0x6a
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0 -- Background 0xbb
    "00000000", -- 3545 - 0xdd9  :    0 - 0x0
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Background 0xbc
    "11111110", -- 3553 - 0xde1  :  254 - 0xfe
    "11111110", -- 3554 - 0xde2  :  254 - 0xfe
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "10011110", -- 3556 - 0xde4  :  158 - 0x9e
    "11011100", -- 3557 - 0xde5  :  220 - 0xdc
    "10011010", -- 3558 - 0xde6  :  154 - 0x9a
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "00000000", -- 3560 - 0xde8  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 3569 - 0xdf1  :    0 - 0x0
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "00000000", -- 3573 - 0xdf5  :    0 - 0x0
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00000000", -- 3592 - 0xe08  :    0 - 0x0 -- Background 0xc1
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00000000", -- 3594 - 0xe0a  :    0 - 0x0
    "00000000", -- 3595 - 0xe0b  :    0 - 0x0
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00000000", -- 3608 - 0xe18  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00000000", -- 3611 - 0xe1b  :    0 - 0x0
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "00000000", -- 3624 - 0xe28  :    0 - 0x0 -- Background 0xc5
    "00000000", -- 3625 - 0xe29  :    0 - 0x0
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "00000001", -- 3627 - 0xe2b  :    1 - 0x1
    "00000111", -- 3628 - 0xe2c  :    7 - 0x7
    "00001111", -- 3629 - 0xe2d  :   15 - 0xf
    "00001111", -- 3630 - 0xe2e  :   15 - 0xf
    "00011111", -- 3631 - 0xe2f  :   31 - 0x1f
    "00000000", -- 3632 - 0xe30  :    0 - 0x0 -- Background 0xc6
    "00011111", -- 3633 - 0xe31  :   31 - 0x1f
    "01111111", -- 3634 - 0xe32  :  127 - 0x7f
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "11111111", -- 3636 - 0xe34  :  255 - 0xff
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "00011111", -- 3640 - 0xe38  :   31 - 0x1f -- Background 0xc7
    "00111111", -- 3641 - 0xe39  :   63 - 0x3f
    "00111111", -- 3642 - 0xe3a  :   63 - 0x3f
    "01111111", -- 3643 - 0xe3b  :  127 - 0x7f
    "01111111", -- 3644 - 0xe3c  :  127 - 0x7f
    "01111111", -- 3645 - 0xe3d  :  127 - 0x7f
    "01111111", -- 3646 - 0xe3e  :  127 - 0x7f
    "01111111", -- 3647 - 0xe3f  :  127 - 0x7f
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xc8
    "11111111", -- 3649 - 0xe41  :  255 - 0xff
    "11111111", -- 3650 - 0xe42  :  255 - 0xff
    "11111111", -- 3651 - 0xe43  :  255 - 0xff
    "11111111", -- 3652 - 0xe44  :  255 - 0xff
    "11111111", -- 3653 - 0xe45  :  255 - 0xff
    "11111111", -- 3654 - 0xe46  :  255 - 0xff
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11101000", -- 3656 - 0xe48  :  232 - 0xe8 -- Background 0xc9
    "11010100", -- 3657 - 0xe49  :  212 - 0xd4
    "11101000", -- 3658 - 0xe4a  :  232 - 0xe8
    "11010100", -- 3659 - 0xe4b  :  212 - 0xd4
    "11101010", -- 3660 - 0xe4c  :  234 - 0xea
    "11010100", -- 3661 - 0xe4d  :  212 - 0xd4
    "11101010", -- 3662 - 0xe4e  :  234 - 0xea
    "11010100", -- 3663 - 0xe4f  :  212 - 0xd4
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Background 0xca
    "00000000", -- 3665 - 0xe51  :    0 - 0x0
    "00000000", -- 3666 - 0xe52  :    0 - 0x0
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00000000", -- 3669 - 0xe55  :    0 - 0x0
    "00000000", -- 3670 - 0xe56  :    0 - 0x0
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00000000", -- 3677 - 0xe5d  :    0 - 0x0
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000101", -- 3684 - 0xe64  :    5 - 0x5
    "00000010", -- 3685 - 0xe65  :    2 - 0x2
    "00000001", -- 3686 - 0xe66  :    1 - 0x1
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "10000000", -- 3691 - 0xe6b  :  128 - 0x80
    "01010000", -- 3692 - 0xe6c  :   80 - 0x50
    "10100000", -- 3693 - 0xe6d  :  160 - 0xa0
    "01000000", -- 3694 - 0xe6e  :   64 - 0x40
    "10000000", -- 3695 - 0xe6f  :  128 - 0x80
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00110000", -- 3700 - 0xe74  :   48 - 0x30
    "01111111", -- 3701 - 0xe75  :  127 - 0x7f
    "00110000", -- 3702 - 0xe76  :   48 - 0x30
    "00110000", -- 3703 - 0xe77  :   48 - 0x30
    "00000000", -- 3704 - 0xe78  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00001100", -- 3708 - 0xe7c  :   12 - 0xc
    "11111110", -- 3709 - 0xe7d  :  254 - 0xfe
    "00001100", -- 3710 - 0xe7e  :   12 - 0xc
    "00001100", -- 3711 - 0xe7f  :   12 - 0xc
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000111", -- 3728 - 0xe90  :    7 - 0x7 -- Background 0xd2
    "00000111", -- 3729 - 0xe91  :    7 - 0x7
    "00000111", -- 3730 - 0xe92  :    7 - 0x7
    "00000111", -- 3731 - 0xe93  :    7 - 0x7
    "00000111", -- 3732 - 0xe94  :    7 - 0x7
    "00000111", -- 3733 - 0xe95  :    7 - 0x7
    "00000111", -- 3734 - 0xe96  :    7 - 0x7
    "00000111", -- 3735 - 0xe97  :    7 - 0x7
    "11100000", -- 3736 - 0xe98  :  224 - 0xe0 -- Background 0xd3
    "11100000", -- 3737 - 0xe99  :  224 - 0xe0
    "11000000", -- 3738 - 0xe9a  :  192 - 0xc0
    "11100000", -- 3739 - 0xe9b  :  224 - 0xe0
    "10100000", -- 3740 - 0xe9c  :  160 - 0xa0
    "11100000", -- 3741 - 0xe9d  :  224 - 0xe0
    "11000000", -- 3742 - 0xe9e  :  192 - 0xc0
    "11100000", -- 3743 - 0xe9f  :  224 - 0xe0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0 -- Background 0xd5
    "11111000", -- 3753 - 0xea9  :  248 - 0xf8
    "11111110", -- 3754 - 0xeaa  :  254 - 0xfe
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "10000000", -- 3763 - 0xeb3  :  128 - 0x80
    "10100000", -- 3764 - 0xeb4  :  160 - 0xa0
    "01010000", -- 3765 - 0xeb5  :   80 - 0x50
    "10100000", -- 3766 - 0xeb6  :  160 - 0xa0
    "11010000", -- 3767 - 0xeb7  :  208 - 0xd0
    "01111111", -- 3768 - 0xeb8  :  127 - 0x7f -- Background 0xd7
    "01111111", -- 3769 - 0xeb9  :  127 - 0x7f
    "01111111", -- 3770 - 0xeba  :  127 - 0x7f
    "00111111", -- 3771 - 0xebb  :   63 - 0x3f
    "00111111", -- 3772 - 0xebc  :   63 - 0x3f
    "00001111", -- 3773 - 0xebd  :   15 - 0xf
    "00000111", -- 3774 - 0xebe  :    7 - 0x7
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "11111111", -- 3776 - 0xec0  :  255 - 0xff -- Background 0xd8
    "11111111", -- 3777 - 0xec1  :  255 - 0xff
    "11111111", -- 3778 - 0xec2  :  255 - 0xff
    "11111111", -- 3779 - 0xec3  :  255 - 0xff
    "11111111", -- 3780 - 0xec4  :  255 - 0xff
    "11111111", -- 3781 - 0xec5  :  255 - 0xff
    "11111111", -- 3782 - 0xec6  :  255 - 0xff
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "11101010", -- 3784 - 0xec8  :  234 - 0xea -- Background 0xd9
    "11010100", -- 3785 - 0xec9  :  212 - 0xd4
    "11101010", -- 3786 - 0xeca  :  234 - 0xea
    "11010100", -- 3787 - 0xecb  :  212 - 0xd4
    "10101000", -- 3788 - 0xecc  :  168 - 0xa8
    "01010000", -- 3789 - 0xecd  :   80 - 0x50
    "10100000", -- 3790 - 0xece  :  160 - 0xa0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00001100", -- 3794 - 0xed2  :   12 - 0xc
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0 -- Background 0xdb
    "10000000", -- 3801 - 0xed9  :  128 - 0x80
    "10000000", -- 3802 - 0xeda  :  128 - 0x80
    "10000000", -- 3803 - 0xedb  :  128 - 0x80
    "10011000", -- 3804 - 0xedc  :  152 - 0x98
    "10000000", -- 3805 - 0xedd  :  128 - 0x80
    "10000000", -- 3806 - 0xede  :  128 - 0x80
    "10000000", -- 3807 - 0xedf  :  128 - 0x80
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000010", -- 3812 - 0xee4  :    2 - 0x2
    "00000011", -- 3813 - 0xee5  :    3 - 0x3
    "00000011", -- 3814 - 0xee6  :    3 - 0x3
    "00000001", -- 3815 - 0xee7  :    1 - 0x1
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "10100000", -- 3820 - 0xeec  :  160 - 0xa0
    "11100000", -- 3821 - 0xeed  :  224 - 0xe0
    "11100000", -- 3822 - 0xeee  :  224 - 0xe0
    "11000000", -- 3823 - 0xeef  :  192 - 0xc0
    "00110000", -- 3824 - 0xef0  :   48 - 0x30 -- Background 0xde
    "01111111", -- 3825 - 0xef1  :  127 - 0x7f
    "00110000", -- 3826 - 0xef2  :   48 - 0x30
    "00110000", -- 3827 - 0xef3  :   48 - 0x30
    "00110000", -- 3828 - 0xef4  :   48 - 0x30
    "00110000", -- 3829 - 0xef5  :   48 - 0x30
    "00110000", -- 3830 - 0xef6  :   48 - 0x30
    "00110000", -- 3831 - 0xef7  :   48 - 0x30
    "00001100", -- 3832 - 0xef8  :   12 - 0xc -- Background 0xdf
    "11111110", -- 3833 - 0xef9  :  254 - 0xfe
    "00001100", -- 3834 - 0xefa  :   12 - 0xc
    "00001100", -- 3835 - 0xefb  :   12 - 0xc
    "00001100", -- 3836 - 0xefc  :   12 - 0xc
    "00001100", -- 3837 - 0xefd  :   12 - 0xc
    "00001100", -- 3838 - 0xefe  :   12 - 0xc
    "00001100", -- 3839 - 0xeff  :   12 - 0xc
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- Background 0xe1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0 -- Background 0xe3
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000000", -- 3866 - 0xf1a  :    0 - 0x0
    "00000000", -- 3867 - 0xf1b  :    0 - 0x0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "00000000", -- 3880 - 0xf28  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000000", -- 3896 - 0xf38  :    0 - 0x0 -- Background 0xe7
    "00000000", -- 3897 - 0xf39  :    0 - 0x0
    "00000000", -- 3898 - 0xf3a  :    0 - 0x0
    "00000000", -- 3899 - 0xf3b  :    0 - 0x0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "00000000", -- 3915 - 0xf4b  :    0 - 0x0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Background 0xea
    "00000000", -- 3921 - 0xf51  :    0 - 0x0
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 3929 - 0xf59  :    0 - 0x0
    "00000000", -- 3930 - 0xf5a  :    0 - 0x0
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- Background 0xed
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0 -- Background 0xef
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00000000", -- 3976 - 0xf88  :    0 - 0x0 -- Background 0xf1
    "00000000", -- 3977 - 0xf89  :    0 - 0x0
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000000", -- 3979 - 0xf8b  :    0 - 0x0
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Background 0xf4
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- Background 0xf5
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- Background 0xf7
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "00000000", -- 4028 - 0xfbc  :    0 - 0x0
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00000000", -- 4030 - 0xfbe  :    0 - 0x0
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Background 0xf8
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "00000000", -- 4034 - 0xfc2  :    0 - 0x0
    "00000000", -- 4035 - 0xfc3  :    0 - 0x0
    "00000000", -- 4036 - 0xfc4  :    0 - 0x0
    "00000000", -- 4037 - 0xfc5  :    0 - 0x0
    "00000000", -- 4038 - 0xfc6  :    0 - 0x0
    "00000000", -- 4039 - 0xfc7  :    0 - 0x0
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0 -- Background 0xf9
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "00000000", -- 4053 - 0xfd5  :    0 - 0x0
    "00000000", -- 4054 - 0xfd6  :    0 - 0x0
    "00000000", -- 4055 - 0xfd7  :    0 - 0x0
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0 -- Background 0xfb
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "00000000", -- 4059 - 0xfdb  :    0 - 0x0
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "00000000", -- 4069 - 0xfe5  :    0 - 0x0
    "00000000", -- 4070 - 0xfe6  :    0 - 0x0
    "00000000", -- 4071 - 0xfe7  :    0 - 0x0
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "00000000", -- 4075 - 0xfeb  :    0 - 0x0
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "00000000", -- 4082 - 0xff2  :    0 - 0x0
    "00000000", -- 4083 - 0xff3  :    0 - 0x0
    "00000000", -- 4084 - 0xff4  :    0 - 0x0
    "00000000", -- 4085 - 0xff5  :    0 - 0x0
    "00000000", -- 4086 - 0xff6  :    0 - 0x0
    "00000000", -- 4087 - 0xff7  :    0 - 0x0
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
