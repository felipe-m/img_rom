//-   Background Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_DONKEYKONG_BG
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table both color planes
      12'h0: dout <= 8'b00111000; //    0 :  56 - 0x38 -- Background 0x0
      12'h1: dout <= 8'b01001100; //    1 :  76 - 0x4c
      12'h2: dout <= 8'b11000110; //    2 : 198 - 0xc6
      12'h3: dout <= 8'b11000110; //    3 : 198 - 0xc6
      12'h4: dout <= 8'b11000110; //    4 : 198 - 0xc6
      12'h5: dout <= 8'b01100100; //    5 : 100 - 0x64
      12'h6: dout <= 8'b00111000; //    6 :  56 - 0x38
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b00011000; //   16 :  24 - 0x18 -- Background 0x1
      12'h11: dout <= 8'b00111000; //   17 :  56 - 0x38
      12'h12: dout <= 8'b00011000; //   18 :  24 - 0x18
      12'h13: dout <= 8'b00011000; //   19 :  24 - 0x18
      12'h14: dout <= 8'b00011000; //   20 :  24 - 0x18
      12'h15: dout <= 8'b00011000; //   21 :  24 - 0x18
      12'h16: dout <= 8'b01111110; //   22 : 126 - 0x7e
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout <= 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b01111100; //   32 : 124 - 0x7c -- Background 0x2
      12'h21: dout <= 8'b11000110; //   33 : 198 - 0xc6
      12'h22: dout <= 8'b00001110; //   34 :  14 - 0xe
      12'h23: dout <= 8'b00111100; //   35 :  60 - 0x3c
      12'h24: dout <= 8'b01111000; //   36 : 120 - 0x78
      12'h25: dout <= 8'b11100000; //   37 : 224 - 0xe0
      12'h26: dout <= 8'b11111110; //   38 : 254 - 0xfe
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b01111110; //   48 : 126 - 0x7e -- Background 0x3
      12'h31: dout <= 8'b00001100; //   49 :  12 - 0xc
      12'h32: dout <= 8'b00011000; //   50 :  24 - 0x18
      12'h33: dout <= 8'b00111100; //   51 :  60 - 0x3c
      12'h34: dout <= 8'b00000110; //   52 :   6 - 0x6
      12'h35: dout <= 8'b11000110; //   53 : 198 - 0xc6
      12'h36: dout <= 8'b01111100; //   54 : 124 - 0x7c
      12'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b00011100; //   64 :  28 - 0x1c -- Background 0x4
      12'h41: dout <= 8'b00111100; //   65 :  60 - 0x3c
      12'h42: dout <= 8'b01101100; //   66 : 108 - 0x6c
      12'h43: dout <= 8'b11001100; //   67 : 204 - 0xcc
      12'h44: dout <= 8'b11111110; //   68 : 254 - 0xfe
      12'h45: dout <= 8'b00001100; //   69 :  12 - 0xc
      12'h46: dout <= 8'b00001100; //   70 :  12 - 0xc
      12'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- plane 1
      12'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout <= 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout <= 8'b11111100; //   80 : 252 - 0xfc -- Background 0x5
      12'h51: dout <= 8'b11000000; //   81 : 192 - 0xc0
      12'h52: dout <= 8'b11111100; //   82 : 252 - 0xfc
      12'h53: dout <= 8'b00000110; //   83 :   6 - 0x6
      12'h54: dout <= 8'b00000110; //   84 :   6 - 0x6
      12'h55: dout <= 8'b11000110; //   85 : 198 - 0xc6
      12'h56: dout <= 8'b01111100; //   86 : 124 - 0x7c
      12'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- plane 1
      12'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b00111100; //   96 :  60 - 0x3c -- Background 0x6
      12'h61: dout <= 8'b01100000; //   97 :  96 - 0x60
      12'h62: dout <= 8'b11000000; //   98 : 192 - 0xc0
      12'h63: dout <= 8'b11111100; //   99 : 252 - 0xfc
      12'h64: dout <= 8'b11000110; //  100 : 198 - 0xc6
      12'h65: dout <= 8'b11000110; //  101 : 198 - 0xc6
      12'h66: dout <= 8'b01111100; //  102 : 124 - 0x7c
      12'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- plane 1
      12'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout <= 8'b11111110; //  112 : 254 - 0xfe -- Background 0x7
      12'h71: dout <= 8'b11000110; //  113 : 198 - 0xc6
      12'h72: dout <= 8'b00001100; //  114 :  12 - 0xc
      12'h73: dout <= 8'b00011000; //  115 :  24 - 0x18
      12'h74: dout <= 8'b00110000; //  116 :  48 - 0x30
      12'h75: dout <= 8'b00110000; //  117 :  48 - 0x30
      12'h76: dout <= 8'b00110000; //  118 :  48 - 0x30
      12'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- plane 1
      12'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b01111000; //  128 : 120 - 0x78 -- Background 0x8
      12'h81: dout <= 8'b11000100; //  129 : 196 - 0xc4
      12'h82: dout <= 8'b11100100; //  130 : 228 - 0xe4
      12'h83: dout <= 8'b01111000; //  131 : 120 - 0x78
      12'h84: dout <= 8'b10000110; //  132 : 134 - 0x86
      12'h85: dout <= 8'b10000110; //  133 : 134 - 0x86
      12'h86: dout <= 8'b01111100; //  134 : 124 - 0x7c
      12'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout <= 8'b01111100; //  144 : 124 - 0x7c -- Background 0x9
      12'h91: dout <= 8'b11000110; //  145 : 198 - 0xc6
      12'h92: dout <= 8'b11000110; //  146 : 198 - 0xc6
      12'h93: dout <= 8'b01111110; //  147 : 126 - 0x7e
      12'h94: dout <= 8'b00000110; //  148 :   6 - 0x6
      12'h95: dout <= 8'b00001100; //  149 :  12 - 0xc
      12'h96: dout <= 8'b01111000; //  150 : 120 - 0x78
      12'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- plane 1
      12'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b00111000; //  160 :  56 - 0x38 -- Background 0xa
      12'hA1: dout <= 8'b01101100; //  161 : 108 - 0x6c
      12'hA2: dout <= 8'b11000110; //  162 : 198 - 0xc6
      12'hA3: dout <= 8'b11000110; //  163 : 198 - 0xc6
      12'hA4: dout <= 8'b11111110; //  164 : 254 - 0xfe
      12'hA5: dout <= 8'b11000110; //  165 : 198 - 0xc6
      12'hA6: dout <= 8'b11000110; //  166 : 198 - 0xc6
      12'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- plane 1
      12'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      12'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b11111100; //  176 : 252 - 0xfc -- Background 0xb
      12'hB1: dout <= 8'b11000110; //  177 : 198 - 0xc6
      12'hB2: dout <= 8'b11000110; //  178 : 198 - 0xc6
      12'hB3: dout <= 8'b11111100; //  179 : 252 - 0xfc
      12'hB4: dout <= 8'b11000110; //  180 : 198 - 0xc6
      12'hB5: dout <= 8'b11000110; //  181 : 198 - 0xc6
      12'hB6: dout <= 8'b11111100; //  182 : 252 - 0xfc
      12'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- plane 1
      12'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      12'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      12'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b00111100; //  192 :  60 - 0x3c -- Background 0xc
      12'hC1: dout <= 8'b01100110; //  193 : 102 - 0x66
      12'hC2: dout <= 8'b11000000; //  194 : 192 - 0xc0
      12'hC3: dout <= 8'b11000000; //  195 : 192 - 0xc0
      12'hC4: dout <= 8'b11000000; //  196 : 192 - 0xc0
      12'hC5: dout <= 8'b01100110; //  197 : 102 - 0x66
      12'hC6: dout <= 8'b00111100; //  198 :  60 - 0x3c
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- plane 1
      12'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      12'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      12'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b11111000; //  208 : 248 - 0xf8 -- Background 0xd
      12'hD1: dout <= 8'b11001100; //  209 : 204 - 0xcc
      12'hD2: dout <= 8'b11000110; //  210 : 198 - 0xc6
      12'hD3: dout <= 8'b11000110; //  211 : 198 - 0xc6
      12'hD4: dout <= 8'b11000110; //  212 : 198 - 0xc6
      12'hD5: dout <= 8'b11001100; //  213 : 204 - 0xcc
      12'hD6: dout <= 8'b11111000; //  214 : 248 - 0xf8
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- plane 1
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      12'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      12'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b11111110; //  224 : 254 - 0xfe -- Background 0xe
      12'hE1: dout <= 8'b11000000; //  225 : 192 - 0xc0
      12'hE2: dout <= 8'b11000000; //  226 : 192 - 0xc0
      12'hE3: dout <= 8'b11111100; //  227 : 252 - 0xfc
      12'hE4: dout <= 8'b11000000; //  228 : 192 - 0xc0
      12'hE5: dout <= 8'b11000000; //  229 : 192 - 0xc0
      12'hE6: dout <= 8'b11111110; //  230 : 254 - 0xfe
      12'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- plane 1
      12'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      12'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      12'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout <= 8'b11111110; //  240 : 254 - 0xfe -- Background 0xf
      12'hF1: dout <= 8'b11000000; //  241 : 192 - 0xc0
      12'hF2: dout <= 8'b11000000; //  242 : 192 - 0xc0
      12'hF3: dout <= 8'b11111100; //  243 : 252 - 0xfc
      12'hF4: dout <= 8'b11000000; //  244 : 192 - 0xc0
      12'hF5: dout <= 8'b11000000; //  245 : 192 - 0xc0
      12'hF6: dout <= 8'b11000000; //  246 : 192 - 0xc0
      12'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00111110; //  256 :  62 - 0x3e -- Background 0x10
      12'h101: dout <= 8'b01100000; //  257 :  96 - 0x60
      12'h102: dout <= 8'b11000000; //  258 : 192 - 0xc0
      12'h103: dout <= 8'b11011110; //  259 : 222 - 0xde
      12'h104: dout <= 8'b11000110; //  260 : 198 - 0xc6
      12'h105: dout <= 8'b01100110; //  261 : 102 - 0x66
      12'h106: dout <= 8'b01111110; //  262 : 126 - 0x7e
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b11000110; //  272 : 198 - 0xc6 -- Background 0x11
      12'h111: dout <= 8'b11000110; //  273 : 198 - 0xc6
      12'h112: dout <= 8'b11000110; //  274 : 198 - 0xc6
      12'h113: dout <= 8'b11111110; //  275 : 254 - 0xfe
      12'h114: dout <= 8'b11000110; //  276 : 198 - 0xc6
      12'h115: dout <= 8'b11000110; //  277 : 198 - 0xc6
      12'h116: dout <= 8'b11000110; //  278 : 198 - 0xc6
      12'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      12'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b01111110; //  288 : 126 - 0x7e -- Background 0x12
      12'h121: dout <= 8'b00011000; //  289 :  24 - 0x18
      12'h122: dout <= 8'b00011000; //  290 :  24 - 0x18
      12'h123: dout <= 8'b00011000; //  291 :  24 - 0x18
      12'h124: dout <= 8'b00011000; //  292 :  24 - 0x18
      12'h125: dout <= 8'b00011000; //  293 :  24 - 0x18
      12'h126: dout <= 8'b01111110; //  294 : 126 - 0x7e
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      12'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      12'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout <= 8'b00011110; //  304 :  30 - 0x1e -- Background 0x13
      12'h131: dout <= 8'b00000110; //  305 :   6 - 0x6
      12'h132: dout <= 8'b00000110; //  306 :   6 - 0x6
      12'h133: dout <= 8'b00000110; //  307 :   6 - 0x6
      12'h134: dout <= 8'b11000110; //  308 : 198 - 0xc6
      12'h135: dout <= 8'b11000110; //  309 : 198 - 0xc6
      12'h136: dout <= 8'b01111100; //  310 : 124 - 0x7c
      12'h137: dout <= 8'b00000000; //  311 :   0 - 0x0
      12'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- plane 1
      12'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b11000110; //  320 : 198 - 0xc6 -- Background 0x14
      12'h141: dout <= 8'b11001100; //  321 : 204 - 0xcc
      12'h142: dout <= 8'b11011000; //  322 : 216 - 0xd8
      12'h143: dout <= 8'b11110000; //  323 : 240 - 0xf0
      12'h144: dout <= 8'b11111000; //  324 : 248 - 0xf8
      12'h145: dout <= 8'b11011100; //  325 : 220 - 0xdc
      12'h146: dout <= 8'b11001110; //  326 : 206 - 0xce
      12'h147: dout <= 8'b00000000; //  327 :   0 - 0x0
      12'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- plane 1
      12'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      12'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout <= 8'b01100000; //  336 :  96 - 0x60 -- Background 0x15
      12'h151: dout <= 8'b01100000; //  337 :  96 - 0x60
      12'h152: dout <= 8'b01100000; //  338 :  96 - 0x60
      12'h153: dout <= 8'b01100000; //  339 :  96 - 0x60
      12'h154: dout <= 8'b01100000; //  340 :  96 - 0x60
      12'h155: dout <= 8'b01100000; //  341 :  96 - 0x60
      12'h156: dout <= 8'b01111110; //  342 : 126 - 0x7e
      12'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- plane 1
      12'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b11000110; //  352 : 198 - 0xc6 -- Background 0x16
      12'h161: dout <= 8'b11101110; //  353 : 238 - 0xee
      12'h162: dout <= 8'b11111110; //  354 : 254 - 0xfe
      12'h163: dout <= 8'b11111110; //  355 : 254 - 0xfe
      12'h164: dout <= 8'b11010110; //  356 : 214 - 0xd6
      12'h165: dout <= 8'b11000110; //  357 : 198 - 0xc6
      12'h166: dout <= 8'b11000110; //  358 : 198 - 0xc6
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- plane 1
      12'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout <= 8'b11000110; //  368 : 198 - 0xc6 -- Background 0x17
      12'h171: dout <= 8'b11100110; //  369 : 230 - 0xe6
      12'h172: dout <= 8'b11110110; //  370 : 246 - 0xf6
      12'h173: dout <= 8'b11111110; //  371 : 254 - 0xfe
      12'h174: dout <= 8'b11011110; //  372 : 222 - 0xde
      12'h175: dout <= 8'b11001110; //  373 : 206 - 0xce
      12'h176: dout <= 8'b11000110; //  374 : 198 - 0xc6
      12'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- plane 1
      12'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      12'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b01111100; //  384 : 124 - 0x7c -- Background 0x18
      12'h181: dout <= 8'b11000110; //  385 : 198 - 0xc6
      12'h182: dout <= 8'b11000110; //  386 : 198 - 0xc6
      12'h183: dout <= 8'b11000110; //  387 : 198 - 0xc6
      12'h184: dout <= 8'b11000110; //  388 : 198 - 0xc6
      12'h185: dout <= 8'b11000110; //  389 : 198 - 0xc6
      12'h186: dout <= 8'b01111100; //  390 : 124 - 0x7c
      12'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      12'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      12'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      12'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b11111100; //  400 : 252 - 0xfc -- Background 0x19
      12'h191: dout <= 8'b11000110; //  401 : 198 - 0xc6
      12'h192: dout <= 8'b11000110; //  402 : 198 - 0xc6
      12'h193: dout <= 8'b11000110; //  403 : 198 - 0xc6
      12'h194: dout <= 8'b11111100; //  404 : 252 - 0xfc
      12'h195: dout <= 8'b11000000; //  405 : 192 - 0xc0
      12'h196: dout <= 8'b11000000; //  406 : 192 - 0xc0
      12'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout <= 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout <= 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout <= 8'b00000000; //  412 :   0 - 0x0
      12'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b01111100; //  416 : 124 - 0x7c -- Background 0x1a
      12'h1A1: dout <= 8'b11000110; //  417 : 198 - 0xc6
      12'h1A2: dout <= 8'b11000110; //  418 : 198 - 0xc6
      12'h1A3: dout <= 8'b11000110; //  419 : 198 - 0xc6
      12'h1A4: dout <= 8'b11011110; //  420 : 222 - 0xde
      12'h1A5: dout <= 8'b11001100; //  421 : 204 - 0xcc
      12'h1A6: dout <= 8'b01111010; //  422 : 122 - 0x7a
      12'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0 -- plane 1
      12'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      12'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b11111100; //  432 : 252 - 0xfc -- Background 0x1b
      12'h1B1: dout <= 8'b11000110; //  433 : 198 - 0xc6
      12'h1B2: dout <= 8'b11000110; //  434 : 198 - 0xc6
      12'h1B3: dout <= 8'b11001110; //  435 : 206 - 0xce
      12'h1B4: dout <= 8'b11111000; //  436 : 248 - 0xf8
      12'h1B5: dout <= 8'b11011100; //  437 : 220 - 0xdc
      12'h1B6: dout <= 8'b11001110; //  438 : 206 - 0xce
      12'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      12'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      12'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b01111000; //  448 : 120 - 0x78 -- Background 0x1c
      12'h1C1: dout <= 8'b11001100; //  449 : 204 - 0xcc
      12'h1C2: dout <= 8'b11000000; //  450 : 192 - 0xc0
      12'h1C3: dout <= 8'b01111100; //  451 : 124 - 0x7c
      12'h1C4: dout <= 8'b00000110; //  452 :   6 - 0x6
      12'h1C5: dout <= 8'b11000110; //  453 : 198 - 0xc6
      12'h1C6: dout <= 8'b01111100; //  454 : 124 - 0x7c
      12'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- plane 1
      12'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b01111110; //  464 : 126 - 0x7e -- Background 0x1d
      12'h1D1: dout <= 8'b00011000; //  465 :  24 - 0x18
      12'h1D2: dout <= 8'b00011000; //  466 :  24 - 0x18
      12'h1D3: dout <= 8'b00011000; //  467 :  24 - 0x18
      12'h1D4: dout <= 8'b00011000; //  468 :  24 - 0x18
      12'h1D5: dout <= 8'b00011000; //  469 :  24 - 0x18
      12'h1D6: dout <= 8'b00011000; //  470 :  24 - 0x18
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- plane 1
      12'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b11000110; //  480 : 198 - 0xc6 -- Background 0x1e
      12'h1E1: dout <= 8'b11000110; //  481 : 198 - 0xc6
      12'h1E2: dout <= 8'b11000110; //  482 : 198 - 0xc6
      12'h1E3: dout <= 8'b11000110; //  483 : 198 - 0xc6
      12'h1E4: dout <= 8'b11000110; //  484 : 198 - 0xc6
      12'h1E5: dout <= 8'b11000110; //  485 : 198 - 0xc6
      12'h1E6: dout <= 8'b01111100; //  486 : 124 - 0x7c
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- plane 1
      12'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b11000110; //  496 : 198 - 0xc6 -- Background 0x1f
      12'h1F1: dout <= 8'b11000110; //  497 : 198 - 0xc6
      12'h1F2: dout <= 8'b11000110; //  498 : 198 - 0xc6
      12'h1F3: dout <= 8'b11101110; //  499 : 238 - 0xee
      12'h1F4: dout <= 8'b01111100; //  500 : 124 - 0x7c
      12'h1F5: dout <= 8'b00111000; //  501 :  56 - 0x38
      12'h1F6: dout <= 8'b00010000; //  502 :  16 - 0x10
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- plane 1
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b11000110; //  512 : 198 - 0xc6 -- Background 0x20
      12'h201: dout <= 8'b11000110; //  513 : 198 - 0xc6
      12'h202: dout <= 8'b11010110; //  514 : 214 - 0xd6
      12'h203: dout <= 8'b11111110; //  515 : 254 - 0xfe
      12'h204: dout <= 8'b11111110; //  516 : 254 - 0xfe
      12'h205: dout <= 8'b11101110; //  517 : 238 - 0xee
      12'h206: dout <= 8'b11000110; //  518 : 198 - 0xc6
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b11000110; //  528 : 198 - 0xc6 -- Background 0x21
      12'h211: dout <= 8'b11101110; //  529 : 238 - 0xee
      12'h212: dout <= 8'b01111100; //  530 : 124 - 0x7c
      12'h213: dout <= 8'b00111000; //  531 :  56 - 0x38
      12'h214: dout <= 8'b01111100; //  532 : 124 - 0x7c
      12'h215: dout <= 8'b11101110; //  533 : 238 - 0xee
      12'h216: dout <= 8'b11000110; //  534 : 198 - 0xc6
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b01100110; //  544 : 102 - 0x66 -- Background 0x22
      12'h221: dout <= 8'b01100110; //  545 : 102 - 0x66
      12'h222: dout <= 8'b01100110; //  546 : 102 - 0x66
      12'h223: dout <= 8'b00111100; //  547 :  60 - 0x3c
      12'h224: dout <= 8'b00011000; //  548 :  24 - 0x18
      12'h225: dout <= 8'b00011000; //  549 :  24 - 0x18
      12'h226: dout <= 8'b00011000; //  550 :  24 - 0x18
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b00000000; //  552 :   0 - 0x0 -- plane 1
      12'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      12'h22A: dout <= 8'b00000000; //  554 :   0 - 0x0
      12'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      12'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      12'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b11111110; //  560 : 254 - 0xfe -- Background 0x23
      12'h231: dout <= 8'b00001110; //  561 :  14 - 0xe
      12'h232: dout <= 8'b00011100; //  562 :  28 - 0x1c
      12'h233: dout <= 8'b00111000; //  563 :  56 - 0x38
      12'h234: dout <= 8'b01110000; //  564 : 112 - 0x70
      12'h235: dout <= 8'b11100000; //  565 : 224 - 0xe0
      12'h236: dout <= 8'b11111110; //  566 : 254 - 0xfe
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- plane 1
      12'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Background 0x24
      12'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      12'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      12'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      12'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- plane 1
      12'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00000000; //  592 :   0 - 0x0 -- Background 0x25
      12'h251: dout <= 8'b00000000; //  593 :   0 - 0x0
      12'h252: dout <= 8'b00000110; //  594 :   6 - 0x6
      12'h253: dout <= 8'b00001110; //  595 :  14 - 0xe
      12'h254: dout <= 8'b00001000; //  596 :   8 - 0x8
      12'h255: dout <= 8'b00001000; //  597 :   8 - 0x8
      12'h256: dout <= 8'b00001000; //  598 :   8 - 0x8
      12'h257: dout <= 8'b00001000; //  599 :   8 - 0x8
      12'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- plane 1
      12'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout <= 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout <= 8'b00000000; //  605 :   0 - 0x0
      12'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Background 0x26
      12'h261: dout <= 8'b01111000; //  609 : 120 - 0x78
      12'h262: dout <= 8'b01100101; //  610 : 101 - 0x65
      12'h263: dout <= 8'b01111001; //  611 : 121 - 0x79
      12'h264: dout <= 8'b01100101; //  612 : 101 - 0x65
      12'h265: dout <= 8'b01100101; //  613 : 101 - 0x65
      12'h266: dout <= 8'b01111000; //  614 : 120 - 0x78
      12'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- plane 1
      12'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout <= 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b00000000; //  621 :   0 - 0x0
      12'h26E: dout <= 8'b00000000; //  622 :   0 - 0x0
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Background 0x27
      12'h271: dout <= 8'b11100100; //  625 : 228 - 0xe4
      12'h272: dout <= 8'b10010110; //  626 : 150 - 0x96
      12'h273: dout <= 8'b10010110; //  627 : 150 - 0x96
      12'h274: dout <= 8'b10010111; //  628 : 151 - 0x97
      12'h275: dout <= 8'b10010110; //  629 : 150 - 0x96
      12'h276: dout <= 8'b11100110; //  630 : 230 - 0xe6
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00000000; //  632 :   0 - 0x0 -- plane 1
      12'h279: dout <= 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout <= 8'b00000000; //  634 :   0 - 0x0
      12'h27B: dout <= 8'b00000000; //  635 :   0 - 0x0
      12'h27C: dout <= 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout <= 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout <= 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Background 0x28
      12'h281: dout <= 8'b01011001; //  641 :  89 - 0x59
      12'h282: dout <= 8'b01011001; //  642 :  89 - 0x59
      12'h283: dout <= 8'b01011001; //  643 :  89 - 0x59
      12'h284: dout <= 8'b01011001; //  644 :  89 - 0x59
      12'h285: dout <= 8'b11011001; //  645 : 217 - 0xd9
      12'h286: dout <= 8'b01001110; //  646 :  78 - 0x4e
      12'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout <= 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout <= 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout <= 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout <= 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Background 0x29
      12'h291: dout <= 8'b00111100; //  657 :  60 - 0x3c
      12'h292: dout <= 8'b01110000; //  658 : 112 - 0x70
      12'h293: dout <= 8'b01110000; //  659 : 112 - 0x70
      12'h294: dout <= 8'b00111100; //  660 :  60 - 0x3c
      12'h295: dout <= 8'b00001100; //  661 :  12 - 0xc
      12'h296: dout <= 8'b01111000; //  662 : 120 - 0x78
      12'h297: dout <= 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- plane 1
      12'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout <= 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout <= 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout <= 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout <= 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout <= 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Background 0x2a
      12'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      12'h2A2: dout <= 8'b11000110; //  674 : 198 - 0xc6
      12'h2A3: dout <= 8'b11101110; //  675 : 238 - 0xee
      12'h2A4: dout <= 8'b00101000; //  676 :  40 - 0x28
      12'h2A5: dout <= 8'b00101000; //  677 :  40 - 0x28
      12'h2A6: dout <= 8'b00101000; //  678 :  40 - 0x28
      12'h2A7: dout <= 8'b00101000; //  679 :  40 - 0x28
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- plane 1
      12'h2A9: dout <= 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout <= 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout <= 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout <= 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout <= 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout <= 8'b00000000; //  686 :   0 - 0x0
      12'h2AF: dout <= 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout <= 8'b00001000; //  688 :   8 - 0x8 -- Background 0x2b
      12'h2B1: dout <= 8'b00001000; //  689 :   8 - 0x8
      12'h2B2: dout <= 8'b00001000; //  690 :   8 - 0x8
      12'h2B3: dout <= 8'b00001000; //  691 :   8 - 0x8
      12'h2B4: dout <= 8'b00001110; //  692 :  14 - 0xe
      12'h2B5: dout <= 8'b00000110; //  693 :   6 - 0x6
      12'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- plane 1
      12'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b00101000; //  704 :  40 - 0x28 -- Background 0x2c
      12'h2C1: dout <= 8'b00101000; //  705 :  40 - 0x28
      12'h2C2: dout <= 8'b00101000; //  706 :  40 - 0x28
      12'h2C3: dout <= 8'b00101000; //  707 :  40 - 0x28
      12'h2C4: dout <= 8'b11101110; //  708 : 238 - 0xee
      12'h2C5: dout <= 8'b11000110; //  709 : 198 - 0xc6
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Background 0x2d
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b01100000; //  722 :  96 - 0x60
      12'h2D3: dout <= 8'b01110000; //  723 : 112 - 0x70
      12'h2D4: dout <= 8'b00010000; //  724 :  16 - 0x10
      12'h2D5: dout <= 8'b00010000; //  725 :  16 - 0x10
      12'h2D6: dout <= 8'b00010000; //  726 :  16 - 0x10
      12'h2D7: dout <= 8'b00010000; //  727 :  16 - 0x10
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- plane 1
      12'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      12'h2DD: dout <= 8'b00000000; //  733 :   0 - 0x0
      12'h2DE: dout <= 8'b00000000; //  734 :   0 - 0x0
      12'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout <= 8'b00011100; //  736 :  28 - 0x1c -- Background 0x2e
      12'h2E1: dout <= 8'b00111110; //  737 :  62 - 0x3e
      12'h2E2: dout <= 8'b00111100; //  738 :  60 - 0x3c
      12'h2E3: dout <= 8'b00111000; //  739 :  56 - 0x38
      12'h2E4: dout <= 8'b00110000; //  740 :  48 - 0x30
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b01100000; //  742 :  96 - 0x60
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout <= 8'b00010000; //  752 :  16 - 0x10 -- Background 0x2f
      12'h2F1: dout <= 8'b00010000; //  753 :  16 - 0x10
      12'h2F2: dout <= 8'b00010000; //  754 :  16 - 0x10
      12'h2F3: dout <= 8'b00010000; //  755 :  16 - 0x10
      12'h2F4: dout <= 8'b01110000; //  756 : 112 - 0x70
      12'h2F5: dout <= 8'b01100000; //  757 :  96 - 0x60
      12'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- plane 1
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b00000000; //  763 :   0 - 0x0
      12'h2FC: dout <= 8'b00000000; //  764 :   0 - 0x0
      12'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b11111111; //  768 : 255 - 0xff -- Background 0x30
      12'h301: dout <= 8'b11111111; //  769 : 255 - 0xff
      12'h302: dout <= 8'b00111000; //  770 :  56 - 0x38
      12'h303: dout <= 8'b01101100; //  771 : 108 - 0x6c
      12'h304: dout <= 8'b11000110; //  772 : 198 - 0xc6
      12'h305: dout <= 8'b10000011; //  773 : 131 - 0x83
      12'h306: dout <= 8'b11111111; //  774 : 255 - 0xff
      12'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- plane 1
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      12'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      12'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      12'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      12'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b11111111; //  784 : 255 - 0xff -- Background 0x31
      12'h311: dout <= 8'b00111000; //  785 :  56 - 0x38
      12'h312: dout <= 8'b01101100; //  786 : 108 - 0x6c
      12'h313: dout <= 8'b11000110; //  787 : 198 - 0xc6
      12'h314: dout <= 8'b10000011; //  788 : 131 - 0x83
      12'h315: dout <= 8'b11111111; //  789 : 255 - 0xff
      12'h316: dout <= 8'b11111111; //  790 : 255 - 0xff
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00111000; //  800 :  56 - 0x38 -- Background 0x32
      12'h321: dout <= 8'b01101100; //  801 : 108 - 0x6c
      12'h322: dout <= 8'b11000110; //  802 : 198 - 0xc6
      12'h323: dout <= 8'b10000011; //  803 : 131 - 0x83
      12'h324: dout <= 8'b11111111; //  804 : 255 - 0xff
      12'h325: dout <= 8'b11111111; //  805 : 255 - 0xff
      12'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout <= 8'b01101100; //  816 : 108 - 0x6c -- Background 0x33
      12'h331: dout <= 8'b11000110; //  817 : 198 - 0xc6
      12'h332: dout <= 8'b10000011; //  818 : 131 - 0x83
      12'h333: dout <= 8'b11111111; //  819 : 255 - 0xff
      12'h334: dout <= 8'b11111111; //  820 : 255 - 0xff
      12'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- plane 1
      12'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b11000110; //  832 : 198 - 0xc6 -- Background 0x34
      12'h341: dout <= 8'b10000011; //  833 : 131 - 0x83
      12'h342: dout <= 8'b11111111; //  834 : 255 - 0xff
      12'h343: dout <= 8'b11111111; //  835 : 255 - 0xff
      12'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b10000011; //  848 : 131 - 0x83 -- Background 0x35
      12'h351: dout <= 8'b11111111; //  849 : 255 - 0xff
      12'h352: dout <= 8'b11111111; //  850 : 255 - 0xff
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- plane 1
      12'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- Background 0x36
      12'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      12'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b11111111; //  880 : 255 - 0xff -- Background 0x37
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b00000000; //  888 :   0 - 0x0 -- plane 1
      12'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Background 0x38
      12'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Background 0x39
      12'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      12'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      12'h398: dout <= 8'b00000000; //  920 :   0 - 0x0 -- plane 1
      12'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Background 0x3a
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b11111111; //  933 : 255 - 0xff
      12'h3A6: dout <= 8'b11111111; //  934 : 255 - 0xff
      12'h3A7: dout <= 8'b00111000; //  935 :  56 - 0x38
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Background 0x3b
      12'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout <= 8'b11111111; //  948 : 255 - 0xff
      12'h3B5: dout <= 8'b11111111; //  949 : 255 - 0xff
      12'h3B6: dout <= 8'b00111000; //  950 :  56 - 0x38
      12'h3B7: dout <= 8'b01101100; //  951 : 108 - 0x6c
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Background 0x3c
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      12'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      12'h3C5: dout <= 8'b00111000; //  965 :  56 - 0x38
      12'h3C6: dout <= 8'b01101100; //  966 : 108 - 0x6c
      12'h3C7: dout <= 8'b11000110; //  967 : 198 - 0xc6
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Background 0x3d
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      12'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      12'h3D4: dout <= 8'b00111000; //  980 :  56 - 0x38
      12'h3D5: dout <= 8'b01101100; //  981 : 108 - 0x6c
      12'h3D6: dout <= 8'b11000110; //  982 : 198 - 0xc6
      12'h3D7: dout <= 8'b10000011; //  983 : 131 - 0x83
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Background 0x3e
      12'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      12'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      12'h3E3: dout <= 8'b00111000; //  995 :  56 - 0x38
      12'h3E4: dout <= 8'b01101100; //  996 : 108 - 0x6c
      12'h3E5: dout <= 8'b11000110; //  997 : 198 - 0xc6
      12'h3E6: dout <= 8'b10000011; //  998 : 131 - 0x83
      12'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout <= 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout <= 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout <= 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x3f
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b10000001; // 1016 : 129 - 0x81 -- plane 1
      12'h3F9: dout <= 8'b11111111; // 1017 : 255 - 0xff
      12'h3FA: dout <= 8'b10000001; // 1018 : 129 - 0x81
      12'h3FB: dout <= 8'b10000001; // 1019 : 129 - 0x81
      12'h3FC: dout <= 8'b10000001; // 1020 : 129 - 0x81
      12'h3FD: dout <= 8'b11111111; // 1021 : 255 - 0xff
      12'h3FE: dout <= 8'b10000001; // 1022 : 129 - 0x81
      12'h3FF: dout <= 8'b10000001; // 1023 : 129 - 0x81
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Background 0x40
      12'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout <= 8'b11111111; // 1031 : 255 - 0xff
      12'h408: dout <= 8'b10000001; // 1032 : 129 - 0x81 -- plane 1
      12'h409: dout <= 8'b11111111; // 1033 : 255 - 0xff
      12'h40A: dout <= 8'b10000001; // 1034 : 129 - 0x81
      12'h40B: dout <= 8'b10000001; // 1035 : 129 - 0x81
      12'h40C: dout <= 8'b10000001; // 1036 : 129 - 0x81
      12'h40D: dout <= 8'b11111111; // 1037 : 255 - 0xff
      12'h40E: dout <= 8'b10000001; // 1038 : 129 - 0x81
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x41
      12'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      12'h415: dout <= 8'b11111111; // 1045 : 255 - 0xff
      12'h416: dout <= 8'b11111111; // 1046 : 255 - 0xff
      12'h417: dout <= 8'b00111000; // 1047 :  56 - 0x38
      12'h418: dout <= 8'b10000001; // 1048 : 129 - 0x81 -- plane 1
      12'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout <= 8'b10000001; // 1050 : 129 - 0x81
      12'h41B: dout <= 8'b10000001; // 1051 : 129 - 0x81
      12'h41C: dout <= 8'b10000001; // 1052 : 129 - 0x81
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Background 0x42
      12'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      12'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      12'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout <= 8'b11111111; // 1060 : 255 - 0xff
      12'h425: dout <= 8'b11111111; // 1061 : 255 - 0xff
      12'h426: dout <= 8'b00111000; // 1062 :  56 - 0x38
      12'h427: dout <= 8'b01101100; // 1063 : 108 - 0x6c
      12'h428: dout <= 8'b10000001; // 1064 : 129 - 0x81 -- plane 1
      12'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      12'h42A: dout <= 8'b10000001; // 1066 : 129 - 0x81
      12'h42B: dout <= 8'b10000001; // 1067 : 129 - 0x81
      12'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x43
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b11111111; // 1075 : 255 - 0xff
      12'h434: dout <= 8'b11111111; // 1076 : 255 - 0xff
      12'h435: dout <= 8'b00111000; // 1077 :  56 - 0x38
      12'h436: dout <= 8'b01101100; // 1078 : 108 - 0x6c
      12'h437: dout <= 8'b11000110; // 1079 : 198 - 0xc6
      12'h438: dout <= 8'b10000001; // 1080 : 129 - 0x81 -- plane 1
      12'h439: dout <= 8'b11111111; // 1081 : 255 - 0xff
      12'h43A: dout <= 8'b10000001; // 1082 : 129 - 0x81
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x44
      12'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      12'h442: dout <= 8'b11111111; // 1090 : 255 - 0xff
      12'h443: dout <= 8'b11111111; // 1091 : 255 - 0xff
      12'h444: dout <= 8'b00111000; // 1092 :  56 - 0x38
      12'h445: dout <= 8'b01101100; // 1093 : 108 - 0x6c
      12'h446: dout <= 8'b11000110; // 1094 : 198 - 0xc6
      12'h447: dout <= 8'b10000011; // 1095 : 131 - 0x83
      12'h448: dout <= 8'b10000001; // 1096 : 129 - 0x81 -- plane 1
      12'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      12'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      12'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x45
      12'h451: dout <= 8'b11111111; // 1105 : 255 - 0xff
      12'h452: dout <= 8'b11111111; // 1106 : 255 - 0xff
      12'h453: dout <= 8'b00111000; // 1107 :  56 - 0x38
      12'h454: dout <= 8'b01101100; // 1108 : 108 - 0x6c
      12'h455: dout <= 8'b11000110; // 1109 : 198 - 0xc6
      12'h456: dout <= 8'b10000011; // 1110 : 131 - 0x83
      12'h457: dout <= 8'b11111111; // 1111 : 255 - 0xff
      12'h458: dout <= 8'b10000001; // 1112 : 129 - 0x81 -- plane 1
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b11111111; // 1120 : 255 - 0xff -- Background 0x46
      12'h461: dout <= 8'b00111000; // 1121 :  56 - 0x38
      12'h462: dout <= 8'b01101100; // 1122 : 108 - 0x6c
      12'h463: dout <= 8'b11000110; // 1123 : 198 - 0xc6
      12'h464: dout <= 8'b10000011; // 1124 : 131 - 0x83
      12'h465: dout <= 8'b11111111; // 1125 : 255 - 0xff
      12'h466: dout <= 8'b11111111; // 1126 : 255 - 0xff
      12'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0 -- plane 1
      12'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      12'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b10000001; // 1135 : 129 - 0x81
      12'h470: dout <= 8'b00111000; // 1136 :  56 - 0x38 -- Background 0x47
      12'h471: dout <= 8'b01101100; // 1137 : 108 - 0x6c
      12'h472: dout <= 8'b11000110; // 1138 : 198 - 0xc6
      12'h473: dout <= 8'b10000011; // 1139 : 131 - 0x83
      12'h474: dout <= 8'b11111111; // 1140 : 255 - 0xff
      12'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      12'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0 -- plane 1
      12'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      12'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b10000001; // 1150 : 129 - 0x81
      12'h47F: dout <= 8'b10000001; // 1151 : 129 - 0x81
      12'h480: dout <= 8'b01101100; // 1152 : 108 - 0x6c -- Background 0x48
      12'h481: dout <= 8'b11000110; // 1153 : 198 - 0xc6
      12'h482: dout <= 8'b10000011; // 1154 : 131 - 0x83
      12'h483: dout <= 8'b11111111; // 1155 : 255 - 0xff
      12'h484: dout <= 8'b11111111; // 1156 : 255 - 0xff
      12'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout <= 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout <= 8'b10000001; // 1166 : 129 - 0x81
      12'h48F: dout <= 8'b10000001; // 1167 : 129 - 0x81
      12'h490: dout <= 8'b11000110; // 1168 : 198 - 0xc6 -- Background 0x49
      12'h491: dout <= 8'b10000011; // 1169 : 131 - 0x83
      12'h492: dout <= 8'b11111111; // 1170 : 255 - 0xff
      12'h493: dout <= 8'b11111111; // 1171 : 255 - 0xff
      12'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b10000001; // 1180 : 129 - 0x81
      12'h49D: dout <= 8'b11111111; // 1181 : 255 - 0xff
      12'h49E: dout <= 8'b10000001; // 1182 : 129 - 0x81
      12'h49F: dout <= 8'b10000001; // 1183 : 129 - 0x81
      12'h4A0: dout <= 8'b10000011; // 1184 : 131 - 0x83 -- Background 0x4a
      12'h4A1: dout <= 8'b11111111; // 1185 : 255 - 0xff
      12'h4A2: dout <= 8'b11111111; // 1186 : 255 - 0xff
      12'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout <= 8'b00000000; // 1188 :   0 - 0x0
      12'h4A5: dout <= 8'b00000000; // 1189 :   0 - 0x0
      12'h4A6: dout <= 8'b00000000; // 1190 :   0 - 0x0
      12'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout <= 8'b10000001; // 1195 : 129 - 0x81
      12'h4AC: dout <= 8'b10000001; // 1196 : 129 - 0x81
      12'h4AD: dout <= 8'b11111111; // 1197 : 255 - 0xff
      12'h4AE: dout <= 8'b10000001; // 1198 : 129 - 0x81
      12'h4AF: dout <= 8'b10000001; // 1199 : 129 - 0x81
      12'h4B0: dout <= 8'b11111111; // 1200 : 255 - 0xff -- Background 0x4b
      12'h4B1: dout <= 8'b11111111; // 1201 : 255 - 0xff
      12'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout <= 8'b00000000; // 1204 :   0 - 0x0
      12'h4B5: dout <= 8'b00000000; // 1205 :   0 - 0x0
      12'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      12'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout <= 8'b10000001; // 1210 : 129 - 0x81
      12'h4BB: dout <= 8'b10000001; // 1211 : 129 - 0x81
      12'h4BC: dout <= 8'b10000001; // 1212 : 129 - 0x81
      12'h4BD: dout <= 8'b11111111; // 1213 : 255 - 0xff
      12'h4BE: dout <= 8'b10000001; // 1214 : 129 - 0x81
      12'h4BF: dout <= 8'b10000001; // 1215 : 129 - 0x81
      12'h4C0: dout <= 8'b10111111; // 1216 : 191 - 0xbf -- Background 0x4c
      12'h4C1: dout <= 8'b01011111; // 1217 :  95 - 0x5f
      12'h4C2: dout <= 8'b01011111; // 1218 :  95 - 0x5f
      12'h4C3: dout <= 8'b01011111; // 1219 :  95 - 0x5f
      12'h4C4: dout <= 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout <= 8'b01011111; // 1221 :  95 - 0x5f
      12'h4C6: dout <= 8'b01010001; // 1222 :  81 - 0x51
      12'h4C7: dout <= 8'b01010101; // 1223 :  85 - 0x55
      12'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- plane 1
      12'h4C9: dout <= 8'b01111111; // 1225 : 127 - 0x7f
      12'h4CA: dout <= 8'b01111111; // 1226 : 127 - 0x7f
      12'h4CB: dout <= 8'b01111111; // 1227 : 127 - 0x7f
      12'h4CC: dout <= 8'b01111111; // 1228 : 127 - 0x7f
      12'h4CD: dout <= 8'b01111111; // 1229 : 127 - 0x7f
      12'h4CE: dout <= 8'b01111111; // 1230 : 127 - 0x7f
      12'h4CF: dout <= 8'b01111111; // 1231 : 127 - 0x7f
      12'h4D0: dout <= 8'b01010001; // 1232 :  81 - 0x51 -- Background 0x4d
      12'h4D1: dout <= 8'b01011111; // 1233 :  95 - 0x5f
      12'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout <= 8'b01011111; // 1235 :  95 - 0x5f
      12'h4D4: dout <= 8'b01011111; // 1236 :  95 - 0x5f
      12'h4D5: dout <= 8'b01011111; // 1237 :  95 - 0x5f
      12'h4D6: dout <= 8'b01011111; // 1238 :  95 - 0x5f
      12'h4D7: dout <= 8'b10111111; // 1239 : 191 - 0xbf
      12'h4D8: dout <= 8'b01111111; // 1240 : 127 - 0x7f -- plane 1
      12'h4D9: dout <= 8'b01111111; // 1241 : 127 - 0x7f
      12'h4DA: dout <= 8'b01111111; // 1242 : 127 - 0x7f
      12'h4DB: dout <= 8'b01111111; // 1243 : 127 - 0x7f
      12'h4DC: dout <= 8'b01110010; // 1244 : 114 - 0x72
      12'h4DD: dout <= 8'b01111111; // 1245 : 127 - 0x7f
      12'h4DE: dout <= 8'b01111111; // 1246 : 127 - 0x7f
      12'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      12'h4E0: dout <= 8'b11111111; // 1248 : 255 - 0xff -- Background 0x4e
      12'h4E1: dout <= 8'b11111110; // 1249 : 254 - 0xfe
      12'h4E2: dout <= 8'b11111110; // 1250 : 254 - 0xfe
      12'h4E3: dout <= 8'b11111110; // 1251 : 254 - 0xfe
      12'h4E4: dout <= 8'b00000000; // 1252 :   0 - 0x0
      12'h4E5: dout <= 8'b11111110; // 1253 : 254 - 0xfe
      12'h4E6: dout <= 8'b00100110; // 1254 :  38 - 0x26
      12'h4E7: dout <= 8'b00100110; // 1255 :  38 - 0x26
      12'h4E8: dout <= 8'b11111111; // 1256 : 255 - 0xff -- plane 1
      12'h4E9: dout <= 8'b11111110; // 1257 : 254 - 0xfe
      12'h4EA: dout <= 8'b11111110; // 1258 : 254 - 0xfe
      12'h4EB: dout <= 8'b11111110; // 1259 : 254 - 0xfe
      12'h4EC: dout <= 8'b11111110; // 1260 : 254 - 0xfe
      12'h4ED: dout <= 8'b11111110; // 1261 : 254 - 0xfe
      12'h4EE: dout <= 8'b11111110; // 1262 : 254 - 0xfe
      12'h4EF: dout <= 8'b11111110; // 1263 : 254 - 0xfe
      12'h4F0: dout <= 8'b00100010; // 1264 :  34 - 0x22 -- Background 0x4f
      12'h4F1: dout <= 8'b11111110; // 1265 : 254 - 0xfe
      12'h4F2: dout <= 8'b00000000; // 1266 :   0 - 0x0
      12'h4F3: dout <= 8'b11111110; // 1267 : 254 - 0xfe
      12'h4F4: dout <= 8'b11111110; // 1268 : 254 - 0xfe
      12'h4F5: dout <= 8'b11111110; // 1269 : 254 - 0xfe
      12'h4F6: dout <= 8'b11111110; // 1270 : 254 - 0xfe
      12'h4F7: dout <= 8'b11111111; // 1271 : 255 - 0xff
      12'h4F8: dout <= 8'b11111110; // 1272 : 254 - 0xfe -- plane 1
      12'h4F9: dout <= 8'b11111110; // 1273 : 254 - 0xfe
      12'h4FA: dout <= 8'b11111110; // 1274 : 254 - 0xfe
      12'h4FB: dout <= 8'b11111110; // 1275 : 254 - 0xfe
      12'h4FC: dout <= 8'b01001010; // 1276 :  74 - 0x4a
      12'h4FD: dout <= 8'b11111110; // 1277 : 254 - 0xfe
      12'h4FE: dout <= 8'b11111110; // 1278 : 254 - 0xfe
      12'h4FF: dout <= 8'b11111111; // 1279 : 255 - 0xff
      12'h500: dout <= 8'b00000111; // 1280 :   7 - 0x7 -- Background 0x50
      12'h501: dout <= 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout <= 8'b00001111; // 1282 :  15 - 0xf
      12'h503: dout <= 8'b00011111; // 1283 :  31 - 0x1f
      12'h504: dout <= 8'b00011111; // 1284 :  31 - 0x1f
      12'h505: dout <= 8'b00011111; // 1285 :  31 - 0x1f
      12'h506: dout <= 8'b00011111; // 1286 :  31 - 0x1f
      12'h507: dout <= 8'b00011111; // 1287 :  31 - 0x1f
      12'h508: dout <= 8'b00000101; // 1288 :   5 - 0x5 -- plane 1
      12'h509: dout <= 8'b00001111; // 1289 :  15 - 0xf
      12'h50A: dout <= 8'b00001011; // 1290 :  11 - 0xb
      12'h50B: dout <= 8'b00011011; // 1291 :  27 - 0x1b
      12'h50C: dout <= 8'b00010011; // 1292 :  19 - 0x13
      12'h50D: dout <= 8'b00010011; // 1293 :  19 - 0x13
      12'h50E: dout <= 8'b00010011; // 1294 :  19 - 0x13
      12'h50F: dout <= 8'b00010011; // 1295 :  19 - 0x13
      12'h510: dout <= 8'b00011111; // 1296 :  31 - 0x1f -- Background 0x51
      12'h511: dout <= 8'b00011111; // 1297 :  31 - 0x1f
      12'h512: dout <= 8'b00011111; // 1298 :  31 - 0x1f
      12'h513: dout <= 8'b00011111; // 1299 :  31 - 0x1f
      12'h514: dout <= 8'b00011111; // 1300 :  31 - 0x1f
      12'h515: dout <= 8'b00001111; // 1301 :  15 - 0xf
      12'h516: dout <= 8'b00000000; // 1302 :   0 - 0x0
      12'h517: dout <= 8'b00000111; // 1303 :   7 - 0x7
      12'h518: dout <= 8'b00010011; // 1304 :  19 - 0x13 -- plane 1
      12'h519: dout <= 8'b00010011; // 1305 :  19 - 0x13
      12'h51A: dout <= 8'b00010011; // 1306 :  19 - 0x13
      12'h51B: dout <= 8'b00010011; // 1307 :  19 - 0x13
      12'h51C: dout <= 8'b00011011; // 1308 :  27 - 0x1b
      12'h51D: dout <= 8'b00001011; // 1309 :  11 - 0xb
      12'h51E: dout <= 8'b00001111; // 1310 :  15 - 0xf
      12'h51F: dout <= 8'b00000101; // 1311 :   5 - 0x5
      12'h520: dout <= 8'b00000111; // 1312 :   7 - 0x7 -- Background 0x52
      12'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout <= 8'b00001111; // 1314 :  15 - 0xf
      12'h523: dout <= 8'b00011111; // 1315 :  31 - 0x1f
      12'h524: dout <= 8'b00011111; // 1316 :  31 - 0x1f
      12'h525: dout <= 8'b00011111; // 1317 :  31 - 0x1f
      12'h526: dout <= 8'b00011111; // 1318 :  31 - 0x1f
      12'h527: dout <= 8'b00011111; // 1319 :  31 - 0x1f
      12'h528: dout <= 8'b00000101; // 1320 :   5 - 0x5 -- plane 1
      12'h529: dout <= 8'b00001111; // 1321 :  15 - 0xf
      12'h52A: dout <= 8'b00001011; // 1322 :  11 - 0xb
      12'h52B: dout <= 8'b00011011; // 1323 :  27 - 0x1b
      12'h52C: dout <= 8'b00010011; // 1324 :  19 - 0x13
      12'h52D: dout <= 8'b00010011; // 1325 :  19 - 0x13
      12'h52E: dout <= 8'b00010011; // 1326 :  19 - 0x13
      12'h52F: dout <= 8'b00010011; // 1327 :  19 - 0x13
      12'h530: dout <= 8'b00011111; // 1328 :  31 - 0x1f -- Background 0x53
      12'h531: dout <= 8'b00011111; // 1329 :  31 - 0x1f
      12'h532: dout <= 8'b00011111; // 1330 :  31 - 0x1f
      12'h533: dout <= 8'b00011111; // 1331 :  31 - 0x1f
      12'h534: dout <= 8'b00011111; // 1332 :  31 - 0x1f
      12'h535: dout <= 8'b00001111; // 1333 :  15 - 0xf
      12'h536: dout <= 8'b00000000; // 1334 :   0 - 0x0
      12'h537: dout <= 8'b00000111; // 1335 :   7 - 0x7
      12'h538: dout <= 8'b00010011; // 1336 :  19 - 0x13 -- plane 1
      12'h539: dout <= 8'b00010011; // 1337 :  19 - 0x13
      12'h53A: dout <= 8'b00010011; // 1338 :  19 - 0x13
      12'h53B: dout <= 8'b00010011; // 1339 :  19 - 0x13
      12'h53C: dout <= 8'b00011011; // 1340 :  27 - 0x1b
      12'h53D: dout <= 8'b00001011; // 1341 :  11 - 0xb
      12'h53E: dout <= 8'b00001111; // 1342 :  15 - 0xf
      12'h53F: dout <= 8'b00000101; // 1343 :   5 - 0x5
      12'h540: dout <= 8'b11100000; // 1344 : 224 - 0xe0 -- Background 0x54
      12'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout <= 8'b11110001; // 1346 : 241 - 0xf1
      12'h543: dout <= 8'b11111011; // 1347 : 251 - 0xfb
      12'h544: dout <= 8'b11111011; // 1348 : 251 - 0xfb
      12'h545: dout <= 8'b11111011; // 1349 : 251 - 0xfb
      12'h546: dout <= 8'b11111011; // 1350 : 251 - 0xfb
      12'h547: dout <= 8'b11111011; // 1351 : 251 - 0xfb
      12'h548: dout <= 8'b10100000; // 1352 : 160 - 0xa0 -- plane 1
      12'h549: dout <= 8'b11110001; // 1353 : 241 - 0xf1
      12'h54A: dout <= 8'b11010001; // 1354 : 209 - 0xd1
      12'h54B: dout <= 8'b11011011; // 1355 : 219 - 0xdb
      12'h54C: dout <= 8'b11001010; // 1356 : 202 - 0xca
      12'h54D: dout <= 8'b11001010; // 1357 : 202 - 0xca
      12'h54E: dout <= 8'b11001010; // 1358 : 202 - 0xca
      12'h54F: dout <= 8'b11001010; // 1359 : 202 - 0xca
      12'h550: dout <= 8'b11111011; // 1360 : 251 - 0xfb -- Background 0x55
      12'h551: dout <= 8'b11111011; // 1361 : 251 - 0xfb
      12'h552: dout <= 8'b11111011; // 1362 : 251 - 0xfb
      12'h553: dout <= 8'b11111011; // 1363 : 251 - 0xfb
      12'h554: dout <= 8'b11111011; // 1364 : 251 - 0xfb
      12'h555: dout <= 8'b11110001; // 1365 : 241 - 0xf1
      12'h556: dout <= 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout <= 8'b11100000; // 1367 : 224 - 0xe0
      12'h558: dout <= 8'b11001010; // 1368 : 202 - 0xca -- plane 1
      12'h559: dout <= 8'b11001010; // 1369 : 202 - 0xca
      12'h55A: dout <= 8'b11001010; // 1370 : 202 - 0xca
      12'h55B: dout <= 8'b11001010; // 1371 : 202 - 0xca
      12'h55C: dout <= 8'b11011011; // 1372 : 219 - 0xdb
      12'h55D: dout <= 8'b11010001; // 1373 : 209 - 0xd1
      12'h55E: dout <= 8'b11110001; // 1374 : 241 - 0xf1
      12'h55F: dout <= 8'b10100000; // 1375 : 160 - 0xa0
      12'h560: dout <= 8'b11100000; // 1376 : 224 - 0xe0 -- Background 0x56
      12'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout <= 8'b11110001; // 1378 : 241 - 0xf1
      12'h563: dout <= 8'b11111011; // 1379 : 251 - 0xfb
      12'h564: dout <= 8'b11111011; // 1380 : 251 - 0xfb
      12'h565: dout <= 8'b11111011; // 1381 : 251 - 0xfb
      12'h566: dout <= 8'b11111011; // 1382 : 251 - 0xfb
      12'h567: dout <= 8'b11111011; // 1383 : 251 - 0xfb
      12'h568: dout <= 8'b10100000; // 1384 : 160 - 0xa0 -- plane 1
      12'h569: dout <= 8'b11110001; // 1385 : 241 - 0xf1
      12'h56A: dout <= 8'b11010001; // 1386 : 209 - 0xd1
      12'h56B: dout <= 8'b11011011; // 1387 : 219 - 0xdb
      12'h56C: dout <= 8'b11001010; // 1388 : 202 - 0xca
      12'h56D: dout <= 8'b11001010; // 1389 : 202 - 0xca
      12'h56E: dout <= 8'b11001010; // 1390 : 202 - 0xca
      12'h56F: dout <= 8'b11001010; // 1391 : 202 - 0xca
      12'h570: dout <= 8'b11111011; // 1392 : 251 - 0xfb -- Background 0x57
      12'h571: dout <= 8'b11111011; // 1393 : 251 - 0xfb
      12'h572: dout <= 8'b11111011; // 1394 : 251 - 0xfb
      12'h573: dout <= 8'b11111011; // 1395 : 251 - 0xfb
      12'h574: dout <= 8'b11111011; // 1396 : 251 - 0xfb
      12'h575: dout <= 8'b11110001; // 1397 : 241 - 0xf1
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b11100000; // 1399 : 224 - 0xe0
      12'h578: dout <= 8'b11001010; // 1400 : 202 - 0xca -- plane 1
      12'h579: dout <= 8'b11001010; // 1401 : 202 - 0xca
      12'h57A: dout <= 8'b11001010; // 1402 : 202 - 0xca
      12'h57B: dout <= 8'b11001010; // 1403 : 202 - 0xca
      12'h57C: dout <= 8'b11011011; // 1404 : 219 - 0xdb
      12'h57D: dout <= 8'b11010001; // 1405 : 209 - 0xd1
      12'h57E: dout <= 8'b11110000; // 1406 : 240 - 0xf0
      12'h57F: dout <= 8'b10100000; // 1407 : 160 - 0xa0
      12'h580: dout <= 8'b11111100; // 1408 : 252 - 0xfc -- Background 0x58
      12'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout <= 8'b11111110; // 1410 : 254 - 0xfe
      12'h583: dout <= 8'b11111111; // 1411 : 255 - 0xff
      12'h584: dout <= 8'b11111111; // 1412 : 255 - 0xff
      12'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout <= 8'b11111111; // 1414 : 255 - 0xff
      12'h587: dout <= 8'b11111111; // 1415 : 255 - 0xff
      12'h588: dout <= 8'b10110100; // 1416 : 180 - 0xb4 -- plane 1
      12'h589: dout <= 8'b11111110; // 1417 : 254 - 0xfe
      12'h58A: dout <= 8'b01111010; // 1418 : 122 - 0x7a
      12'h58B: dout <= 8'b01111011; // 1419 : 123 - 0x7b
      12'h58C: dout <= 8'b01111001; // 1420 : 121 - 0x79
      12'h58D: dout <= 8'b01111001; // 1421 : 121 - 0x79
      12'h58E: dout <= 8'b01111001; // 1422 : 121 - 0x79
      12'h58F: dout <= 8'b01111001; // 1423 : 121 - 0x79
      12'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Background 0x59
      12'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      12'h592: dout <= 8'b11111111; // 1426 : 255 - 0xff
      12'h593: dout <= 8'b11111111; // 1427 : 255 - 0xff
      12'h594: dout <= 8'b11111111; // 1428 : 255 - 0xff
      12'h595: dout <= 8'b11111110; // 1429 : 254 - 0xfe
      12'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout <= 8'b11111100; // 1431 : 252 - 0xfc
      12'h598: dout <= 8'b01111001; // 1432 : 121 - 0x79 -- plane 1
      12'h599: dout <= 8'b01111001; // 1433 : 121 - 0x79
      12'h59A: dout <= 8'b01111001; // 1434 : 121 - 0x79
      12'h59B: dout <= 8'b01111001; // 1435 : 121 - 0x79
      12'h59C: dout <= 8'b01111011; // 1436 : 123 - 0x7b
      12'h59D: dout <= 8'b01111010; // 1437 : 122 - 0x7a
      12'h59E: dout <= 8'b11111110; // 1438 : 254 - 0xfe
      12'h59F: dout <= 8'b10110100; // 1439 : 180 - 0xb4
      12'h5A0: dout <= 8'b11111100; // 1440 : 252 - 0xfc -- Background 0x5a
      12'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout <= 8'b11111110; // 1442 : 254 - 0xfe
      12'h5A3: dout <= 8'b11111111; // 1443 : 255 - 0xff
      12'h5A4: dout <= 8'b11111111; // 1444 : 255 - 0xff
      12'h5A5: dout <= 8'b11111111; // 1445 : 255 - 0xff
      12'h5A6: dout <= 8'b11111111; // 1446 : 255 - 0xff
      12'h5A7: dout <= 8'b11111111; // 1447 : 255 - 0xff
      12'h5A8: dout <= 8'b10110100; // 1448 : 180 - 0xb4 -- plane 1
      12'h5A9: dout <= 8'b11111110; // 1449 : 254 - 0xfe
      12'h5AA: dout <= 8'b01111010; // 1450 : 122 - 0x7a
      12'h5AB: dout <= 8'b01111011; // 1451 : 123 - 0x7b
      12'h5AC: dout <= 8'b01111001; // 1452 : 121 - 0x79
      12'h5AD: dout <= 8'b01111001; // 1453 : 121 - 0x79
      12'h5AE: dout <= 8'b01111001; // 1454 : 121 - 0x79
      12'h5AF: dout <= 8'b01111001; // 1455 : 121 - 0x79
      12'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Background 0x5b
      12'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      12'h5B2: dout <= 8'b11111111; // 1458 : 255 - 0xff
      12'h5B3: dout <= 8'b11111111; // 1459 : 255 - 0xff
      12'h5B4: dout <= 8'b11111111; // 1460 : 255 - 0xff
      12'h5B5: dout <= 8'b11111110; // 1461 : 254 - 0xfe
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b11111100; // 1463 : 252 - 0xfc
      12'h5B8: dout <= 8'b01111001; // 1464 : 121 - 0x79 -- plane 1
      12'h5B9: dout <= 8'b01111001; // 1465 : 121 - 0x79
      12'h5BA: dout <= 8'b01111001; // 1466 : 121 - 0x79
      12'h5BB: dout <= 8'b01111001; // 1467 : 121 - 0x79
      12'h5BC: dout <= 8'b01111011; // 1468 : 123 - 0x7b
      12'h5BD: dout <= 8'b01111010; // 1469 : 122 - 0x7a
      12'h5BE: dout <= 8'b11111110; // 1470 : 254 - 0xfe
      12'h5BF: dout <= 8'b10110100; // 1471 : 180 - 0xb4
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Background 0x5c
      12'h5C1: dout <= 8'b00000000; // 1473 :   0 - 0x0
      12'h5C2: dout <= 8'b00011111; // 1474 :  31 - 0x1f
      12'h5C3: dout <= 8'b00010000; // 1475 :  16 - 0x10
      12'h5C4: dout <= 8'b00010000; // 1476 :  16 - 0x10
      12'h5C5: dout <= 8'b00011111; // 1477 :  31 - 0x1f
      12'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b01111111; // 1480 : 127 - 0x7f -- plane 1
      12'h5C9: dout <= 8'b10111111; // 1481 : 191 - 0xbf
      12'h5CA: dout <= 8'b11111111; // 1482 : 255 - 0xff
      12'h5CB: dout <= 8'b10110010; // 1483 : 178 - 0xb2
      12'h5CC: dout <= 8'b10110001; // 1484 : 177 - 0xb1
      12'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      12'h5CE: dout <= 8'b10111111; // 1486 : 191 - 0xbf
      12'h5CF: dout <= 8'b01111111; // 1487 : 127 - 0x7f
      12'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Background 0x5d
      12'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout <= 8'b11111000; // 1490 : 248 - 0xf8
      12'h5D3: dout <= 8'b00001000; // 1491 :   8 - 0x8
      12'h5D4: dout <= 8'b00001000; // 1492 :   8 - 0x8
      12'h5D5: dout <= 8'b11111000; // 1493 : 248 - 0xf8
      12'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b11111110; // 1496 : 254 - 0xfe -- plane 1
      12'h5D9: dout <= 8'b11111101; // 1497 : 253 - 0xfd
      12'h5DA: dout <= 8'b11111111; // 1498 : 255 - 0xff
      12'h5DB: dout <= 8'b11001101; // 1499 : 205 - 0xcd
      12'h5DC: dout <= 8'b01101101; // 1500 : 109 - 0x6d
      12'h5DD: dout <= 8'b11111111; // 1501 : 255 - 0xff
      12'h5DE: dout <= 8'b11111101; // 1502 : 253 - 0xfd
      12'h5DF: dout <= 8'b11111110; // 1503 : 254 - 0xfe
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Background 0x5e
      12'h5E1: dout <= 8'b00000001; // 1505 :   1 - 0x1
      12'h5E2: dout <= 8'b00000010; // 1506 :   2 - 0x2
      12'h5E3: dout <= 8'b00000010; // 1507 :   2 - 0x2
      12'h5E4: dout <= 8'b11110001; // 1508 : 241 - 0xf1
      12'h5E5: dout <= 8'b00001000; // 1509 :   8 - 0x8
      12'h5E6: dout <= 8'b00000100; // 1510 :   4 - 0x4
      12'h5E7: dout <= 8'b00000011; // 1511 :   3 - 0x3
      12'h5E8: dout <= 8'b11111111; // 1512 : 255 - 0xff -- plane 1
      12'h5E9: dout <= 8'b11111111; // 1513 : 255 - 0xff
      12'h5EA: dout <= 8'b10101110; // 1514 : 174 - 0xae
      12'h5EB: dout <= 8'b11111110; // 1515 : 254 - 0xfe
      12'h5EC: dout <= 8'b11111111; // 1516 : 255 - 0xff
      12'h5ED: dout <= 8'b00001111; // 1517 :  15 - 0xf
      12'h5EE: dout <= 8'b00000111; // 1518 :   7 - 0x7
      12'h5EF: dout <= 8'b00000011; // 1519 :   3 - 0x3
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Background 0x5f
      12'h5F1: dout <= 8'b10000000; // 1521 : 128 - 0x80
      12'h5F2: dout <= 8'b01000000; // 1522 :  64 - 0x40
      12'h5F3: dout <= 8'b01000000; // 1523 :  64 - 0x40
      12'h5F4: dout <= 8'b10001111; // 1524 : 143 - 0x8f
      12'h5F5: dout <= 8'b00010000; // 1525 :  16 - 0x10
      12'h5F6: dout <= 8'b00100000; // 1526 :  32 - 0x20
      12'h5F7: dout <= 8'b11000000; // 1527 : 192 - 0xc0
      12'h5F8: dout <= 8'b11111111; // 1528 : 255 - 0xff -- plane 1
      12'h5F9: dout <= 8'b11111111; // 1529 : 255 - 0xff
      12'h5FA: dout <= 8'b01110101; // 1530 : 117 - 0x75
      12'h5FB: dout <= 8'b01111111; // 1531 : 127 - 0x7f
      12'h5FC: dout <= 8'b11111111; // 1532 : 255 - 0xff
      12'h5FD: dout <= 8'b11110000; // 1533 : 240 - 0xf0
      12'h5FE: dout <= 8'b11100000; // 1534 : 224 - 0xe0
      12'h5FF: dout <= 8'b11000000; // 1535 : 192 - 0xc0
      12'h600: dout <= 8'b00000011; // 1536 :   3 - 0x3 -- Background 0x60
      12'h601: dout <= 8'b00000100; // 1537 :   4 - 0x4
      12'h602: dout <= 8'b00001000; // 1538 :   8 - 0x8
      12'h603: dout <= 8'b11110001; // 1539 : 241 - 0xf1
      12'h604: dout <= 8'b00000010; // 1540 :   2 - 0x2
      12'h605: dout <= 8'b00000010; // 1541 :   2 - 0x2
      12'h606: dout <= 8'b00000001; // 1542 :   1 - 0x1
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00000011; // 1544 :   3 - 0x3 -- plane 1
      12'h609: dout <= 8'b00000111; // 1545 :   7 - 0x7
      12'h60A: dout <= 8'b00001111; // 1546 :  15 - 0xf
      12'h60B: dout <= 8'b11111111; // 1547 : 255 - 0xff
      12'h60C: dout <= 8'b11111110; // 1548 : 254 - 0xfe
      12'h60D: dout <= 8'b10101110; // 1549 : 174 - 0xae
      12'h60E: dout <= 8'b11111111; // 1550 : 255 - 0xff
      12'h60F: dout <= 8'b11111111; // 1551 : 255 - 0xff
      12'h610: dout <= 8'b11000000; // 1552 : 192 - 0xc0 -- Background 0x61
      12'h611: dout <= 8'b00100000; // 1553 :  32 - 0x20
      12'h612: dout <= 8'b00010000; // 1554 :  16 - 0x10
      12'h613: dout <= 8'b10001111; // 1555 : 143 - 0x8f
      12'h614: dout <= 8'b01000000; // 1556 :  64 - 0x40
      12'h615: dout <= 8'b01000000; // 1557 :  64 - 0x40
      12'h616: dout <= 8'b10000000; // 1558 : 128 - 0x80
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b11000000; // 1560 : 192 - 0xc0 -- plane 1
      12'h619: dout <= 8'b11100000; // 1561 : 224 - 0xe0
      12'h61A: dout <= 8'b11110000; // 1562 : 240 - 0xf0
      12'h61B: dout <= 8'b11111111; // 1563 : 255 - 0xff
      12'h61C: dout <= 8'b01111111; // 1564 : 127 - 0x7f
      12'h61D: dout <= 8'b01110101; // 1565 : 117 - 0x75
      12'h61E: dout <= 8'b11111111; // 1566 : 255 - 0xff
      12'h61F: dout <= 8'b11111111; // 1567 : 255 - 0xff
      12'h620: dout <= 8'b11111111; // 1568 : 255 - 0xff -- Background 0x62
      12'h621: dout <= 8'b11111111; // 1569 : 255 - 0xff
      12'h622: dout <= 8'b11000011; // 1570 : 195 - 0xc3
      12'h623: dout <= 8'b10000001; // 1571 : 129 - 0x81
      12'h624: dout <= 8'b10000001; // 1572 : 129 - 0x81
      12'h625: dout <= 8'b11000011; // 1573 : 195 - 0xc3
      12'h626: dout <= 8'b11111111; // 1574 : 255 - 0xff
      12'h627: dout <= 8'b11111111; // 1575 : 255 - 0xff
      12'h628: dout <= 8'b11111111; // 1576 : 255 - 0xff -- plane 1
      12'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout <= 8'b11000011; // 1578 : 195 - 0xc3
      12'h62B: dout <= 8'b10000001; // 1579 : 129 - 0x81
      12'h62C: dout <= 8'b10000001; // 1580 : 129 - 0x81
      12'h62D: dout <= 8'b11000011; // 1581 : 195 - 0xc3
      12'h62E: dout <= 8'b11111111; // 1582 : 255 - 0xff
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b11111111; // 1584 : 255 - 0xff -- Background 0x63
      12'h631: dout <= 8'b10011001; // 1585 : 153 - 0x99
      12'h632: dout <= 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout <= 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout <= 8'b10000001; // 1589 : 129 - 0x81
      12'h636: dout <= 8'b10000001; // 1590 : 129 - 0x81
      12'h637: dout <= 8'b10000001; // 1591 : 129 - 0x81
      12'h638: dout <= 8'b10000001; // 1592 : 129 - 0x81 -- plane 1
      12'h639: dout <= 8'b01100110; // 1593 : 102 - 0x66
      12'h63A: dout <= 8'b01111110; // 1594 : 126 - 0x7e
      12'h63B: dout <= 8'b01111110; // 1595 : 126 - 0x7e
      12'h63C: dout <= 8'b01111110; // 1596 : 126 - 0x7e
      12'h63D: dout <= 8'b11111111; // 1597 : 255 - 0xff
      12'h63E: dout <= 8'b11111111; // 1598 : 255 - 0xff
      12'h63F: dout <= 8'b01111110; // 1599 : 126 - 0x7e
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Background 0x64
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b01100000; // 1604 :  96 - 0x60
      12'h645: dout <= 8'b01100000; // 1605 :  96 - 0x60
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Background 0x65
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout <= 8'b01101100; // 1620 : 108 - 0x6c
      12'h655: dout <= 8'b01101100; // 1621 : 108 - 0x6c
      12'h656: dout <= 8'b00001000; // 1622 :   8 - 0x8
      12'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00111100; // 1632 :  60 - 0x3c -- Background 0x66
      12'h661: dout <= 8'b00011000; // 1633 :  24 - 0x18
      12'h662: dout <= 8'b00011000; // 1634 :  24 - 0x18
      12'h663: dout <= 8'b00011000; // 1635 :  24 - 0x18
      12'h664: dout <= 8'b00011000; // 1636 :  24 - 0x18
      12'h665: dout <= 8'b00011000; // 1637 :  24 - 0x18
      12'h666: dout <= 8'b00111100; // 1638 :  60 - 0x3c
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b11111111; // 1648 : 255 - 0xff -- Background 0x67
      12'h671: dout <= 8'b01100110; // 1649 : 102 - 0x66
      12'h672: dout <= 8'b01100110; // 1650 : 102 - 0x66
      12'h673: dout <= 8'b01100110; // 1651 : 102 - 0x66
      12'h674: dout <= 8'b01100110; // 1652 : 102 - 0x66
      12'h675: dout <= 8'b01100110; // 1653 : 102 - 0x66
      12'h676: dout <= 8'b01100110; // 1654 : 102 - 0x66
      12'h677: dout <= 8'b11111111; // 1655 : 255 - 0xff
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b00000011; // 1664 :   3 - 0x3 -- Background 0x68
      12'h681: dout <= 8'b00000001; // 1665 :   1 - 0x1
      12'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000011; // 1672 :   3 - 0x3 -- plane 1
      12'h689: dout <= 8'b00000001; // 1673 :   1 - 0x1
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b10000011; // 1680 : 131 - 0x83 -- Background 0x69
      12'h691: dout <= 8'b11010001; // 1681 : 209 - 0xd1
      12'h692: dout <= 8'b11100001; // 1682 : 225 - 0xe1
      12'h693: dout <= 8'b11010001; // 1683 : 209 - 0xd1
      12'h694: dout <= 8'b00000010; // 1684 :   2 - 0x2
      12'h695: dout <= 8'b10000100; // 1685 : 132 - 0x84
      12'h696: dout <= 8'b11110000; // 1686 : 240 - 0xf0
      12'h697: dout <= 8'b11001110; // 1687 : 206 - 0xce
      12'h698: dout <= 8'b11111111; // 1688 : 255 - 0xff -- plane 1
      12'h699: dout <= 8'b11111111; // 1689 : 255 - 0xff
      12'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      12'h69B: dout <= 8'b11111111; // 1691 : 255 - 0xff
      12'h69C: dout <= 8'b11111111; // 1692 : 255 - 0xff
      12'h69D: dout <= 8'b11111111; // 1693 : 255 - 0xff
      12'h69E: dout <= 8'b11111111; // 1694 : 255 - 0xff
      12'h69F: dout <= 8'b11111111; // 1695 : 255 - 0xff
      12'h6A0: dout <= 8'b11000000; // 1696 : 192 - 0xc0 -- Background 0x6a
      12'h6A1: dout <= 8'b10000000; // 1697 : 128 - 0x80
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b11000000; // 1704 : 192 - 0xc0 -- plane 1
      12'h6A9: dout <= 8'b10000000; // 1705 : 128 - 0x80
      12'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b11000001; // 1712 : 193 - 0xc1 -- Background 0x6b
      12'h6B1: dout <= 8'b10001011; // 1713 : 139 - 0x8b
      12'h6B2: dout <= 8'b10000111; // 1714 : 135 - 0x87
      12'h6B3: dout <= 8'b10001011; // 1715 : 139 - 0x8b
      12'h6B4: dout <= 8'b01000000; // 1716 :  64 - 0x40
      12'h6B5: dout <= 8'b00100001; // 1717 :  33 - 0x21
      12'h6B6: dout <= 8'b00001111; // 1718 :  15 - 0xf
      12'h6B7: dout <= 8'b11010011; // 1719 : 211 - 0xd3
      12'h6B8: dout <= 8'b11111111; // 1720 : 255 - 0xff -- plane 1
      12'h6B9: dout <= 8'b11111111; // 1721 : 255 - 0xff
      12'h6BA: dout <= 8'b11111111; // 1722 : 255 - 0xff
      12'h6BB: dout <= 8'b11111111; // 1723 : 255 - 0xff
      12'h6BC: dout <= 8'b11111111; // 1724 : 255 - 0xff
      12'h6BD: dout <= 8'b11111111; // 1725 : 255 - 0xff
      12'h6BE: dout <= 8'b11111111; // 1726 : 255 - 0xff
      12'h6BF: dout <= 8'b11111111; // 1727 : 255 - 0xff
      12'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Background 0x6c
      12'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      12'h6C3: dout <= 8'b00011111; // 1731 :  31 - 0x1f
      12'h6C4: dout <= 8'b00001111; // 1732 :  15 - 0xf
      12'h6C5: dout <= 8'b00011110; // 1733 :  30 - 0x1e
      12'h6C6: dout <= 8'b00111111; // 1734 :  63 - 0x3f
      12'h6C7: dout <= 8'b01111111; // 1735 : 127 - 0x7f
      12'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff -- plane 1
      12'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      12'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      12'h6CB: dout <= 8'b00011111; // 1739 :  31 - 0x1f
      12'h6CC: dout <= 8'b00011111; // 1740 :  31 - 0x1f
      12'h6CD: dout <= 8'b00111111; // 1741 :  63 - 0x3f
      12'h6CE: dout <= 8'b01111111; // 1742 : 127 - 0x7f
      12'h6CF: dout <= 8'b11111111; // 1743 : 255 - 0xff
      12'h6D0: dout <= 8'b11111111; // 1744 : 255 - 0xff -- Background 0x6d
      12'h6D1: dout <= 8'b11111111; // 1745 : 255 - 0xff
      12'h6D2: dout <= 8'b11111111; // 1746 : 255 - 0xff
      12'h6D3: dout <= 8'b11111000; // 1747 : 248 - 0xf8
      12'h6D4: dout <= 8'b11110000; // 1748 : 240 - 0xf0
      12'h6D5: dout <= 8'b01111000; // 1749 : 120 - 0x78
      12'h6D6: dout <= 8'b11111100; // 1750 : 252 - 0xfc
      12'h6D7: dout <= 8'b11111110; // 1751 : 254 - 0xfe
      12'h6D8: dout <= 8'b11111111; // 1752 : 255 - 0xff -- plane 1
      12'h6D9: dout <= 8'b11111111; // 1753 : 255 - 0xff
      12'h6DA: dout <= 8'b11111111; // 1754 : 255 - 0xff
      12'h6DB: dout <= 8'b11111000; // 1755 : 248 - 0xf8
      12'h6DC: dout <= 8'b11111000; // 1756 : 248 - 0xf8
      12'h6DD: dout <= 8'b11111100; // 1757 : 252 - 0xfc
      12'h6DE: dout <= 8'b11111110; // 1758 : 254 - 0xfe
      12'h6DF: dout <= 8'b11111111; // 1759 : 255 - 0xff
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Background 0x6e
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b00111100; // 1765 :  60 - 0x3c
      12'h6E6: dout <= 8'b01000010; // 1766 :  66 - 0x42
      12'h6E7: dout <= 8'b10000001; // 1767 : 129 - 0x81
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b00111100; // 1773 :  60 - 0x3c
      12'h6EE: dout <= 8'b01000010; // 1774 :  66 - 0x42
      12'h6EF: dout <= 8'b10000001; // 1775 : 129 - 0x81
      12'h6F0: dout <= 8'b10000001; // 1776 : 129 - 0x81 -- Background 0x6f
      12'h6F1: dout <= 8'b10111101; // 1777 : 189 - 0xbd
      12'h6F2: dout <= 8'b01111110; // 1778 : 126 - 0x7e
      12'h6F3: dout <= 8'b11111111; // 1779 : 255 - 0xff
      12'h6F4: dout <= 8'b11100111; // 1780 : 231 - 0xe7
      12'h6F5: dout <= 8'b11111111; // 1781 : 255 - 0xff
      12'h6F6: dout <= 8'b11111111; // 1782 : 255 - 0xff
      12'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      12'h6F8: dout <= 8'b10000001; // 1784 : 129 - 0x81 -- plane 1
      12'h6F9: dout <= 8'b10111101; // 1785 : 189 - 0xbd
      12'h6FA: dout <= 8'b01111110; // 1786 : 126 - 0x7e
      12'h6FB: dout <= 8'b10100101; // 1787 : 165 - 0xa5
      12'h6FC: dout <= 8'b11011011; // 1788 : 219 - 0xdb
      12'h6FD: dout <= 8'b11100111; // 1789 : 231 - 0xe7
      12'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      12'h6FF: dout <= 8'b11111111; // 1791 : 255 - 0xff
      12'h700: dout <= 8'b00000001; // 1792 :   1 - 0x1 -- Background 0x70
      12'h701: dout <= 8'b00000111; // 1793 :   7 - 0x7
      12'h702: dout <= 8'b00011111; // 1794 :  31 - 0x1f
      12'h703: dout <= 8'b00111111; // 1795 :  63 - 0x3f
      12'h704: dout <= 8'b01111111; // 1796 : 127 - 0x7f
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout <= 8'b11011101; // 1799 : 221 - 0xdd
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout <= 8'b00000101; // 1801 :   5 - 0x5
      12'h70A: dout <= 8'b00011001; // 1802 :  25 - 0x19
      12'h70B: dout <= 8'b00110011; // 1803 :  51 - 0x33
      12'h70C: dout <= 8'b01100011; // 1804 :  99 - 0x63
      12'h70D: dout <= 8'b11000111; // 1805 : 199 - 0xc7
      12'h70E: dout <= 8'b11000111; // 1806 : 199 - 0xc7
      12'h70F: dout <= 8'b11000100; // 1807 : 196 - 0xc4
      12'h710: dout <= 8'b10001001; // 1808 : 137 - 0x89 -- Background 0x71
      12'h711: dout <= 8'b00000001; // 1809 :   1 - 0x1
      12'h712: dout <= 8'b00000001; // 1810 :   1 - 0x1
      12'h713: dout <= 8'b00000001; // 1811 :   1 - 0x1
      12'h714: dout <= 8'b00000001; // 1812 :   1 - 0x1
      12'h715: dout <= 8'b00000001; // 1813 :   1 - 0x1
      12'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout <= 8'b10000000; // 1816 : 128 - 0x80 -- plane 1
      12'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout <= 8'b00000001; // 1819 :   1 - 0x1
      12'h71C: dout <= 8'b00000001; // 1820 :   1 - 0x1
      12'h71D: dout <= 8'b00000001; // 1821 :   1 - 0x1
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b10000000; // 1824 : 128 - 0x80 -- Background 0x72
      12'h721: dout <= 8'b11100000; // 1825 : 224 - 0xe0
      12'h722: dout <= 8'b11111000; // 1826 : 248 - 0xf8
      12'h723: dout <= 8'b11111100; // 1827 : 252 - 0xfc
      12'h724: dout <= 8'b11111110; // 1828 : 254 - 0xfe
      12'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout <= 8'b00111011; // 1831 :  59 - 0x3b
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout <= 8'b10100000; // 1833 : 160 - 0xa0
      12'h72A: dout <= 8'b10011000; // 1834 : 152 - 0x98
      12'h72B: dout <= 8'b11001100; // 1835 : 204 - 0xcc
      12'h72C: dout <= 8'b11000110; // 1836 : 198 - 0xc6
      12'h72D: dout <= 8'b11100011; // 1837 : 227 - 0xe3
      12'h72E: dout <= 8'b11100011; // 1838 : 227 - 0xe3
      12'h72F: dout <= 8'b00100011; // 1839 :  35 - 0x23
      12'h730: dout <= 8'b00010001; // 1840 :  17 - 0x11 -- Background 0x73
      12'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout <= 8'b01000000; // 1845 :  64 - 0x40
      12'h736: dout <= 8'b10000000; // 1846 : 128 - 0x80
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00000001; // 1848 :   1 - 0x1 -- plane 1
      12'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b01000000; // 1853 :  64 - 0x40
      12'h73E: dout <= 8'b10000000; // 1854 : 128 - 0x80
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000001; // 1856 :   1 - 0x1 -- Background 0x74
      12'h741: dout <= 8'b00000001; // 1857 :   1 - 0x1
      12'h742: dout <= 8'b00000001; // 1858 :   1 - 0x1
      12'h743: dout <= 8'b00000001; // 1859 :   1 - 0x1
      12'h744: dout <= 8'b00000001; // 1860 :   1 - 0x1
      12'h745: dout <= 8'b00000001; // 1861 :   1 - 0x1
      12'h746: dout <= 8'b00000001; // 1862 :   1 - 0x1
      12'h747: dout <= 8'b00000001; // 1863 :   1 - 0x1
      12'h748: dout <= 8'b00000001; // 1864 :   1 - 0x1 -- plane 1
      12'h749: dout <= 8'b00000001; // 1865 :   1 - 0x1
      12'h74A: dout <= 8'b00000001; // 1866 :   1 - 0x1
      12'h74B: dout <= 8'b00000001; // 1867 :   1 - 0x1
      12'h74C: dout <= 8'b00000001; // 1868 :   1 - 0x1
      12'h74D: dout <= 8'b00000001; // 1869 :   1 - 0x1
      12'h74E: dout <= 8'b00000001; // 1870 :   1 - 0x1
      12'h74F: dout <= 8'b00000001; // 1871 :   1 - 0x1
      12'h750: dout <= 8'b10000000; // 1872 : 128 - 0x80 -- Background 0x75
      12'h751: dout <= 8'b10000000; // 1873 : 128 - 0x80
      12'h752: dout <= 8'b10000000; // 1874 : 128 - 0x80
      12'h753: dout <= 8'b10000000; // 1875 : 128 - 0x80
      12'h754: dout <= 8'b10000000; // 1876 : 128 - 0x80
      12'h755: dout <= 8'b10000000; // 1877 : 128 - 0x80
      12'h756: dout <= 8'b10000000; // 1878 : 128 - 0x80
      12'h757: dout <= 8'b10000000; // 1879 : 128 - 0x80
      12'h758: dout <= 8'b10000000; // 1880 : 128 - 0x80 -- plane 1
      12'h759: dout <= 8'b10000000; // 1881 : 128 - 0x80
      12'h75A: dout <= 8'b10000000; // 1882 : 128 - 0x80
      12'h75B: dout <= 8'b10000000; // 1883 : 128 - 0x80
      12'h75C: dout <= 8'b10000000; // 1884 : 128 - 0x80
      12'h75D: dout <= 8'b10000000; // 1885 : 128 - 0x80
      12'h75E: dout <= 8'b10000000; // 1886 : 128 - 0x80
      12'h75F: dout <= 8'b10000000; // 1887 : 128 - 0x80
      12'h760: dout <= 8'b00000001; // 1888 :   1 - 0x1 -- Background 0x76
      12'h761: dout <= 8'b00000011; // 1889 :   3 - 0x3
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000011; // 1892 :   3 - 0x3
      12'h765: dout <= 8'b00011001; // 1893 :  25 - 0x19
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00000001; // 1896 :   1 - 0x1 -- plane 1
      12'h769: dout <= 8'b00000011; // 1897 :   3 - 0x3
      12'h76A: dout <= 8'b00000011; // 1898 :   3 - 0x3
      12'h76B: dout <= 8'b00000111; // 1899 :   7 - 0x7
      12'h76C: dout <= 8'b00000100; // 1900 :   4 - 0x4
      12'h76D: dout <= 8'b00011100; // 1901 :  28 - 0x1c
      12'h76E: dout <= 8'b00111111; // 1902 :  63 - 0x3f
      12'h76F: dout <= 8'b01111111; // 1903 : 127 - 0x7f
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Background 0x77
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b01111100; // 1906 : 124 - 0x7c
      12'h773: dout <= 8'b00000010; // 1907 :   2 - 0x2
      12'h774: dout <= 8'b00000001; // 1908 :   1 - 0x1
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b01111111; // 1912 : 127 - 0x7f -- plane 1
      12'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      12'h77A: dout <= 8'b11111111; // 1914 : 255 - 0xff
      12'h77B: dout <= 8'b01111111; // 1915 : 127 - 0x7f
      12'h77C: dout <= 8'b01111111; // 1916 : 127 - 0x7f
      12'h77D: dout <= 8'b00011111; // 1917 :  31 - 0x1f
      12'h77E: dout <= 8'b00000011; // 1918 :   3 - 0x3
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Background 0x78
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000001; // 1922 :   1 - 0x1
      12'h783: dout <= 8'b00000001; // 1923 :   1 - 0x1
      12'h784: dout <= 8'b00000011; // 1924 :   3 - 0x3
      12'h785: dout <= 8'b00000111; // 1925 :   7 - 0x7
      12'h786: dout <= 8'b00000111; // 1926 :   7 - 0x7
      12'h787: dout <= 8'b00001111; // 1927 :  15 - 0xf
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000001; // 1930 :   1 - 0x1
      12'h78B: dout <= 8'b00000001; // 1931 :   1 - 0x1
      12'h78C: dout <= 8'b00000011; // 1932 :   3 - 0x3
      12'h78D: dout <= 8'b00000111; // 1933 :   7 - 0x7
      12'h78E: dout <= 8'b00000111; // 1934 :   7 - 0x7
      12'h78F: dout <= 8'b00001111; // 1935 :  15 - 0xf
      12'h790: dout <= 8'b00001111; // 1936 :  15 - 0xf -- Background 0x79
      12'h791: dout <= 8'b00000111; // 1937 :   7 - 0x7
      12'h792: dout <= 8'b00001111; // 1938 :  15 - 0xf
      12'h793: dout <= 8'b00000111; // 1939 :   7 - 0x7
      12'h794: dout <= 8'b00000001; // 1940 :   1 - 0x1
      12'h795: dout <= 8'b00010000; // 1941 :  16 - 0x10
      12'h796: dout <= 8'b00100000; // 1942 :  32 - 0x20
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b11111111; // 1944 : 255 - 0xff -- plane 1
      12'h799: dout <= 8'b11111111; // 1945 : 255 - 0xff
      12'h79A: dout <= 8'b00111111; // 1946 :  63 - 0x3f
      12'h79B: dout <= 8'b00111111; // 1947 :  63 - 0x3f
      12'h79C: dout <= 8'b01111111; // 1948 : 127 - 0x7f
      12'h79D: dout <= 8'b11111110; // 1949 : 254 - 0xfe
      12'h79E: dout <= 8'b11111100; // 1950 : 252 - 0xfc
      12'h79F: dout <= 8'b00110000; // 1951 :  48 - 0x30
      12'h7A0: dout <= 8'b11111000; // 1952 : 248 - 0xf8 -- Background 0x7a
      12'h7A1: dout <= 8'b11111110; // 1953 : 254 - 0xfe
      12'h7A2: dout <= 8'b01111111; // 1954 : 127 - 0x7f
      12'h7A3: dout <= 8'b00011111; // 1955 :  31 - 0x1f
      12'h7A4: dout <= 8'b00001111; // 1956 :  15 - 0xf
      12'h7A5: dout <= 8'b00011001; // 1957 :  25 - 0x19
      12'h7A6: dout <= 8'b00110000; // 1958 :  48 - 0x30
      12'h7A7: dout <= 8'b01110000; // 1959 : 112 - 0x70
      12'h7A8: dout <= 8'b11111000; // 1960 : 248 - 0xf8 -- plane 1
      12'h7A9: dout <= 8'b11111110; // 1961 : 254 - 0xfe
      12'h7AA: dout <= 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout <= 8'b11111111; // 1963 : 255 - 0xff
      12'h7AC: dout <= 8'b11111111; // 1964 : 255 - 0xff
      12'h7AD: dout <= 8'b11111111; // 1965 : 255 - 0xff
      12'h7AE: dout <= 8'b11111111; // 1966 : 255 - 0xff
      12'h7AF: dout <= 8'b11111111; // 1967 : 255 - 0xff
      12'h7B0: dout <= 8'b11111011; // 1968 : 251 - 0xfb -- Background 0x7b
      12'h7B1: dout <= 8'b01110011; // 1969 : 115 - 0x73
      12'h7B2: dout <= 8'b00100111; // 1970 :  39 - 0x27
      12'h7B3: dout <= 8'b00001111; // 1971 :  15 - 0xf
      12'h7B4: dout <= 8'b00011111; // 1972 :  31 - 0x1f
      12'h7B5: dout <= 8'b00011111; // 1973 :  31 - 0x1f
      12'h7B6: dout <= 8'b00111111; // 1974 :  63 - 0x3f
      12'h7B7: dout <= 8'b01111111; // 1975 : 127 - 0x7f
      12'h7B8: dout <= 8'b11111111; // 1976 : 255 - 0xff -- plane 1
      12'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      12'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      12'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      12'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      12'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      12'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      12'h7BF: dout <= 8'b01111111; // 1983 : 127 - 0x7f
      12'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Background 0x7c
      12'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout <= 8'b11111110; // 1988 : 254 - 0xfe
      12'h7C5: dout <= 8'b11111101; // 1989 : 253 - 0xfd
      12'h7C6: dout <= 8'b11111000; // 1990 : 248 - 0xf8
      12'h7C7: dout <= 8'b11110110; // 1991 : 246 - 0xf6
      12'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- plane 1
      12'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      12'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      12'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      12'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      12'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout <= 8'b11101111; // 2000 : 239 - 0xef -- Background 0x7d
      12'h7D1: dout <= 8'b11001111; // 2001 : 207 - 0xcf
      12'h7D2: dout <= 8'b10011111; // 2002 : 159 - 0x9f
      12'h7D3: dout <= 8'b00011111; // 2003 :  31 - 0x1f
      12'h7D4: dout <= 8'b00001111; // 2004 :  15 - 0xf
      12'h7D5: dout <= 8'b00101101; // 2005 :  45 - 0x2d
      12'h7D6: dout <= 8'b01010000; // 2006 :  80 - 0x50
      12'h7D7: dout <= 8'b01000000; // 2007 :  64 - 0x40
      12'h7D8: dout <= 8'b11101111; // 2008 : 239 - 0xef -- plane 1
      12'h7D9: dout <= 8'b11001111; // 2009 : 207 - 0xcf
      12'h7DA: dout <= 8'b10011111; // 2010 : 159 - 0x9f
      12'h7DB: dout <= 8'b00011111; // 2011 :  31 - 0x1f
      12'h7DC: dout <= 8'b00001111; // 2012 :  15 - 0xf
      12'h7DD: dout <= 8'b01111111; // 2013 : 127 - 0x7f
      12'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      12'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Background 0x7e
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout <= 8'b11100000; // 2020 : 224 - 0xe0
      12'h7E5: dout <= 8'b11111110; // 2021 : 254 - 0xfe
      12'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout <= 8'b11110011; // 2023 : 243 - 0xf3
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- plane 1
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout <= 8'b11110000; // 2027 : 240 - 0xf0
      12'h7EC: dout <= 8'b11111110; // 2028 : 254 - 0xfe
      12'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      12'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      12'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout <= 8'b11111011; // 2032 : 251 - 0xfb -- Background 0x7f
      12'h7F1: dout <= 8'b11111011; // 2033 : 251 - 0xfb
      12'h7F2: dout <= 8'b11111011; // 2034 : 251 - 0xfb
      12'h7F3: dout <= 8'b11111011; // 2035 : 251 - 0xfb
      12'h7F4: dout <= 8'b11111011; // 2036 : 251 - 0xfb
      12'h7F5: dout <= 8'b11110011; // 2037 : 243 - 0xf3
      12'h7F6: dout <= 8'b11110111; // 2038 : 247 - 0xf7
      12'h7F7: dout <= 8'b11100111; // 2039 : 231 - 0xe7
      12'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- plane 1
      12'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      12'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      12'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      12'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      12'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      12'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
      12'h800: dout <= 8'b11001111; // 2048 : 207 - 0xcf -- Background 0x80
      12'h801: dout <= 8'b10011111; // 2049 : 159 - 0x9f
      12'h802: dout <= 8'b00111111; // 2050 :  63 - 0x3f
      12'h803: dout <= 8'b00111111; // 2051 :  63 - 0x3f
      12'h804: dout <= 8'b00111111; // 2052 :  63 - 0x3f
      12'h805: dout <= 8'b00001111; // 2053 :  15 - 0xf
      12'h806: dout <= 8'b00000011; // 2054 :   3 - 0x3
      12'h807: dout <= 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout <= 8'b11111111; // 2056 : 255 - 0xff -- plane 1
      12'h809: dout <= 8'b11111111; // 2057 : 255 - 0xff
      12'h80A: dout <= 8'b11111111; // 2058 : 255 - 0xff
      12'h80B: dout <= 8'b11111111; // 2059 : 255 - 0xff
      12'h80C: dout <= 8'b11111111; // 2060 : 255 - 0xff
      12'h80D: dout <= 8'b11111111; // 2061 : 255 - 0xff
      12'h80E: dout <= 8'b11111111; // 2062 : 255 - 0xff
      12'h80F: dout <= 8'b11111111; // 2063 : 255 - 0xff
      12'h810: dout <= 8'b11000000; // 2064 : 192 - 0xc0 -- Background 0x81
      12'h811: dout <= 8'b11110000; // 2065 : 240 - 0xf0
      12'h812: dout <= 8'b11111100; // 2066 : 252 - 0xfc
      12'h813: dout <= 8'b11110000; // 2067 : 240 - 0xf0
      12'h814: dout <= 8'b11110000; // 2068 : 240 - 0xf0
      12'h815: dout <= 8'b10011000; // 2069 : 152 - 0x98
      12'h816: dout <= 8'b00001000; // 2070 :   8 - 0x8
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b11111111; // 2072 : 255 - 0xff -- plane 1
      12'h819: dout <= 8'b11111111; // 2073 : 255 - 0xff
      12'h81A: dout <= 8'b11111111; // 2074 : 255 - 0xff
      12'h81B: dout <= 8'b11110000; // 2075 : 240 - 0xf0
      12'h81C: dout <= 8'b11110000; // 2076 : 240 - 0xf0
      12'h81D: dout <= 8'b11111000; // 2077 : 248 - 0xf8
      12'h81E: dout <= 8'b11111000; // 2078 : 248 - 0xf8
      12'h81F: dout <= 8'b11111000; // 2079 : 248 - 0xf8
      12'h820: dout <= 8'b00000000; // 2080 :   0 - 0x0 -- Background 0x82
      12'h821: dout <= 8'b00000000; // 2081 :   0 - 0x0
      12'h822: dout <= 8'b00000000; // 2082 :   0 - 0x0
      12'h823: dout <= 8'b00000000; // 2083 :   0 - 0x0
      12'h824: dout <= 8'b00000000; // 2084 :   0 - 0x0
      12'h825: dout <= 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout <= 8'b10000000; // 2086 : 128 - 0x80
      12'h827: dout <= 8'b11000000; // 2087 : 192 - 0xc0
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout <= 8'b10000000; // 2093 : 128 - 0x80
      12'h82E: dout <= 8'b11000000; // 2094 : 192 - 0xc0
      12'h82F: dout <= 8'b11100000; // 2095 : 224 - 0xe0
      12'h830: dout <= 8'b11100000; // 2096 : 224 - 0xe0 -- Background 0x83
      12'h831: dout <= 8'b11100000; // 2097 : 224 - 0xe0
      12'h832: dout <= 8'b11110000; // 2098 : 240 - 0xf0
      12'h833: dout <= 8'b11110000; // 2099 : 240 - 0xf0
      12'h834: dout <= 8'b11110000; // 2100 : 240 - 0xf0
      12'h835: dout <= 8'b11110000; // 2101 : 240 - 0xf0
      12'h836: dout <= 8'b11111000; // 2102 : 248 - 0xf8
      12'h837: dout <= 8'b11111000; // 2103 : 248 - 0xf8
      12'h838: dout <= 8'b11110000; // 2104 : 240 - 0xf0 -- plane 1
      12'h839: dout <= 8'b11110000; // 2105 : 240 - 0xf0
      12'h83A: dout <= 8'b11111000; // 2106 : 248 - 0xf8
      12'h83B: dout <= 8'b11111000; // 2107 : 248 - 0xf8
      12'h83C: dout <= 8'b11111000; // 2108 : 248 - 0xf8
      12'h83D: dout <= 8'b11111100; // 2109 : 252 - 0xfc
      12'h83E: dout <= 8'b11111100; // 2110 : 252 - 0xfc
      12'h83F: dout <= 8'b11111110; // 2111 : 254 - 0xfe
      12'h840: dout <= 8'b11111110; // 2112 : 254 - 0xfe -- Background 0x84
      12'h841: dout <= 8'b11111111; // 2113 : 255 - 0xff
      12'h842: dout <= 8'b11111111; // 2114 : 255 - 0xff
      12'h843: dout <= 8'b11111111; // 2115 : 255 - 0xff
      12'h844: dout <= 8'b11111111; // 2116 : 255 - 0xff
      12'h845: dout <= 8'b11111111; // 2117 : 255 - 0xff
      12'h846: dout <= 8'b11111111; // 2118 : 255 - 0xff
      12'h847: dout <= 8'b11111111; // 2119 : 255 - 0xff
      12'h848: dout <= 8'b11111111; // 2120 : 255 - 0xff -- plane 1
      12'h849: dout <= 8'b11111111; // 2121 : 255 - 0xff
      12'h84A: dout <= 8'b11111111; // 2122 : 255 - 0xff
      12'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      12'h84C: dout <= 8'b11111111; // 2124 : 255 - 0xff
      12'h84D: dout <= 8'b11111111; // 2125 : 255 - 0xff
      12'h84E: dout <= 8'b11111111; // 2126 : 255 - 0xff
      12'h84F: dout <= 8'b11111111; // 2127 : 255 - 0xff
      12'h850: dout <= 8'b00111111; // 2128 :  63 - 0x3f -- Background 0x85
      12'h851: dout <= 8'b00011111; // 2129 :  31 - 0x1f
      12'h852: dout <= 8'b00011111; // 2130 :  31 - 0x1f
      12'h853: dout <= 8'b00001111; // 2131 :  15 - 0xf
      12'h854: dout <= 8'b00000111; // 2132 :   7 - 0x7
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b11111111; // 2136 : 255 - 0xff -- plane 1
      12'h859: dout <= 8'b11111111; // 2137 : 255 - 0xff
      12'h85A: dout <= 8'b11111111; // 2138 : 255 - 0xff
      12'h85B: dout <= 8'b00001111; // 2139 :  15 - 0xf
      12'h85C: dout <= 8'b00000111; // 2140 :   7 - 0x7
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b00000000; // 2144 :   0 - 0x0 -- Background 0x86
      12'h861: dout <= 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout <= 8'b11000000; // 2146 : 192 - 0xc0
      12'h863: dout <= 8'b11100000; // 2147 : 224 - 0xe0
      12'h864: dout <= 8'b11110000; // 2148 : 240 - 0xf0
      12'h865: dout <= 8'b11110000; // 2149 : 240 - 0xf0
      12'h866: dout <= 8'b11110000; // 2150 : 240 - 0xf0
      12'h867: dout <= 8'b11111000; // 2151 : 248 - 0xf8
      12'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout <= 8'b10000000; // 2153 : 128 - 0x80
      12'h86A: dout <= 8'b11000000; // 2154 : 192 - 0xc0
      12'h86B: dout <= 8'b11100000; // 2155 : 224 - 0xe0
      12'h86C: dout <= 8'b11110000; // 2156 : 240 - 0xf0
      12'h86D: dout <= 8'b11110000; // 2157 : 240 - 0xf0
      12'h86E: dout <= 8'b11110000; // 2158 : 240 - 0xf0
      12'h86F: dout <= 8'b11111100; // 2159 : 252 - 0xfc
      12'h870: dout <= 8'b11111001; // 2160 : 249 - 0xf9 -- Background 0x87
      12'h871: dout <= 8'b11111111; // 2161 : 255 - 0xff
      12'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout <= 8'b11111111; // 2164 : 255 - 0xff
      12'h875: dout <= 8'b00001110; // 2165 :  14 - 0xe
      12'h876: dout <= 8'b00000010; // 2166 :   2 - 0x2
      12'h877: dout <= 8'b00010100; // 2167 :  20 - 0x14
      12'h878: dout <= 8'b11111111; // 2168 : 255 - 0xff -- plane 1
      12'h879: dout <= 8'b11111111; // 2169 : 255 - 0xff
      12'h87A: dout <= 8'b11111111; // 2170 : 255 - 0xff
      12'h87B: dout <= 8'b11111111; // 2171 : 255 - 0xff
      12'h87C: dout <= 8'b11111111; // 2172 : 255 - 0xff
      12'h87D: dout <= 8'b00001111; // 2173 :  15 - 0xf
      12'h87E: dout <= 8'b00011111; // 2174 :  31 - 0x1f
      12'h87F: dout <= 8'b00111111; // 2175 :  63 - 0x3f
      12'h880: dout <= 8'b10000000; // 2176 : 128 - 0x80 -- Background 0x88
      12'h881: dout <= 8'b10100000; // 2177 : 160 - 0xa0
      12'h882: dout <= 8'b00100000; // 2178 :  32 - 0x20
      12'h883: dout <= 8'b00100000; // 2179 :  32 - 0x20
      12'h884: dout <= 8'b10100000; // 2180 : 160 - 0xa0
      12'h885: dout <= 8'b10000000; // 2181 : 128 - 0x80
      12'h886: dout <= 8'b00000000; // 2182 :   0 - 0x0
      12'h887: dout <= 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout <= 8'b11000000; // 2184 : 192 - 0xc0 -- plane 1
      12'h889: dout <= 8'b11100000; // 2185 : 224 - 0xe0
      12'h88A: dout <= 8'b11100000; // 2186 : 224 - 0xe0
      12'h88B: dout <= 8'b11100000; // 2187 : 224 - 0xe0
      12'h88C: dout <= 8'b11100000; // 2188 : 224 - 0xe0
      12'h88D: dout <= 8'b11000000; // 2189 : 192 - 0xc0
      12'h88E: dout <= 8'b11000000; // 2190 : 192 - 0xc0
      12'h88F: dout <= 8'b10000000; // 2191 : 128 - 0x80
      12'h890: dout <= 8'b00000001; // 2192 :   1 - 0x1 -- Background 0x89
      12'h891: dout <= 8'b00000101; // 2193 :   5 - 0x5
      12'h892: dout <= 8'b00000100; // 2194 :   4 - 0x4
      12'h893: dout <= 8'b00000100; // 2195 :   4 - 0x4
      12'h894: dout <= 8'b00000101; // 2196 :   5 - 0x5
      12'h895: dout <= 8'b00000001; // 2197 :   1 - 0x1
      12'h896: dout <= 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00000011; // 2200 :   3 - 0x3 -- plane 1
      12'h899: dout <= 8'b00000111; // 2201 :   7 - 0x7
      12'h89A: dout <= 8'b00000111; // 2202 :   7 - 0x7
      12'h89B: dout <= 8'b00000111; // 2203 :   7 - 0x7
      12'h89C: dout <= 8'b00000111; // 2204 :   7 - 0x7
      12'h89D: dout <= 8'b00000011; // 2205 :   3 - 0x3
      12'h89E: dout <= 8'b00000011; // 2206 :   3 - 0x3
      12'h89F: dout <= 8'b00000001; // 2207 :   1 - 0x1
      12'h8A0: dout <= 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x8a
      12'h8A1: dout <= 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout <= 8'b00000011; // 2210 :   3 - 0x3
      12'h8A3: dout <= 8'b00000111; // 2211 :   7 - 0x7
      12'h8A4: dout <= 8'b00001111; // 2212 :  15 - 0xf
      12'h8A5: dout <= 8'b00001111; // 2213 :  15 - 0xf
      12'h8A6: dout <= 8'b00001111; // 2214 :  15 - 0xf
      12'h8A7: dout <= 8'b00001111; // 2215 :  15 - 0xf
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout <= 8'b00000001; // 2217 :   1 - 0x1
      12'h8AA: dout <= 8'b00000011; // 2218 :   3 - 0x3
      12'h8AB: dout <= 8'b00000111; // 2219 :   7 - 0x7
      12'h8AC: dout <= 8'b00001111; // 2220 :  15 - 0xf
      12'h8AD: dout <= 8'b00001111; // 2221 :  15 - 0xf
      12'h8AE: dout <= 8'b00001111; // 2222 :  15 - 0xf
      12'h8AF: dout <= 8'b00111111; // 2223 :  63 - 0x3f
      12'h8B0: dout <= 8'b10011111; // 2224 : 159 - 0x9f -- Background 0x8b
      12'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout <= 8'b11111111; // 2226 : 255 - 0xff
      12'h8B3: dout <= 8'b11111111; // 2227 : 255 - 0xff
      12'h8B4: dout <= 8'b11111111; // 2228 : 255 - 0xff
      12'h8B5: dout <= 8'b01110000; // 2229 : 112 - 0x70
      12'h8B6: dout <= 8'b01000000; // 2230 :  64 - 0x40
      12'h8B7: dout <= 8'b00101000; // 2231 :  40 - 0x28
      12'h8B8: dout <= 8'b11111111; // 2232 : 255 - 0xff -- plane 1
      12'h8B9: dout <= 8'b11111111; // 2233 : 255 - 0xff
      12'h8BA: dout <= 8'b11111111; // 2234 : 255 - 0xff
      12'h8BB: dout <= 8'b11111111; // 2235 : 255 - 0xff
      12'h8BC: dout <= 8'b11111111; // 2236 : 255 - 0xff
      12'h8BD: dout <= 8'b11110000; // 2237 : 240 - 0xf0
      12'h8BE: dout <= 8'b11111000; // 2238 : 248 - 0xf8
      12'h8BF: dout <= 8'b11111100; // 2239 : 252 - 0xfc
      12'h8C0: dout <= 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x8c
      12'h8C1: dout <= 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout <= 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00000000; // 2244 :   0 - 0x0
      12'h8C5: dout <= 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout <= 8'b00000001; // 2246 :   1 - 0x1
      12'h8C7: dout <= 8'b00000011; // 2247 :   3 - 0x3
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout <= 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout <= 8'b00000001; // 2253 :   1 - 0x1
      12'h8CE: dout <= 8'b00000011; // 2254 :   3 - 0x3
      12'h8CF: dout <= 8'b00000111; // 2255 :   7 - 0x7
      12'h8D0: dout <= 8'b00000111; // 2256 :   7 - 0x7 -- Background 0x8d
      12'h8D1: dout <= 8'b00000111; // 2257 :   7 - 0x7
      12'h8D2: dout <= 8'b00001111; // 2258 :  15 - 0xf
      12'h8D3: dout <= 8'b00001111; // 2259 :  15 - 0xf
      12'h8D4: dout <= 8'b00001111; // 2260 :  15 - 0xf
      12'h8D5: dout <= 8'b00001111; // 2261 :  15 - 0xf
      12'h8D6: dout <= 8'b00011111; // 2262 :  31 - 0x1f
      12'h8D7: dout <= 8'b00011111; // 2263 :  31 - 0x1f
      12'h8D8: dout <= 8'b00001111; // 2264 :  15 - 0xf -- plane 1
      12'h8D9: dout <= 8'b00001111; // 2265 :  15 - 0xf
      12'h8DA: dout <= 8'b00011111; // 2266 :  31 - 0x1f
      12'h8DB: dout <= 8'b00011111; // 2267 :  31 - 0x1f
      12'h8DC: dout <= 8'b00011111; // 2268 :  31 - 0x1f
      12'h8DD: dout <= 8'b00111111; // 2269 :  63 - 0x3f
      12'h8DE: dout <= 8'b00111111; // 2270 :  63 - 0x3f
      12'h8DF: dout <= 8'b01111111; // 2271 : 127 - 0x7f
      12'h8E0: dout <= 8'b01111111; // 2272 : 127 - 0x7f -- Background 0x8e
      12'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout <= 8'b11111111; // 2274 : 255 - 0xff
      12'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      12'h8E4: dout <= 8'b11111111; // 2276 : 255 - 0xff
      12'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      12'h8E6: dout <= 8'b11111111; // 2278 : 255 - 0xff
      12'h8E7: dout <= 8'b11111111; // 2279 : 255 - 0xff
      12'h8E8: dout <= 8'b11111111; // 2280 : 255 - 0xff -- plane 1
      12'h8E9: dout <= 8'b11111111; // 2281 : 255 - 0xff
      12'h8EA: dout <= 8'b11111111; // 2282 : 255 - 0xff
      12'h8EB: dout <= 8'b11111111; // 2283 : 255 - 0xff
      12'h8EC: dout <= 8'b11111111; // 2284 : 255 - 0xff
      12'h8ED: dout <= 8'b11111111; // 2285 : 255 - 0xff
      12'h8EE: dout <= 8'b11111111; // 2286 : 255 - 0xff
      12'h8EF: dout <= 8'b11111111; // 2287 : 255 - 0xff
      12'h8F0: dout <= 8'b11111100; // 2288 : 252 - 0xfc -- Background 0x8f
      12'h8F1: dout <= 8'b11111000; // 2289 : 248 - 0xf8
      12'h8F2: dout <= 8'b11111000; // 2290 : 248 - 0xf8
      12'h8F3: dout <= 8'b11110000; // 2291 : 240 - 0xf0
      12'h8F4: dout <= 8'b11100000; // 2292 : 224 - 0xe0
      12'h8F5: dout <= 8'b00000000; // 2293 :   0 - 0x0
      12'h8F6: dout <= 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout <= 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout <= 8'b11111111; // 2296 : 255 - 0xff -- plane 1
      12'h8F9: dout <= 8'b11111111; // 2297 : 255 - 0xff
      12'h8FA: dout <= 8'b11111111; // 2298 : 255 - 0xff
      12'h8FB: dout <= 8'b11110000; // 2299 : 240 - 0xf0
      12'h8FC: dout <= 8'b11100000; // 2300 : 224 - 0xe0
      12'h8FD: dout <= 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout <= 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x90
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout <= 8'b00000111; // 2308 :   7 - 0x7
      12'h905: dout <= 8'b01111111; // 2309 : 127 - 0x7f
      12'h906: dout <= 8'b11111111; // 2310 : 255 - 0xff
      12'h907: dout <= 8'b11001111; // 2311 : 207 - 0xcf
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00001111; // 2315 :  15 - 0xf
      12'h90C: dout <= 8'b01111111; // 2316 : 127 - 0x7f
      12'h90D: dout <= 8'b11111111; // 2317 : 255 - 0xff
      12'h90E: dout <= 8'b11111111; // 2318 : 255 - 0xff
      12'h90F: dout <= 8'b11111111; // 2319 : 255 - 0xff
      12'h910: dout <= 8'b11011111; // 2320 : 223 - 0xdf -- Background 0x91
      12'h911: dout <= 8'b11011111; // 2321 : 223 - 0xdf
      12'h912: dout <= 8'b11011111; // 2322 : 223 - 0xdf
      12'h913: dout <= 8'b11011111; // 2323 : 223 - 0xdf
      12'h914: dout <= 8'b11011111; // 2324 : 223 - 0xdf
      12'h915: dout <= 8'b11001111; // 2325 : 207 - 0xcf
      12'h916: dout <= 8'b11101111; // 2326 : 239 - 0xef
      12'h917: dout <= 8'b11100111; // 2327 : 231 - 0xe7
      12'h918: dout <= 8'b11111111; // 2328 : 255 - 0xff -- plane 1
      12'h919: dout <= 8'b11111111; // 2329 : 255 - 0xff
      12'h91A: dout <= 8'b11111111; // 2330 : 255 - 0xff
      12'h91B: dout <= 8'b11111111; // 2331 : 255 - 0xff
      12'h91C: dout <= 8'b11111111; // 2332 : 255 - 0xff
      12'h91D: dout <= 8'b11111111; // 2333 : 255 - 0xff
      12'h91E: dout <= 8'b11111111; // 2334 : 255 - 0xff
      12'h91F: dout <= 8'b11111111; // 2335 : 255 - 0xff
      12'h920: dout <= 8'b11110011; // 2336 : 243 - 0xf3 -- Background 0x92
      12'h921: dout <= 8'b11111001; // 2337 : 249 - 0xf9
      12'h922: dout <= 8'b11111100; // 2338 : 252 - 0xfc
      12'h923: dout <= 8'b11111100; // 2339 : 252 - 0xfc
      12'h924: dout <= 8'b11111100; // 2340 : 252 - 0xfc
      12'h925: dout <= 8'b11110000; // 2341 : 240 - 0xf0
      12'h926: dout <= 8'b11000000; // 2342 : 192 - 0xc0
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b11111111; // 2344 : 255 - 0xff -- plane 1
      12'h929: dout <= 8'b11111111; // 2345 : 255 - 0xff
      12'h92A: dout <= 8'b11111111; // 2346 : 255 - 0xff
      12'h92B: dout <= 8'b11111111; // 2347 : 255 - 0xff
      12'h92C: dout <= 8'b11111111; // 2348 : 255 - 0xff
      12'h92D: dout <= 8'b11111111; // 2349 : 255 - 0xff
      12'h92E: dout <= 8'b11111111; // 2350 : 255 - 0xff
      12'h92F: dout <= 8'b11111111; // 2351 : 255 - 0xff
      12'h930: dout <= 8'b00000011; // 2352 :   3 - 0x3 -- Background 0x93
      12'h931: dout <= 8'b00001111; // 2353 :  15 - 0xf
      12'h932: dout <= 8'b00111111; // 2354 :  63 - 0x3f
      12'h933: dout <= 8'b00001111; // 2355 :  15 - 0xf
      12'h934: dout <= 8'b00001111; // 2356 :  15 - 0xf
      12'h935: dout <= 8'b00011001; // 2357 :  25 - 0x19
      12'h936: dout <= 8'b00010000; // 2358 :  16 - 0x10
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b11111111; // 2360 : 255 - 0xff -- plane 1
      12'h939: dout <= 8'b11111111; // 2361 : 255 - 0xff
      12'h93A: dout <= 8'b11111111; // 2362 : 255 - 0xff
      12'h93B: dout <= 8'b00001111; // 2363 :  15 - 0xf
      12'h93C: dout <= 8'b00001111; // 2364 :  15 - 0xf
      12'h93D: dout <= 8'b00011111; // 2365 :  31 - 0x1f
      12'h93E: dout <= 8'b00011111; // 2366 :  31 - 0x1f
      12'h93F: dout <= 8'b00011111; // 2367 :  31 - 0x1f
      12'h940: dout <= 8'b00011111; // 2368 :  31 - 0x1f -- Background 0x94
      12'h941: dout <= 8'b01111111; // 2369 : 127 - 0x7f
      12'h942: dout <= 8'b11111110; // 2370 : 254 - 0xfe
      12'h943: dout <= 8'b11111000; // 2371 : 248 - 0xf8
      12'h944: dout <= 8'b11110000; // 2372 : 240 - 0xf0
      12'h945: dout <= 8'b10011000; // 2373 : 152 - 0x98
      12'h946: dout <= 8'b00001100; // 2374 :  12 - 0xc
      12'h947: dout <= 8'b00001110; // 2375 :  14 - 0xe
      12'h948: dout <= 8'b00011111; // 2376 :  31 - 0x1f -- plane 1
      12'h949: dout <= 8'b01111111; // 2377 : 127 - 0x7f
      12'h94A: dout <= 8'b11111111; // 2378 : 255 - 0xff
      12'h94B: dout <= 8'b11111111; // 2379 : 255 - 0xff
      12'h94C: dout <= 8'b11111111; // 2380 : 255 - 0xff
      12'h94D: dout <= 8'b11111111; // 2381 : 255 - 0xff
      12'h94E: dout <= 8'b11111111; // 2382 : 255 - 0xff
      12'h94F: dout <= 8'b11111111; // 2383 : 255 - 0xff
      12'h950: dout <= 8'b11011111; // 2384 : 223 - 0xdf -- Background 0x95
      12'h951: dout <= 8'b11001110; // 2385 : 206 - 0xce
      12'h952: dout <= 8'b11100100; // 2386 : 228 - 0xe4
      12'h953: dout <= 8'b11110000; // 2387 : 240 - 0xf0
      12'h954: dout <= 8'b11111000; // 2388 : 248 - 0xf8
      12'h955: dout <= 8'b11111000; // 2389 : 248 - 0xf8
      12'h956: dout <= 8'b11111100; // 2390 : 252 - 0xfc
      12'h957: dout <= 8'b11111110; // 2391 : 254 - 0xfe
      12'h958: dout <= 8'b11111111; // 2392 : 255 - 0xff -- plane 1
      12'h959: dout <= 8'b11111111; // 2393 : 255 - 0xff
      12'h95A: dout <= 8'b11111111; // 2394 : 255 - 0xff
      12'h95B: dout <= 8'b11111111; // 2395 : 255 - 0xff
      12'h95C: dout <= 8'b11111111; // 2396 : 255 - 0xff
      12'h95D: dout <= 8'b11111111; // 2397 : 255 - 0xff
      12'h95E: dout <= 8'b11111111; // 2398 : 255 - 0xff
      12'h95F: dout <= 8'b11111110; // 2399 : 254 - 0xfe
      12'h960: dout <= 8'b11111111; // 2400 : 255 - 0xff -- Background 0x96
      12'h961: dout <= 8'b11111111; // 2401 : 255 - 0xff
      12'h962: dout <= 8'b11111111; // 2402 : 255 - 0xff
      12'h963: dout <= 8'b11111111; // 2403 : 255 - 0xff
      12'h964: dout <= 8'b01111111; // 2404 : 127 - 0x7f
      12'h965: dout <= 8'b10111111; // 2405 : 191 - 0xbf
      12'h966: dout <= 8'b00011111; // 2406 :  31 - 0x1f
      12'h967: dout <= 8'b01101111; // 2407 : 111 - 0x6f
      12'h968: dout <= 8'b11111111; // 2408 : 255 - 0xff -- plane 1
      12'h969: dout <= 8'b11111111; // 2409 : 255 - 0xff
      12'h96A: dout <= 8'b11111111; // 2410 : 255 - 0xff
      12'h96B: dout <= 8'b11111111; // 2411 : 255 - 0xff
      12'h96C: dout <= 8'b11111111; // 2412 : 255 - 0xff
      12'h96D: dout <= 8'b11111111; // 2413 : 255 - 0xff
      12'h96E: dout <= 8'b11111111; // 2414 : 255 - 0xff
      12'h96F: dout <= 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout <= 8'b11110111; // 2416 : 247 - 0xf7 -- Background 0x97
      12'h971: dout <= 8'b11110011; // 2417 : 243 - 0xf3
      12'h972: dout <= 8'b11111001; // 2418 : 249 - 0xf9
      12'h973: dout <= 8'b11111000; // 2419 : 248 - 0xf8
      12'h974: dout <= 8'b11110000; // 2420 : 240 - 0xf0
      12'h975: dout <= 8'b10110100; // 2421 : 180 - 0xb4
      12'h976: dout <= 8'b00001010; // 2422 :  10 - 0xa
      12'h977: dout <= 8'b00000010; // 2423 :   2 - 0x2
      12'h978: dout <= 8'b11110111; // 2424 : 247 - 0xf7 -- plane 1
      12'h979: dout <= 8'b11110011; // 2425 : 243 - 0xf3
      12'h97A: dout <= 8'b11111001; // 2426 : 249 - 0xf9
      12'h97B: dout <= 8'b11111000; // 2427 : 248 - 0xf8
      12'h97C: dout <= 8'b11110000; // 2428 : 240 - 0xf0
      12'h97D: dout <= 8'b11111110; // 2429 : 254 - 0xfe
      12'h97E: dout <= 8'b11111111; // 2430 : 255 - 0xff
      12'h97F: dout <= 8'b11111111; // 2431 : 255 - 0xff
      12'h980: dout <= 8'b10000000; // 2432 : 128 - 0x80 -- Background 0x98
      12'h981: dout <= 8'b11000000; // 2433 : 192 - 0xc0
      12'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout <= 8'b00000000; // 2435 :   0 - 0x0
      12'h984: dout <= 8'b11000000; // 2436 : 192 - 0xc0
      12'h985: dout <= 8'b10011000; // 2437 : 152 - 0x98
      12'h986: dout <= 8'b00000000; // 2438 :   0 - 0x0
      12'h987: dout <= 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout <= 8'b10000000; // 2440 : 128 - 0x80 -- plane 1
      12'h989: dout <= 8'b11000000; // 2441 : 192 - 0xc0
      12'h98A: dout <= 8'b11000000; // 2442 : 192 - 0xc0
      12'h98B: dout <= 8'b11100000; // 2443 : 224 - 0xe0
      12'h98C: dout <= 8'b00100000; // 2444 :  32 - 0x20
      12'h98D: dout <= 8'b00111000; // 2445 :  56 - 0x38
      12'h98E: dout <= 8'b11111100; // 2446 : 252 - 0xfc
      12'h98F: dout <= 8'b11111110; // 2447 : 254 - 0xfe
      12'h990: dout <= 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x99
      12'h991: dout <= 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout <= 8'b00111110; // 2450 :  62 - 0x3e
      12'h993: dout <= 8'b01000000; // 2451 :  64 - 0x40
      12'h994: dout <= 8'b10000000; // 2452 : 128 - 0x80
      12'h995: dout <= 8'b00000000; // 2453 :   0 - 0x0
      12'h996: dout <= 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout <= 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout <= 8'b11111110; // 2456 : 254 - 0xfe -- plane 1
      12'h999: dout <= 8'b11111111; // 2457 : 255 - 0xff
      12'h99A: dout <= 8'b11111111; // 2458 : 255 - 0xff
      12'h99B: dout <= 8'b11111110; // 2459 : 254 - 0xfe
      12'h99C: dout <= 8'b11111100; // 2460 : 252 - 0xfc
      12'h99D: dout <= 8'b11111000; // 2461 : 248 - 0xf8
      12'h99E: dout <= 8'b11000000; // 2462 : 192 - 0xc0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x9a
      12'h9A1: dout <= 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout <= 8'b10000000; // 2466 : 128 - 0x80
      12'h9A3: dout <= 8'b10000000; // 2467 : 128 - 0x80
      12'h9A4: dout <= 8'b11000000; // 2468 : 192 - 0xc0
      12'h9A5: dout <= 8'b11100000; // 2469 : 224 - 0xe0
      12'h9A6: dout <= 8'b11100000; // 2470 : 224 - 0xe0
      12'h9A7: dout <= 8'b11110000; // 2471 : 240 - 0xf0
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b10000000; // 2474 : 128 - 0x80
      12'h9AB: dout <= 8'b10000000; // 2475 : 128 - 0x80
      12'h9AC: dout <= 8'b11000000; // 2476 : 192 - 0xc0
      12'h9AD: dout <= 8'b11100000; // 2477 : 224 - 0xe0
      12'h9AE: dout <= 8'b11100000; // 2478 : 224 - 0xe0
      12'h9AF: dout <= 8'b11110000; // 2479 : 240 - 0xf0
      12'h9B0: dout <= 8'b11110000; // 2480 : 240 - 0xf0 -- Background 0x9b
      12'h9B1: dout <= 8'b11100000; // 2481 : 224 - 0xe0
      12'h9B2: dout <= 8'b11110000; // 2482 : 240 - 0xf0
      12'h9B3: dout <= 8'b11100000; // 2483 : 224 - 0xe0
      12'h9B4: dout <= 8'b10000000; // 2484 : 128 - 0x80
      12'h9B5: dout <= 8'b00001000; // 2485 :   8 - 0x8
      12'h9B6: dout <= 8'b00000100; // 2486 :   4 - 0x4
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b11111111; // 2488 : 255 - 0xff -- plane 1
      12'h9B9: dout <= 8'b11111111; // 2489 : 255 - 0xff
      12'h9BA: dout <= 8'b11111100; // 2490 : 252 - 0xfc
      12'h9BB: dout <= 8'b11111100; // 2491 : 252 - 0xfc
      12'h9BC: dout <= 8'b11111110; // 2492 : 254 - 0xfe
      12'h9BD: dout <= 8'b01111110; // 2493 : 126 - 0x7e
      12'h9BE: dout <= 8'b00111111; // 2494 :  63 - 0x3f
      12'h9BF: dout <= 8'b00001100; // 2495 :  12 - 0xc
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x9c
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000001; // 2498 :   1 - 0x1
      12'h9C3: dout <= 8'b00000011; // 2499 :   3 - 0x3
      12'h9C4: dout <= 8'b00000011; // 2500 :   3 - 0x3
      12'h9C5: dout <= 8'b00000011; // 2501 :   3 - 0x3
      12'h9C6: dout <= 8'b00000111; // 2502 :   7 - 0x7
      12'h9C7: dout <= 8'b00000111; // 2503 :   7 - 0x7
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout <= 8'b00000001; // 2505 :   1 - 0x1
      12'h9CA: dout <= 8'b00000011; // 2506 :   3 - 0x3
      12'h9CB: dout <= 8'b00000111; // 2507 :   7 - 0x7
      12'h9CC: dout <= 8'b00000111; // 2508 :   7 - 0x7
      12'h9CD: dout <= 8'b00000111; // 2509 :   7 - 0x7
      12'h9CE: dout <= 8'b00001111; // 2510 :  15 - 0xf
      12'h9CF: dout <= 8'b00001111; // 2511 :  15 - 0xf
      12'h9D0: dout <= 8'b00000111; // 2512 :   7 - 0x7 -- Background 0x9d
      12'h9D1: dout <= 8'b00000011; // 2513 :   3 - 0x3
      12'h9D2: dout <= 8'b00000011; // 2514 :   3 - 0x3
      12'h9D3: dout <= 8'b00000011; // 2515 :   3 - 0x3
      12'h9D4: dout <= 8'b00000011; // 2516 :   3 - 0x3
      12'h9D5: dout <= 8'b00000011; // 2517 :   3 - 0x3
      12'h9D6: dout <= 8'b00000011; // 2518 :   3 - 0x3
      12'h9D7: dout <= 8'b00000001; // 2519 :   1 - 0x1
      12'h9D8: dout <= 8'b00001111; // 2520 :  15 - 0xf -- plane 1
      12'h9D9: dout <= 8'b00001111; // 2521 :  15 - 0xf
      12'h9DA: dout <= 8'b00000111; // 2522 :   7 - 0x7
      12'h9DB: dout <= 8'b00000111; // 2523 :   7 - 0x7
      12'h9DC: dout <= 8'b00000111; // 2524 :   7 - 0x7
      12'h9DD: dout <= 8'b00000011; // 2525 :   3 - 0x3
      12'h9DE: dout <= 8'b00000011; // 2526 :   3 - 0x3
      12'h9DF: dout <= 8'b00000001; // 2527 :   1 - 0x1
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x9e
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000001; // 2533 :   1 - 0x1
      12'h9E6: dout <= 8'b00000010; // 2534 :   2 - 0x2
      12'h9E7: dout <= 8'b00000100; // 2535 :   4 - 0x4
      12'h9E8: dout <= 8'b00000001; // 2536 :   1 - 0x1 -- plane 1
      12'h9E9: dout <= 8'b00000001; // 2537 :   1 - 0x1
      12'h9EA: dout <= 8'b00000001; // 2538 :   1 - 0x1
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000011; // 2541 :   3 - 0x3
      12'h9EE: dout <= 8'b00000111; // 2542 :   7 - 0x7
      12'h9EF: dout <= 8'b00001111; // 2543 :  15 - 0xf
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x9f
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00011100; // 2550 :  28 - 0x1c
      12'h9F7: dout <= 8'b00111011; // 2551 :  59 - 0x3b
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000001; // 2556 :   1 - 0x1
      12'h9FD: dout <= 8'b00000011; // 2557 :   3 - 0x3
      12'h9FE: dout <= 8'b00111111; // 2558 :  63 - 0x3f
      12'h9FF: dout <= 8'b01111111; // 2559 : 127 - 0x7f
      12'hA00: dout <= 8'b01111110; // 2560 : 126 - 0x7e -- Background 0xa0
      12'hA01: dout <= 8'b11111110; // 2561 : 254 - 0xfe
      12'hA02: dout <= 8'b11111111; // 2562 : 255 - 0xff
      12'hA03: dout <= 8'b11111111; // 2563 : 255 - 0xff
      12'hA04: dout <= 8'b11111111; // 2564 : 255 - 0xff
      12'hA05: dout <= 8'b11111111; // 2565 : 255 - 0xff
      12'hA06: dout <= 8'b11111101; // 2566 : 253 - 0xfd
      12'hA07: dout <= 8'b11111001; // 2567 : 249 - 0xf9
      12'hA08: dout <= 8'b11111111; // 2568 : 255 - 0xff -- plane 1
      12'hA09: dout <= 8'b11111111; // 2569 : 255 - 0xff
      12'hA0A: dout <= 8'b11111111; // 2570 : 255 - 0xff
      12'hA0B: dout <= 8'b11111111; // 2571 : 255 - 0xff
      12'hA0C: dout <= 8'b11111111; // 2572 : 255 - 0xff
      12'hA0D: dout <= 8'b11111111; // 2573 : 255 - 0xff
      12'hA0E: dout <= 8'b11111101; // 2574 : 253 - 0xfd
      12'hA0F: dout <= 8'b11111001; // 2575 : 249 - 0xf9
      12'hA10: dout <= 8'b11110011; // 2576 : 243 - 0xf3 -- Background 0xa1
      12'hA11: dout <= 8'b11110111; // 2577 : 247 - 0xf7
      12'hA12: dout <= 8'b11110110; // 2578 : 246 - 0xf6
      12'hA13: dout <= 8'b11101110; // 2579 : 238 - 0xee
      12'hA14: dout <= 8'b11111101; // 2580 : 253 - 0xfd
      12'hA15: dout <= 8'b11111100; // 2581 : 252 - 0xfc
      12'hA16: dout <= 8'b11111000; // 2582 : 248 - 0xf8
      12'hA17: dout <= 8'b11100001; // 2583 : 225 - 0xe1
      12'hA18: dout <= 8'b11110011; // 2584 : 243 - 0xf3 -- plane 1
      12'hA19: dout <= 8'b11111111; // 2585 : 255 - 0xff
      12'hA1A: dout <= 8'b11111111; // 2586 : 255 - 0xff
      12'hA1B: dout <= 8'b11111111; // 2587 : 255 - 0xff
      12'hA1C: dout <= 8'b11111111; // 2588 : 255 - 0xff
      12'hA1D: dout <= 8'b11111111; // 2589 : 255 - 0xff
      12'hA1E: dout <= 8'b11111111; // 2590 : 255 - 0xff
      12'hA1F: dout <= 8'b11111111; // 2591 : 255 - 0xff
      12'hA20: dout <= 8'b11010011; // 2592 : 211 - 0xd3 -- Background 0xa2
      12'hA21: dout <= 8'b11001011; // 2593 : 203 - 0xcb
      12'hA22: dout <= 8'b11000011; // 2594 : 195 - 0xc3
      12'hA23: dout <= 8'b11100001; // 2595 : 225 - 0xe1
      12'hA24: dout <= 8'b11111001; // 2596 : 249 - 0xf9
      12'hA25: dout <= 8'b00111001; // 2597 :  57 - 0x39
      12'hA26: dout <= 8'b01000010; // 2598 :  66 - 0x42
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b11111111; // 2600 : 255 - 0xff -- plane 1
      12'hA29: dout <= 8'b11111111; // 2601 : 255 - 0xff
      12'hA2A: dout <= 8'b11111111; // 2602 : 255 - 0xff
      12'hA2B: dout <= 8'b11111111; // 2603 : 255 - 0xff
      12'hA2C: dout <= 8'b11111111; // 2604 : 255 - 0xff
      12'hA2D: dout <= 8'b11111111; // 2605 : 255 - 0xff
      12'hA2E: dout <= 8'b11111111; // 2606 : 255 - 0xff
      12'hA2F: dout <= 8'b11111111; // 2607 : 255 - 0xff
      12'hA30: dout <= 8'b00000111; // 2608 :   7 - 0x7 -- Background 0xa3
      12'hA31: dout <= 8'b00001111; // 2609 :  15 - 0xf
      12'hA32: dout <= 8'b00011001; // 2610 :  25 - 0x19
      12'hA33: dout <= 8'b00110000; // 2611 :  48 - 0x30
      12'hA34: dout <= 8'b01100011; // 2612 :  99 - 0x63
      12'hA35: dout <= 8'b01110010; // 2613 : 114 - 0x72
      12'hA36: dout <= 8'b01110000; // 2614 : 112 - 0x70
      12'hA37: dout <= 8'b00000001; // 2615 :   1 - 0x1
      12'hA38: dout <= 8'b00000111; // 2616 :   7 - 0x7 -- plane 1
      12'hA39: dout <= 8'b00001111; // 2617 :  15 - 0xf
      12'hA3A: dout <= 8'b00011111; // 2618 :  31 - 0x1f
      12'hA3B: dout <= 8'b00111111; // 2619 :  63 - 0x3f
      12'hA3C: dout <= 8'b11111100; // 2620 : 252 - 0xfc
      12'hA3D: dout <= 8'b11111100; // 2621 : 252 - 0xfc
      12'hA3E: dout <= 8'b11111111; // 2622 : 255 - 0xff
      12'hA3F: dout <= 8'b11111111; // 2623 : 255 - 0xff
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0xa4
      12'hA41: dout <= 8'b00011111; // 2625 :  31 - 0x1f
      12'hA42: dout <= 8'b00100000; // 2626 :  32 - 0x20
      12'hA43: dout <= 8'b11000000; // 2627 : 192 - 0xc0
      12'hA44: dout <= 8'b11000000; // 2628 : 192 - 0xc0
      12'hA45: dout <= 8'b11110000; // 2629 : 240 - 0xf0
      12'hA46: dout <= 8'b11111111; // 2630 : 255 - 0xff
      12'hA47: dout <= 8'b11111111; // 2631 : 255 - 0xff
      12'hA48: dout <= 8'b11111111; // 2632 : 255 - 0xff -- plane 1
      12'hA49: dout <= 8'b11111111; // 2633 : 255 - 0xff
      12'hA4A: dout <= 8'b11111111; // 2634 : 255 - 0xff
      12'hA4B: dout <= 8'b11111111; // 2635 : 255 - 0xff
      12'hA4C: dout <= 8'b11111111; // 2636 : 255 - 0xff
      12'hA4D: dout <= 8'b11111111; // 2637 : 255 - 0xff
      12'hA4E: dout <= 8'b11111111; // 2638 : 255 - 0xff
      12'hA4F: dout <= 8'b11111111; // 2639 : 255 - 0xff
      12'hA50: dout <= 8'b10101011; // 2640 : 171 - 0xab -- Background 0xa5
      12'hA51: dout <= 8'b11000001; // 2641 : 193 - 0xc1
      12'hA52: dout <= 8'b10000001; // 2642 : 129 - 0x81
      12'hA53: dout <= 8'b10010001; // 2643 : 145 - 0x91
      12'hA54: dout <= 8'b10000010; // 2644 : 130 - 0x82
      12'hA55: dout <= 8'b11111100; // 2645 : 252 - 0xfc
      12'hA56: dout <= 8'b11100000; // 2646 : 224 - 0xe0
      12'hA57: dout <= 8'b11001110; // 2647 : 206 - 0xce
      12'hA58: dout <= 8'b11111111; // 2648 : 255 - 0xff -- plane 1
      12'hA59: dout <= 8'b11111111; // 2649 : 255 - 0xff
      12'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      12'hA5B: dout <= 8'b11111111; // 2651 : 255 - 0xff
      12'hA5C: dout <= 8'b11111111; // 2652 : 255 - 0xff
      12'hA5D: dout <= 8'b11111111; // 2653 : 255 - 0xff
      12'hA5E: dout <= 8'b11111111; // 2654 : 255 - 0xff
      12'hA5F: dout <= 8'b11111111; // 2655 : 255 - 0xff
      12'hA60: dout <= 8'b11100101; // 2656 : 229 - 0xe5 -- Background 0xa6
      12'hA61: dout <= 8'b11011010; // 2657 : 218 - 0xda
      12'hA62: dout <= 8'b11110000; // 2658 : 240 - 0xf0
      12'hA63: dout <= 8'b11100000; // 2659 : 224 - 0xe0
      12'hA64: dout <= 8'b11000000; // 2660 : 192 - 0xc0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b11111111; // 2664 : 255 - 0xff -- plane 1
      12'hA69: dout <= 8'b11111111; // 2665 : 255 - 0xff
      12'hA6A: dout <= 8'b11110000; // 2666 : 240 - 0xf0
      12'hA6B: dout <= 8'b11100000; // 2667 : 224 - 0xe0
      12'hA6C: dout <= 8'b11000000; // 2668 : 192 - 0xc0
      12'hA6D: dout <= 8'b10000000; // 2669 : 128 - 0x80
      12'hA6E: dout <= 8'b10000000; // 2670 : 128 - 0x80
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b11110000; // 2672 : 240 - 0xf0 -- Background 0xa7
      12'hA71: dout <= 8'b11111000; // 2673 : 248 - 0xf8
      12'hA72: dout <= 8'b11001100; // 2674 : 204 - 0xcc
      12'hA73: dout <= 8'b10000110; // 2675 : 134 - 0x86
      12'hA74: dout <= 8'b01100010; // 2676 :  98 - 0x62
      12'hA75: dout <= 8'b00100110; // 2677 :  38 - 0x26
      12'hA76: dout <= 8'b00000110; // 2678 :   6 - 0x6
      12'hA77: dout <= 8'b11000000; // 2679 : 192 - 0xc0
      12'hA78: dout <= 8'b11110000; // 2680 : 240 - 0xf0 -- plane 1
      12'hA79: dout <= 8'b11111000; // 2681 : 248 - 0xf8
      12'hA7A: dout <= 8'b11111100; // 2682 : 252 - 0xfc
      12'hA7B: dout <= 8'b11111110; // 2683 : 254 - 0xfe
      12'hA7C: dout <= 8'b10011111; // 2684 : 159 - 0x9f
      12'hA7D: dout <= 8'b10011111; // 2685 : 159 - 0x9f
      12'hA7E: dout <= 8'b11111111; // 2686 : 255 - 0xff
      12'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Background 0xa8
      12'hA81: dout <= 8'b11111100; // 2689 : 252 - 0xfc
      12'hA82: dout <= 8'b00000110; // 2690 :   6 - 0x6
      12'hA83: dout <= 8'b00000011; // 2691 :   3 - 0x3
      12'hA84: dout <= 8'b00000001; // 2692 :   1 - 0x1
      12'hA85: dout <= 8'b00000111; // 2693 :   7 - 0x7
      12'hA86: dout <= 8'b11111111; // 2694 : 255 - 0xff
      12'hA87: dout <= 8'b11111111; // 2695 : 255 - 0xff
      12'hA88: dout <= 8'b11111111; // 2696 : 255 - 0xff -- plane 1
      12'hA89: dout <= 8'b11111111; // 2697 : 255 - 0xff
      12'hA8A: dout <= 8'b11111111; // 2698 : 255 - 0xff
      12'hA8B: dout <= 8'b11111111; // 2699 : 255 - 0xff
      12'hA8C: dout <= 8'b11111111; // 2700 : 255 - 0xff
      12'hA8D: dout <= 8'b11111111; // 2701 : 255 - 0xff
      12'hA8E: dout <= 8'b11111111; // 2702 : 255 - 0xff
      12'hA8F: dout <= 8'b11111111; // 2703 : 255 - 0xff
      12'hA90: dout <= 8'b11010101; // 2704 : 213 - 0xd5 -- Background 0xa9
      12'hA91: dout <= 8'b10000011; // 2705 : 131 - 0x83
      12'hA92: dout <= 8'b10000001; // 2706 : 129 - 0x81
      12'hA93: dout <= 8'b10001001; // 2707 : 137 - 0x89
      12'hA94: dout <= 8'b01000001; // 2708 :  65 - 0x41
      12'hA95: dout <= 8'b00111111; // 2709 :  63 - 0x3f
      12'hA96: dout <= 8'b00000111; // 2710 :   7 - 0x7
      12'hA97: dout <= 8'b11010011; // 2711 : 211 - 0xd3
      12'hA98: dout <= 8'b11111111; // 2712 : 255 - 0xff -- plane 1
      12'hA99: dout <= 8'b11111111; // 2713 : 255 - 0xff
      12'hA9A: dout <= 8'b11111111; // 2714 : 255 - 0xff
      12'hA9B: dout <= 8'b11111111; // 2715 : 255 - 0xff
      12'hA9C: dout <= 8'b11111111; // 2716 : 255 - 0xff
      12'hA9D: dout <= 8'b11111111; // 2717 : 255 - 0xff
      12'hA9E: dout <= 8'b11111111; // 2718 : 255 - 0xff
      12'hA9F: dout <= 8'b11111111; // 2719 : 255 - 0xff
      12'hAA0: dout <= 8'b01101111; // 2720 : 111 - 0x6f -- Background 0xaa
      12'hAA1: dout <= 8'b11011011; // 2721 : 219 - 0xdb
      12'hAA2: dout <= 8'b00001111; // 2722 :  15 - 0xf
      12'hAA3: dout <= 8'b00000111; // 2723 :   7 - 0x7
      12'hAA4: dout <= 8'b00000011; // 2724 :   3 - 0x3
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b11111111; // 2728 : 255 - 0xff -- plane 1
      12'hAA9: dout <= 8'b11111111; // 2729 : 255 - 0xff
      12'hAAA: dout <= 8'b00001111; // 2730 :  15 - 0xf
      12'hAAB: dout <= 8'b00000111; // 2731 :   7 - 0x7
      12'hAAC: dout <= 8'b00000011; // 2732 :   3 - 0x3
      12'hAAD: dout <= 8'b00000001; // 2733 :   1 - 0x1
      12'hAAE: dout <= 8'b00000001; // 2734 :   1 - 0x1
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b00000000; // 2736 :   0 - 0x0 -- Background 0xab
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout <= 8'b00111000; // 2742 :  56 - 0x38
      12'hAB7: dout <= 8'b11011100; // 2743 : 220 - 0xdc
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b10000000; // 2748 : 128 - 0x80
      12'hABD: dout <= 8'b11000000; // 2749 : 192 - 0xc0
      12'hABE: dout <= 8'b11111100; // 2750 : 252 - 0xfc
      12'hABF: dout <= 8'b11111110; // 2751 : 254 - 0xfe
      12'hAC0: dout <= 8'b01111110; // 2752 : 126 - 0x7e -- Background 0xac
      12'hAC1: dout <= 8'b01111111; // 2753 : 127 - 0x7f
      12'hAC2: dout <= 8'b01111111; // 2754 : 127 - 0x7f
      12'hAC3: dout <= 8'b11111111; // 2755 : 255 - 0xff
      12'hAC4: dout <= 8'b11111111; // 2756 : 255 - 0xff
      12'hAC5: dout <= 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout <= 8'b10111111; // 2758 : 191 - 0xbf
      12'hAC7: dout <= 8'b10011111; // 2759 : 159 - 0x9f
      12'hAC8: dout <= 8'b11111111; // 2760 : 255 - 0xff -- plane 1
      12'hAC9: dout <= 8'b11111111; // 2761 : 255 - 0xff
      12'hACA: dout <= 8'b11111111; // 2762 : 255 - 0xff
      12'hACB: dout <= 8'b11111111; // 2763 : 255 - 0xff
      12'hACC: dout <= 8'b11111111; // 2764 : 255 - 0xff
      12'hACD: dout <= 8'b11111111; // 2765 : 255 - 0xff
      12'hACE: dout <= 8'b10111111; // 2766 : 191 - 0xbf
      12'hACF: dout <= 8'b10011111; // 2767 : 159 - 0x9f
      12'hAD0: dout <= 8'b11001111; // 2768 : 207 - 0xcf -- Background 0xad
      12'hAD1: dout <= 8'b11101111; // 2769 : 239 - 0xef
      12'hAD2: dout <= 8'b01101111; // 2770 : 111 - 0x6f
      12'hAD3: dout <= 8'b01110111; // 2771 : 119 - 0x77
      12'hAD4: dout <= 8'b10111111; // 2772 : 191 - 0xbf
      12'hAD5: dout <= 8'b00111111; // 2773 :  63 - 0x3f
      12'hAD6: dout <= 8'b00011111; // 2774 :  31 - 0x1f
      12'hAD7: dout <= 8'b10000111; // 2775 : 135 - 0x87
      12'hAD8: dout <= 8'b11001111; // 2776 : 207 - 0xcf -- plane 1
      12'hAD9: dout <= 8'b11111111; // 2777 : 255 - 0xff
      12'hADA: dout <= 8'b11111111; // 2778 : 255 - 0xff
      12'hADB: dout <= 8'b11111111; // 2779 : 255 - 0xff
      12'hADC: dout <= 8'b11111111; // 2780 : 255 - 0xff
      12'hADD: dout <= 8'b11111111; // 2781 : 255 - 0xff
      12'hADE: dout <= 8'b11111111; // 2782 : 255 - 0xff
      12'hADF: dout <= 8'b11111111; // 2783 : 255 - 0xff
      12'hAE0: dout <= 8'b11001011; // 2784 : 203 - 0xcb -- Background 0xae
      12'hAE1: dout <= 8'b11010011; // 2785 : 211 - 0xd3
      12'hAE2: dout <= 8'b11000011; // 2786 : 195 - 0xc3
      12'hAE3: dout <= 8'b10000111; // 2787 : 135 - 0x87
      12'hAE4: dout <= 8'b10011111; // 2788 : 159 - 0x9f
      12'hAE5: dout <= 8'b10011100; // 2789 : 156 - 0x9c
      12'hAE6: dout <= 8'b01000010; // 2790 :  66 - 0x42
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b11111111; // 2792 : 255 - 0xff -- plane 1
      12'hAE9: dout <= 8'b11111111; // 2793 : 255 - 0xff
      12'hAEA: dout <= 8'b11111111; // 2794 : 255 - 0xff
      12'hAEB: dout <= 8'b11111111; // 2795 : 255 - 0xff
      12'hAEC: dout <= 8'b11111111; // 2796 : 255 - 0xff
      12'hAED: dout <= 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout <= 8'b11111111; // 2798 : 255 - 0xff
      12'hAEF: dout <= 8'b11111111; // 2799 : 255 - 0xff
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0xaf
      12'hAF1: dout <= 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout <= 8'b10000000; // 2802 : 128 - 0x80
      12'hAF3: dout <= 8'b11000000; // 2803 : 192 - 0xc0
      12'hAF4: dout <= 8'b11000000; // 2804 : 192 - 0xc0
      12'hAF5: dout <= 8'b11000000; // 2805 : 192 - 0xc0
      12'hAF6: dout <= 8'b11100000; // 2806 : 224 - 0xe0
      12'hAF7: dout <= 8'b11100000; // 2807 : 224 - 0xe0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout <= 8'b10000000; // 2809 : 128 - 0x80
      12'hAFA: dout <= 8'b11000000; // 2810 : 192 - 0xc0
      12'hAFB: dout <= 8'b11100000; // 2811 : 224 - 0xe0
      12'hAFC: dout <= 8'b11100000; // 2812 : 224 - 0xe0
      12'hAFD: dout <= 8'b11100000; // 2813 : 224 - 0xe0
      12'hAFE: dout <= 8'b11110000; // 2814 : 240 - 0xf0
      12'hAFF: dout <= 8'b11110000; // 2815 : 240 - 0xf0
      12'hB00: dout <= 8'b11100000; // 2816 : 224 - 0xe0 -- Background 0xb0
      12'hB01: dout <= 8'b11000000; // 2817 : 192 - 0xc0
      12'hB02: dout <= 8'b11000000; // 2818 : 192 - 0xc0
      12'hB03: dout <= 8'b11000000; // 2819 : 192 - 0xc0
      12'hB04: dout <= 8'b11000000; // 2820 : 192 - 0xc0
      12'hB05: dout <= 8'b11000000; // 2821 : 192 - 0xc0
      12'hB06: dout <= 8'b11000000; // 2822 : 192 - 0xc0
      12'hB07: dout <= 8'b10000000; // 2823 : 128 - 0x80
      12'hB08: dout <= 8'b11110000; // 2824 : 240 - 0xf0 -- plane 1
      12'hB09: dout <= 8'b11110000; // 2825 : 240 - 0xf0
      12'hB0A: dout <= 8'b11100000; // 2826 : 224 - 0xe0
      12'hB0B: dout <= 8'b11100000; // 2827 : 224 - 0xe0
      12'hB0C: dout <= 8'b11100000; // 2828 : 224 - 0xe0
      12'hB0D: dout <= 8'b11000000; // 2829 : 192 - 0xc0
      12'hB0E: dout <= 8'b11000000; // 2830 : 192 - 0xc0
      12'hB0F: dout <= 8'b10000000; // 2831 : 128 - 0x80
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Background 0xb1
      12'hB11: dout <= 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout <= 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout <= 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout <= 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout <= 8'b10000000; // 2837 : 128 - 0x80
      12'hB16: dout <= 8'b01000000; // 2838 :  64 - 0x40
      12'hB17: dout <= 8'b00100000; // 2839 :  32 - 0x20
      12'hB18: dout <= 8'b10000000; // 2840 : 128 - 0x80 -- plane 1
      12'hB19: dout <= 8'b10000000; // 2841 : 128 - 0x80
      12'hB1A: dout <= 8'b10000000; // 2842 : 128 - 0x80
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b11000000; // 2845 : 192 - 0xc0
      12'hB1E: dout <= 8'b11100000; // 2846 : 224 - 0xe0
      12'hB1F: dout <= 8'b11110000; // 2847 : 240 - 0xf0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0xb2
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000001; // 2851 :   1 - 0x1
      12'hB24: dout <= 8'b00000011; // 2852 :   3 - 0x3
      12'hB25: dout <= 8'b00000111; // 2853 :   7 - 0x7
      12'hB26: dout <= 8'b00000111; // 2854 :   7 - 0x7
      12'hB27: dout <= 8'b00000111; // 2855 :   7 - 0x7
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- plane 1
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000001; // 2858 :   1 - 0x1
      12'hB2B: dout <= 8'b00000011; // 2859 :   3 - 0x3
      12'hB2C: dout <= 8'b00000111; // 2860 :   7 - 0x7
      12'hB2D: dout <= 8'b00000111; // 2861 :   7 - 0x7
      12'hB2E: dout <= 8'b00000111; // 2862 :   7 - 0x7
      12'hB2F: dout <= 8'b00000111; // 2863 :   7 - 0x7
      12'hB30: dout <= 8'b00000011; // 2864 :   3 - 0x3 -- Background 0xb3
      12'hB31: dout <= 8'b00000001; // 2865 :   1 - 0x1
      12'hB32: dout <= 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout <= 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout <= 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout <= 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout <= 8'b00000001; // 2870 :   1 - 0x1
      12'hB37: dout <= 8'b00000001; // 2871 :   1 - 0x1
      12'hB38: dout <= 8'b00000011; // 2872 :   3 - 0x3 -- plane 1
      12'hB39: dout <= 8'b00000001; // 2873 :   1 - 0x1
      12'hB3A: dout <= 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout <= 8'b00000000; // 2875 :   0 - 0x0
      12'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout <= 8'b00000001; // 2877 :   1 - 0x1
      12'hB3E: dout <= 8'b00000011; // 2878 :   3 - 0x3
      12'hB3F: dout <= 8'b00000011; // 2879 :   3 - 0x3
      12'hB40: dout <= 8'b00000001; // 2880 :   1 - 0x1 -- Background 0xb4
      12'hB41: dout <= 8'b00000001; // 2881 :   1 - 0x1
      12'hB42: dout <= 8'b00000111; // 2882 :   7 - 0x7
      12'hB43: dout <= 8'b00000011; // 2883 :   3 - 0x3
      12'hB44: dout <= 8'b00000100; // 2884 :   4 - 0x4
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000011; // 2888 :   3 - 0x3 -- plane 1
      12'hB49: dout <= 8'b00000011; // 2889 :   3 - 0x3
      12'hB4A: dout <= 8'b00000111; // 2890 :   7 - 0x7
      12'hB4B: dout <= 8'b00011111; // 2891 :  31 - 0x1f
      12'hB4C: dout <= 8'b00111111; // 2892 :  63 - 0x3f
      12'hB4D: dout <= 8'b00111111; // 2893 :  63 - 0x3f
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0xb5
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000111; // 2903 :   7 - 0x7
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- plane 1
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000001; // 2908 :   1 - 0x1
      12'hB5D: dout <= 8'b00000011; // 2909 :   3 - 0x3
      12'hB5E: dout <= 8'b00000011; // 2910 :   3 - 0x3
      12'hB5F: dout <= 8'b00001111; // 2911 :  15 - 0xf
      12'hB60: dout <= 8'b00001110; // 2912 :  14 - 0xe -- Background 0xb6
      12'hB61: dout <= 8'b00111110; // 2913 :  62 - 0x3e
      12'hB62: dout <= 8'b01111111; // 2914 : 127 - 0x7f
      12'hB63: dout <= 8'b11111111; // 2915 : 255 - 0xff
      12'hB64: dout <= 8'b11111111; // 2916 : 255 - 0xff
      12'hB65: dout <= 8'b11101111; // 2917 : 239 - 0xef
      12'hB66: dout <= 8'b11110111; // 2918 : 247 - 0xf7
      12'hB67: dout <= 8'b11111000; // 2919 : 248 - 0xf8
      12'hB68: dout <= 8'b00111111; // 2920 :  63 - 0x3f -- plane 1
      12'hB69: dout <= 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout <= 8'b11111111; // 2922 : 255 - 0xff
      12'hB6B: dout <= 8'b11111111; // 2923 : 255 - 0xff
      12'hB6C: dout <= 8'b11111111; // 2924 : 255 - 0xff
      12'hB6D: dout <= 8'b11111111; // 2925 : 255 - 0xff
      12'hB6E: dout <= 8'b11111111; // 2926 : 255 - 0xff
      12'hB6F: dout <= 8'b11111111; // 2927 : 255 - 0xff
      12'hB70: dout <= 8'b11111111; // 2928 : 255 - 0xff -- Background 0xb7
      12'hB71: dout <= 8'b11111111; // 2929 : 255 - 0xff
      12'hB72: dout <= 8'b11111111; // 2930 : 255 - 0xff
      12'hB73: dout <= 8'b00011111; // 2931 :  31 - 0x1f
      12'hB74: dout <= 8'b00011111; // 2932 :  31 - 0x1f
      12'hB75: dout <= 8'b01111111; // 2933 : 127 - 0x7f
      12'hB76: dout <= 8'b11111111; // 2934 : 255 - 0xff
      12'hB77: dout <= 8'b11111110; // 2935 : 254 - 0xfe
      12'hB78: dout <= 8'b11111111; // 2936 : 255 - 0xff -- plane 1
      12'hB79: dout <= 8'b11111111; // 2937 : 255 - 0xff
      12'hB7A: dout <= 8'b11111111; // 2938 : 255 - 0xff
      12'hB7B: dout <= 8'b00011111; // 2939 :  31 - 0x1f
      12'hB7C: dout <= 8'b01111111; // 2940 : 127 - 0x7f
      12'hB7D: dout <= 8'b11111111; // 2941 : 255 - 0xff
      12'hB7E: dout <= 8'b11111111; // 2942 : 255 - 0xff
      12'hB7F: dout <= 8'b11111111; // 2943 : 255 - 0xff
      12'hB80: dout <= 8'b11111111; // 2944 : 255 - 0xff -- Background 0xb8
      12'hB81: dout <= 8'b11111111; // 2945 : 255 - 0xff
      12'hB82: dout <= 8'b11111111; // 2946 : 255 - 0xff
      12'hB83: dout <= 8'b11111100; // 2947 : 252 - 0xfc
      12'hB84: dout <= 8'b11111000; // 2948 : 248 - 0xf8
      12'hB85: dout <= 8'b10000000; // 2949 : 128 - 0x80
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b11111111; // 2952 : 255 - 0xff -- plane 1
      12'hB89: dout <= 8'b11111111; // 2953 : 255 - 0xff
      12'hB8A: dout <= 8'b11111111; // 2954 : 255 - 0xff
      12'hB8B: dout <= 8'b11111100; // 2955 : 252 - 0xfc
      12'hB8C: dout <= 8'b11111000; // 2956 : 248 - 0xf8
      12'hB8D: dout <= 8'b11111000; // 2957 : 248 - 0xf8
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00110000; // 2960 :  48 - 0x30 -- Background 0xb9
      12'hB91: dout <= 8'b01111111; // 2961 : 127 - 0x7f
      12'hB92: dout <= 8'b01111111; // 2962 : 127 - 0x7f
      12'hB93: dout <= 8'b00111111; // 2963 :  63 - 0x3f
      12'hB94: dout <= 8'b10000111; // 2964 : 135 - 0x87
      12'hB95: dout <= 8'b11110000; // 2965 : 240 - 0xf0
      12'hB96: dout <= 8'b11111111; // 2966 : 255 - 0xff
      12'hB97: dout <= 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout <= 8'b11001111; // 2968 : 207 - 0xcf -- plane 1
      12'hB99: dout <= 8'b10001000; // 2969 : 136 - 0x88
      12'hB9A: dout <= 8'b11011101; // 2970 : 221 - 0xdd
      12'hB9B: dout <= 8'b11001000; // 2971 : 200 - 0xc8
      12'hB9C: dout <= 8'b11111000; // 2972 : 248 - 0xf8
      12'hB9D: dout <= 8'b11111111; // 2973 : 255 - 0xff
      12'hB9E: dout <= 8'b11111111; // 2974 : 255 - 0xff
      12'hB9F: dout <= 8'b11111111; // 2975 : 255 - 0xff
      12'hBA0: dout <= 8'b11100101; // 2976 : 229 - 0xe5 -- Background 0xba
      12'hBA1: dout <= 8'b11011010; // 2977 : 218 - 0xda
      12'hBA2: dout <= 8'b11000000; // 2978 : 192 - 0xc0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b11111111; // 2984 : 255 - 0xff -- plane 1
      12'hBA9: dout <= 8'b11111111; // 2985 : 255 - 0xff
      12'hBAA: dout <= 8'b11000000; // 2986 : 192 - 0xc0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000110; // 2992 :   6 - 0x6 -- Background 0xbb
      12'hBB1: dout <= 8'b11111111; // 2993 : 255 - 0xff
      12'hBB2: dout <= 8'b11111111; // 2994 : 255 - 0xff
      12'hBB3: dout <= 8'b11111110; // 2995 : 254 - 0xfe
      12'hBB4: dout <= 8'b11110001; // 2996 : 241 - 0xf1
      12'hBB5: dout <= 8'b00000111; // 2997 :   7 - 0x7
      12'hBB6: dout <= 8'b11111111; // 2998 : 255 - 0xff
      12'hBB7: dout <= 8'b11111111; // 2999 : 255 - 0xff
      12'hBB8: dout <= 8'b11111001; // 3000 : 249 - 0xf9 -- plane 1
      12'hBB9: dout <= 8'b10001000; // 3001 : 136 - 0x88
      12'hBBA: dout <= 8'b11011101; // 3002 : 221 - 0xdd
      12'hBBB: dout <= 8'b10001001; // 3003 : 137 - 0x89
      12'hBBC: dout <= 8'b00001111; // 3004 :  15 - 0xf
      12'hBBD: dout <= 8'b11111111; // 3005 : 255 - 0xff
      12'hBBE: dout <= 8'b11111111; // 3006 : 255 - 0xff
      12'hBBF: dout <= 8'b11111111; // 3007 : 255 - 0xff
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0xbc
      12'hBC1: dout <= 8'b00000001; // 3009 :   1 - 0x1
      12'hBC2: dout <= 8'b00000010; // 3010 :   2 - 0x2
      12'hBC3: dout <= 8'b00000111; // 3011 :   7 - 0x7
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00100000; // 3014 :  32 - 0x20
      12'hBC7: dout <= 8'b11111111; // 3015 : 255 - 0xff
      12'hBC8: dout <= 8'b00000011; // 3016 :   3 - 0x3 -- plane 1
      12'hBC9: dout <= 8'b00000111; // 3017 :   7 - 0x7
      12'hBCA: dout <= 8'b00001111; // 3018 :  15 - 0xf
      12'hBCB: dout <= 8'b00000111; // 3019 :   7 - 0x7
      12'hBCC: dout <= 8'b10000111; // 3020 : 135 - 0x87
      12'hBCD: dout <= 8'b11000011; // 3021 : 195 - 0xc3
      12'hBCE: dout <= 8'b11100000; // 3022 : 224 - 0xe0
      12'hBCF: dout <= 8'b11111111; // 3023 : 255 - 0xff
      12'hBD0: dout <= 8'b01111111; // 3024 : 127 - 0x7f -- Background 0xbd
      12'hBD1: dout <= 8'b01111111; // 3025 : 127 - 0x7f
      12'hBD2: dout <= 8'b01111111; // 3026 : 127 - 0x7f
      12'hBD3: dout <= 8'b11111111; // 3027 : 255 - 0xff
      12'hBD4: dout <= 8'b11111111; // 3028 : 255 - 0xff
      12'hBD5: dout <= 8'b11111111; // 3029 : 255 - 0xff
      12'hBD6: dout <= 8'b11111111; // 3030 : 255 - 0xff
      12'hBD7: dout <= 8'b11111110; // 3031 : 254 - 0xfe
      12'hBD8: dout <= 8'b11111111; // 3032 : 255 - 0xff -- plane 1
      12'hBD9: dout <= 8'b11111111; // 3033 : 255 - 0xff
      12'hBDA: dout <= 8'b11111111; // 3034 : 255 - 0xff
      12'hBDB: dout <= 8'b11111111; // 3035 : 255 - 0xff
      12'hBDC: dout <= 8'b11111111; // 3036 : 255 - 0xff
      12'hBDD: dout <= 8'b11111111; // 3037 : 255 - 0xff
      12'hBDE: dout <= 8'b11111111; // 3038 : 255 - 0xff
      12'hBDF: dout <= 8'b11111110; // 3039 : 254 - 0xfe
      12'hBE0: dout <= 8'b11111100; // 3040 : 252 - 0xfc -- Background 0xbe
      12'hBE1: dout <= 8'b10111000; // 3041 : 184 - 0xb8
      12'hBE2: dout <= 8'b01111000; // 3042 : 120 - 0x78
      12'hBE3: dout <= 8'b01111000; // 3043 : 120 - 0x78
      12'hBE4: dout <= 8'b10110000; // 3044 : 176 - 0xb0
      12'hBE5: dout <= 8'b01111000; // 3045 : 120 - 0x78
      12'hBE6: dout <= 8'b11111100; // 3046 : 252 - 0xfc
      12'hBE7: dout <= 8'b11111110; // 3047 : 254 - 0xfe
      12'hBE8: dout <= 8'b11111100; // 3048 : 252 - 0xfc -- plane 1
      12'hBE9: dout <= 8'b11111000; // 3049 : 248 - 0xf8
      12'hBEA: dout <= 8'b11111000; // 3050 : 248 - 0xf8
      12'hBEB: dout <= 8'b11111000; // 3051 : 248 - 0xf8
      12'hBEC: dout <= 8'b11111000; // 3052 : 248 - 0xf8
      12'hBED: dout <= 8'b11111100; // 3053 : 252 - 0xfc
      12'hBEE: dout <= 8'b11111110; // 3054 : 254 - 0xfe
      12'hBEF: dout <= 8'b11111111; // 3055 : 255 - 0xff
      12'hBF0: dout <= 8'b11111111; // 3056 : 255 - 0xff -- Background 0xbf
      12'hBF1: dout <= 8'b11111111; // 3057 : 255 - 0xff
      12'hBF2: dout <= 8'b11111111; // 3058 : 255 - 0xff
      12'hBF3: dout <= 8'b11111111; // 3059 : 255 - 0xff
      12'hBF4: dout <= 8'b11111111; // 3060 : 255 - 0xff
      12'hBF5: dout <= 8'b10011100; // 3061 : 156 - 0x9c
      12'hBF6: dout <= 8'b01000010; // 3062 :  66 - 0x42
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b11111111; // 3064 : 255 - 0xff -- plane 1
      12'hBF9: dout <= 8'b11111111; // 3065 : 255 - 0xff
      12'hBFA: dout <= 8'b11111111; // 3066 : 255 - 0xff
      12'hBFB: dout <= 8'b11111111; // 3067 : 255 - 0xff
      12'hBFC: dout <= 8'b11111111; // 3068 : 255 - 0xff
      12'hBFD: dout <= 8'b11111111; // 3069 : 255 - 0xff
      12'hBFE: dout <= 8'b11111111; // 3070 : 255 - 0xff
      12'hBFF: dout <= 8'b11111111; // 3071 : 255 - 0xff
      12'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Background 0xc0
      12'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      12'hC02: dout <= 8'b00100000; // 3074 :  32 - 0x20
      12'hC03: dout <= 8'b01000000; // 3075 :  64 - 0x40
      12'hC04: dout <= 8'b10001010; // 3076 : 138 - 0x8a
      12'hC05: dout <= 8'b00011110; // 3077 :  30 - 0x1e
      12'hC06: dout <= 8'b01111110; // 3078 : 126 - 0x7e
      12'hC07: dout <= 8'b10111110; // 3079 : 190 - 0xbe
      12'hC08: dout <= 8'b11000000; // 3080 : 192 - 0xc0 -- plane 1
      12'hC09: dout <= 8'b11110000; // 3081 : 240 - 0xf0
      12'hC0A: dout <= 8'b11111100; // 3082 : 252 - 0xfc
      12'hC0B: dout <= 8'b11111100; // 3083 : 252 - 0xfc
      12'hC0C: dout <= 8'b11111110; // 3084 : 254 - 0xfe
      12'hC0D: dout <= 8'b11111110; // 3085 : 254 - 0xfe
      12'hC0E: dout <= 8'b11111110; // 3086 : 254 - 0xfe
      12'hC0F: dout <= 8'b11111110; // 3087 : 254 - 0xfe
      12'hC10: dout <= 8'b11011111; // 3088 : 223 - 0xdf -- Background 0xc1
      12'hC11: dout <= 8'b11111111; // 3089 : 255 - 0xff
      12'hC12: dout <= 8'b11111110; // 3090 : 254 - 0xfe
      12'hC13: dout <= 8'b11111100; // 3091 : 252 - 0xfc
      12'hC14: dout <= 8'b11110000; // 3092 : 240 - 0xf0
      12'hC15: dout <= 8'b11100000; // 3093 : 224 - 0xe0
      12'hC16: dout <= 8'b10000000; // 3094 : 128 - 0x80
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b11111111; // 3096 : 255 - 0xff -- plane 1
      12'hC19: dout <= 8'b11111111; // 3097 : 255 - 0xff
      12'hC1A: dout <= 8'b11111110; // 3098 : 254 - 0xfe
      12'hC1B: dout <= 8'b11111100; // 3099 : 252 - 0xfc
      12'hC1C: dout <= 8'b11110000; // 3100 : 240 - 0xf0
      12'hC1D: dout <= 8'b11100000; // 3101 : 224 - 0xe0
      12'hC1E: dout <= 8'b10000000; // 3102 : 128 - 0x80
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Background 0xc2
      12'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout <= 8'b00000100; // 3106 :   4 - 0x4
      12'hC23: dout <= 8'b00000010; // 3107 :   2 - 0x2
      12'hC24: dout <= 8'b01010001; // 3108 :  81 - 0x51
      12'hC25: dout <= 8'b01111000; // 3109 : 120 - 0x78
      12'hC26: dout <= 8'b01111110; // 3110 : 126 - 0x7e
      12'hC27: dout <= 8'b11111101; // 3111 : 253 - 0xfd
      12'hC28: dout <= 8'b00000011; // 3112 :   3 - 0x3 -- plane 1
      12'hC29: dout <= 8'b00001111; // 3113 :  15 - 0xf
      12'hC2A: dout <= 8'b00111111; // 3114 :  63 - 0x3f
      12'hC2B: dout <= 8'b00111111; // 3115 :  63 - 0x3f
      12'hC2C: dout <= 8'b01111111; // 3116 : 127 - 0x7f
      12'hC2D: dout <= 8'b01111111; // 3117 : 127 - 0x7f
      12'hC2E: dout <= 8'b01111110; // 3118 : 126 - 0x7e
      12'hC2F: dout <= 8'b11111111; // 3119 : 255 - 0xff
      12'hC30: dout <= 8'b11111011; // 3120 : 251 - 0xfb -- Background 0xc3
      12'hC31: dout <= 8'b11111111; // 3121 : 255 - 0xff
      12'hC32: dout <= 8'b01111111; // 3122 : 127 - 0x7f
      12'hC33: dout <= 8'b00111111; // 3123 :  63 - 0x3f
      12'hC34: dout <= 8'b00001111; // 3124 :  15 - 0xf
      12'hC35: dout <= 8'b00000111; // 3125 :   7 - 0x7
      12'hC36: dout <= 8'b00000001; // 3126 :   1 - 0x1
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b11111111; // 3128 : 255 - 0xff -- plane 1
      12'hC39: dout <= 8'b11111111; // 3129 : 255 - 0xff
      12'hC3A: dout <= 8'b01111111; // 3130 : 127 - 0x7f
      12'hC3B: dout <= 8'b00111111; // 3131 :  63 - 0x3f
      12'hC3C: dout <= 8'b00001111; // 3132 :  15 - 0xf
      12'hC3D: dout <= 8'b00000111; // 3133 :   7 - 0x7
      12'hC3E: dout <= 8'b00000001; // 3134 :   1 - 0x1
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Background 0xc4
      12'hC41: dout <= 8'b10000000; // 3137 : 128 - 0x80
      12'hC42: dout <= 8'b01000000; // 3138 :  64 - 0x40
      12'hC43: dout <= 8'b11100000; // 3139 : 224 - 0xe0
      12'hC44: dout <= 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout <= 8'b00000000; // 3141 :   0 - 0x0
      12'hC46: dout <= 8'b00000100; // 3142 :   4 - 0x4
      12'hC47: dout <= 8'b11111111; // 3143 : 255 - 0xff
      12'hC48: dout <= 8'b11000000; // 3144 : 192 - 0xc0 -- plane 1
      12'hC49: dout <= 8'b11100000; // 3145 : 224 - 0xe0
      12'hC4A: dout <= 8'b11110000; // 3146 : 240 - 0xf0
      12'hC4B: dout <= 8'b11100000; // 3147 : 224 - 0xe0
      12'hC4C: dout <= 8'b11100001; // 3148 : 225 - 0xe1
      12'hC4D: dout <= 8'b11000011; // 3149 : 195 - 0xc3
      12'hC4E: dout <= 8'b00000111; // 3150 :   7 - 0x7
      12'hC4F: dout <= 8'b11111111; // 3151 : 255 - 0xff
      12'hC50: dout <= 8'b11111110; // 3152 : 254 - 0xfe -- Background 0xc5
      12'hC51: dout <= 8'b11111110; // 3153 : 254 - 0xfe
      12'hC52: dout <= 8'b11111110; // 3154 : 254 - 0xfe
      12'hC53: dout <= 8'b11111111; // 3155 : 255 - 0xff
      12'hC54: dout <= 8'b11111111; // 3156 : 255 - 0xff
      12'hC55: dout <= 8'b11111111; // 3157 : 255 - 0xff
      12'hC56: dout <= 8'b11111111; // 3158 : 255 - 0xff
      12'hC57: dout <= 8'b01111111; // 3159 : 127 - 0x7f
      12'hC58: dout <= 8'b11111111; // 3160 : 255 - 0xff -- plane 1
      12'hC59: dout <= 8'b11111111; // 3161 : 255 - 0xff
      12'hC5A: dout <= 8'b11111111; // 3162 : 255 - 0xff
      12'hC5B: dout <= 8'b11111111; // 3163 : 255 - 0xff
      12'hC5C: dout <= 8'b11111111; // 3164 : 255 - 0xff
      12'hC5D: dout <= 8'b11111111; // 3165 : 255 - 0xff
      12'hC5E: dout <= 8'b11111111; // 3166 : 255 - 0xff
      12'hC5F: dout <= 8'b01111111; // 3167 : 127 - 0x7f
      12'hC60: dout <= 8'b00111111; // 3168 :  63 - 0x3f -- Background 0xc6
      12'hC61: dout <= 8'b00011101; // 3169 :  29 - 0x1d
      12'hC62: dout <= 8'b00011110; // 3170 :  30 - 0x1e
      12'hC63: dout <= 8'b00011110; // 3171 :  30 - 0x1e
      12'hC64: dout <= 8'b00001101; // 3172 :  13 - 0xd
      12'hC65: dout <= 8'b00011110; // 3173 :  30 - 0x1e
      12'hC66: dout <= 8'b00111111; // 3174 :  63 - 0x3f
      12'hC67: dout <= 8'b01111111; // 3175 : 127 - 0x7f
      12'hC68: dout <= 8'b00111111; // 3176 :  63 - 0x3f -- plane 1
      12'hC69: dout <= 8'b00011111; // 3177 :  31 - 0x1f
      12'hC6A: dout <= 8'b00011111; // 3178 :  31 - 0x1f
      12'hC6B: dout <= 8'b00011111; // 3179 :  31 - 0x1f
      12'hC6C: dout <= 8'b00011111; // 3180 :  31 - 0x1f
      12'hC6D: dout <= 8'b00111111; // 3181 :  63 - 0x3f
      12'hC6E: dout <= 8'b01111111; // 3182 : 127 - 0x7f
      12'hC6F: dout <= 8'b11111111; // 3183 : 255 - 0xff
      12'hC70: dout <= 8'b11111111; // 3184 : 255 - 0xff -- Background 0xc7
      12'hC71: dout <= 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout <= 8'b11111111; // 3186 : 255 - 0xff
      12'hC73: dout <= 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout <= 8'b11111111; // 3188 : 255 - 0xff
      12'hC75: dout <= 8'b00111001; // 3189 :  57 - 0x39
      12'hC76: dout <= 8'b01000010; // 3190 :  66 - 0x42
      12'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      12'hC78: dout <= 8'b11111111; // 3192 : 255 - 0xff -- plane 1
      12'hC79: dout <= 8'b11111111; // 3193 : 255 - 0xff
      12'hC7A: dout <= 8'b11111111; // 3194 : 255 - 0xff
      12'hC7B: dout <= 8'b11111111; // 3195 : 255 - 0xff
      12'hC7C: dout <= 8'b11111111; // 3196 : 255 - 0xff
      12'hC7D: dout <= 8'b11111111; // 3197 : 255 - 0xff
      12'hC7E: dout <= 8'b11111111; // 3198 : 255 - 0xff
      12'hC7F: dout <= 8'b11111111; // 3199 : 255 - 0xff
      12'hC80: dout <= 8'b01101111; // 3200 : 111 - 0x6f -- Background 0xc8
      12'hC81: dout <= 8'b11011011; // 3201 : 219 - 0xdb
      12'hC82: dout <= 8'b00000011; // 3202 :   3 - 0x3
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      12'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      12'hC88: dout <= 8'b11111111; // 3208 : 255 - 0xff -- plane 1
      12'hC89: dout <= 8'b11111111; // 3209 : 255 - 0xff
      12'hC8A: dout <= 8'b00000011; // 3210 :   3 - 0x3
      12'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00000000; // 3216 :   0 - 0x0 -- Background 0xc9
      12'hC91: dout <= 8'b00000000; // 3217 :   0 - 0x0
      12'hC92: dout <= 8'b00000000; // 3218 :   0 - 0x0
      12'hC93: dout <= 8'b00000000; // 3219 :   0 - 0x0
      12'hC94: dout <= 8'b00000000; // 3220 :   0 - 0x0
      12'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      12'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      12'hC97: dout <= 8'b11100000; // 3223 : 224 - 0xe0
      12'hC98: dout <= 8'b00000000; // 3224 :   0 - 0x0 -- plane 1
      12'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      12'hC9A: dout <= 8'b00000000; // 3226 :   0 - 0x0
      12'hC9B: dout <= 8'b00000000; // 3227 :   0 - 0x0
      12'hC9C: dout <= 8'b10000000; // 3228 : 128 - 0x80
      12'hC9D: dout <= 8'b11000000; // 3229 : 192 - 0xc0
      12'hC9E: dout <= 8'b11000000; // 3230 : 192 - 0xc0
      12'hC9F: dout <= 8'b11110000; // 3231 : 240 - 0xf0
      12'hCA0: dout <= 8'b01110000; // 3232 : 112 - 0x70 -- Background 0xca
      12'hCA1: dout <= 8'b01111100; // 3233 : 124 - 0x7c
      12'hCA2: dout <= 8'b01111110; // 3234 : 126 - 0x7e
      12'hCA3: dout <= 8'b11111111; // 3235 : 255 - 0xff
      12'hCA4: dout <= 8'b11111111; // 3236 : 255 - 0xff
      12'hCA5: dout <= 8'b11110111; // 3237 : 247 - 0xf7
      12'hCA6: dout <= 8'b11101111; // 3238 : 239 - 0xef
      12'hCA7: dout <= 8'b00011111; // 3239 :  31 - 0x1f
      12'hCA8: dout <= 8'b11111100; // 3240 : 252 - 0xfc -- plane 1
      12'hCA9: dout <= 8'b11111110; // 3241 : 254 - 0xfe
      12'hCAA: dout <= 8'b11111111; // 3242 : 255 - 0xff
      12'hCAB: dout <= 8'b11111111; // 3243 : 255 - 0xff
      12'hCAC: dout <= 8'b11111111; // 3244 : 255 - 0xff
      12'hCAD: dout <= 8'b11111111; // 3245 : 255 - 0xff
      12'hCAE: dout <= 8'b11111111; // 3246 : 255 - 0xff
      12'hCAF: dout <= 8'b11111111; // 3247 : 255 - 0xff
      12'hCB0: dout <= 8'b11111111; // 3248 : 255 - 0xff -- Background 0xcb
      12'hCB1: dout <= 8'b11111111; // 3249 : 255 - 0xff
      12'hCB2: dout <= 8'b11111111; // 3250 : 255 - 0xff
      12'hCB3: dout <= 8'b11111000; // 3251 : 248 - 0xf8
      12'hCB4: dout <= 8'b11111000; // 3252 : 248 - 0xf8
      12'hCB5: dout <= 8'b11111110; // 3253 : 254 - 0xfe
      12'hCB6: dout <= 8'b11111111; // 3254 : 255 - 0xff
      12'hCB7: dout <= 8'b11111111; // 3255 : 255 - 0xff
      12'hCB8: dout <= 8'b11111111; // 3256 : 255 - 0xff -- plane 1
      12'hCB9: dout <= 8'b11111111; // 3257 : 255 - 0xff
      12'hCBA: dout <= 8'b11111111; // 3258 : 255 - 0xff
      12'hCBB: dout <= 8'b11111000; // 3259 : 248 - 0xf8
      12'hCBC: dout <= 8'b11111110; // 3260 : 254 - 0xfe
      12'hCBD: dout <= 8'b11111111; // 3261 : 255 - 0xff
      12'hCBE: dout <= 8'b11111111; // 3262 : 255 - 0xff
      12'hCBF: dout <= 8'b11111111; // 3263 : 255 - 0xff
      12'hCC0: dout <= 8'b11111111; // 3264 : 255 - 0xff -- Background 0xcc
      12'hCC1: dout <= 8'b11111111; // 3265 : 255 - 0xff
      12'hCC2: dout <= 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout <= 8'b00111111; // 3267 :  63 - 0x3f
      12'hCC4: dout <= 8'b00011110; // 3268 :  30 - 0x1e
      12'hCC5: dout <= 8'b00000001; // 3269 :   1 - 0x1
      12'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b11111111; // 3272 : 255 - 0xff -- plane 1
      12'hCC9: dout <= 8'b11111111; // 3273 : 255 - 0xff
      12'hCCA: dout <= 8'b11111111; // 3274 : 255 - 0xff
      12'hCCB: dout <= 8'b00111111; // 3275 :  63 - 0x3f
      12'hCCC: dout <= 8'b00011111; // 3276 :  31 - 0x1f
      12'hCCD: dout <= 8'b00011111; // 3277 :  31 - 0x1f
      12'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Background 0xcd
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout <= 8'b10000000; // 3283 : 128 - 0x80
      12'hCD4: dout <= 8'b11000000; // 3284 : 192 - 0xc0
      12'hCD5: dout <= 8'b11100000; // 3285 : 224 - 0xe0
      12'hCD6: dout <= 8'b11100000; // 3286 : 224 - 0xe0
      12'hCD7: dout <= 8'b11100000; // 3287 : 224 - 0xe0
      12'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b10000000; // 3290 : 128 - 0x80
      12'hCDB: dout <= 8'b11000000; // 3291 : 192 - 0xc0
      12'hCDC: dout <= 8'b11100000; // 3292 : 224 - 0xe0
      12'hCDD: dout <= 8'b11100000; // 3293 : 224 - 0xe0
      12'hCDE: dout <= 8'b11100000; // 3294 : 224 - 0xe0
      12'hCDF: dout <= 8'b11100000; // 3295 : 224 - 0xe0
      12'hCE0: dout <= 8'b11000000; // 3296 : 192 - 0xc0 -- Background 0xce
      12'hCE1: dout <= 8'b10000000; // 3297 : 128 - 0x80
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      12'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      12'hCE6: dout <= 8'b10000000; // 3302 : 128 - 0x80
      12'hCE7: dout <= 8'b10000000; // 3303 : 128 - 0x80
      12'hCE8: dout <= 8'b11000000; // 3304 : 192 - 0xc0 -- plane 1
      12'hCE9: dout <= 8'b10000000; // 3305 : 128 - 0x80
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      12'hCEC: dout <= 8'b00000000; // 3308 :   0 - 0x0
      12'hCED: dout <= 8'b10000000; // 3309 : 128 - 0x80
      12'hCEE: dout <= 8'b11000000; // 3310 : 192 - 0xc0
      12'hCEF: dout <= 8'b11000000; // 3311 : 192 - 0xc0
      12'hCF0: dout <= 8'b10000000; // 3312 : 128 - 0x80 -- Background 0xcf
      12'hCF1: dout <= 8'b10000000; // 3313 : 128 - 0x80
      12'hCF2: dout <= 8'b11100000; // 3314 : 224 - 0xe0
      12'hCF3: dout <= 8'b11000000; // 3315 : 192 - 0xc0
      12'hCF4: dout <= 8'b00100000; // 3316 :  32 - 0x20
      12'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      12'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout <= 8'b11000000; // 3320 : 192 - 0xc0 -- plane 1
      12'hCF9: dout <= 8'b11000000; // 3321 : 192 - 0xc0
      12'hCFA: dout <= 8'b11100000; // 3322 : 224 - 0xe0
      12'hCFB: dout <= 8'b11111000; // 3323 : 248 - 0xf8
      12'hCFC: dout <= 8'b11111100; // 3324 : 252 - 0xfc
      12'hCFD: dout <= 8'b11111100; // 3325 : 252 - 0xfc
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b00011111; // 3328 :  31 - 0x1f -- Background 0xd0
      12'hD01: dout <= 8'b00000110; // 3329 :   6 - 0x6
      12'hD02: dout <= 8'b00000110; // 3330 :   6 - 0x6
      12'hD03: dout <= 8'b00000110; // 3331 :   6 - 0x6
      12'hD04: dout <= 8'b00000110; // 3332 :   6 - 0x6
      12'hD05: dout <= 8'b00000110; // 3333 :   6 - 0x6
      12'hD06: dout <= 8'b00000110; // 3334 :   6 - 0x6
      12'hD07: dout <= 8'b00000000; // 3335 :   0 - 0x0
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b00000000; // 3338 :   0 - 0x0
      12'hD0B: dout <= 8'b00000000; // 3339 :   0 - 0x0
      12'hD0C: dout <= 8'b00000000; // 3340 :   0 - 0x0
      12'hD0D: dout <= 8'b00000000; // 3341 :   0 - 0x0
      12'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00111001; // 3344 :  57 - 0x39 -- Background 0xd1
      12'hD11: dout <= 8'b01100101; // 3345 : 101 - 0x65
      12'hD12: dout <= 8'b01100101; // 3346 : 101 - 0x65
      12'hD13: dout <= 8'b01100101; // 3347 : 101 - 0x65
      12'hD14: dout <= 8'b01100101; // 3348 : 101 - 0x65
      12'hD15: dout <= 8'b01100101; // 3349 : 101 - 0x65
      12'hD16: dout <= 8'b00111001; // 3350 :  57 - 0x39
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout <= 8'b00000000; // 3354 :   0 - 0x0
      12'hD1B: dout <= 8'b00000000; // 3355 :   0 - 0x0
      12'hD1C: dout <= 8'b00000000; // 3356 :   0 - 0x0
      12'hD1D: dout <= 8'b00000000; // 3357 :   0 - 0x0
      12'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b11100000; // 3360 : 224 - 0xe0 -- Background 0xd2
      12'hD21: dout <= 8'b10110000; // 3361 : 176 - 0xb0
      12'hD22: dout <= 8'b10110000; // 3362 : 176 - 0xb0
      12'hD23: dout <= 8'b10110110; // 3363 : 182 - 0xb6
      12'hD24: dout <= 8'b11100110; // 3364 : 230 - 0xe6
      12'hD25: dout <= 8'b10000000; // 3365 : 128 - 0x80
      12'hD26: dout <= 8'b10000000; // 3366 : 128 - 0x80
      12'hD27: dout <= 8'b00000000; // 3367 :   0 - 0x0
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout <= 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout <= 8'b00000000; // 3372 :   0 - 0x0
      12'hD2D: dout <= 8'b00000000; // 3373 :   0 - 0x0
      12'hD2E: dout <= 8'b00000000; // 3374 :   0 - 0x0
      12'hD2F: dout <= 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout <= 8'b00111100; // 3376 :  60 - 0x3c -- Background 0xd3
      12'hD31: dout <= 8'b01000010; // 3377 :  66 - 0x42
      12'hD32: dout <= 8'b10011001; // 3378 : 153 - 0x99
      12'hD33: dout <= 8'b10100001; // 3379 : 161 - 0xa1
      12'hD34: dout <= 8'b10100001; // 3380 : 161 - 0xa1
      12'hD35: dout <= 8'b10011001; // 3381 : 153 - 0x99
      12'hD36: dout <= 8'b01000010; // 3382 :  66 - 0x42
      12'hD37: dout <= 8'b00111100; // 3383 :  60 - 0x3c
      12'hD38: dout <= 8'b00000000; // 3384 :   0 - 0x0 -- plane 1
      12'hD39: dout <= 8'b00000000; // 3385 :   0 - 0x0
      12'hD3A: dout <= 8'b00000000; // 3386 :   0 - 0x0
      12'hD3B: dout <= 8'b00000000; // 3387 :   0 - 0x0
      12'hD3C: dout <= 8'b00000000; // 3388 :   0 - 0x0
      12'hD3D: dout <= 8'b00000000; // 3389 :   0 - 0x0
      12'hD3E: dout <= 8'b00000000; // 3390 :   0 - 0x0
      12'hD3F: dout <= 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xd4
      12'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout <= 8'b00000011; // 3395 :   3 - 0x3
      12'hD44: dout <= 8'b00000110; // 3396 :   6 - 0x6
      12'hD45: dout <= 8'b00000000; // 3397 :   0 - 0x0
      12'hD46: dout <= 8'b00000001; // 3398 :   1 - 0x1
      12'hD47: dout <= 8'b00000111; // 3399 :   7 - 0x7
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout <= 8'b00000011; // 3404 :   3 - 0x3
      12'hD4D: dout <= 8'b00000111; // 3405 :   7 - 0x7
      12'hD4E: dout <= 8'b00000011; // 3406 :   3 - 0x3
      12'hD4F: dout <= 8'b00000111; // 3407 :   7 - 0x7
      12'hD50: dout <= 8'b00001111; // 3408 :  15 - 0xf -- Background 0xd5
      12'hD51: dout <= 8'b00011111; // 3409 :  31 - 0x1f
      12'hD52: dout <= 8'b00111111; // 3410 :  63 - 0x3f
      12'hD53: dout <= 8'b01111111; // 3411 : 127 - 0x7f
      12'hD54: dout <= 8'b01111111; // 3412 : 127 - 0x7f
      12'hD55: dout <= 8'b01111111; // 3413 : 127 - 0x7f
      12'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout <= 8'b01111111; // 3415 : 127 - 0x7f
      12'hD58: dout <= 8'b00011111; // 3416 :  31 - 0x1f -- plane 1
      12'hD59: dout <= 8'b00111111; // 3417 :  63 - 0x3f
      12'hD5A: dout <= 8'b01111111; // 3418 : 127 - 0x7f
      12'hD5B: dout <= 8'b11111111; // 3419 : 255 - 0xff
      12'hD5C: dout <= 8'b11111111; // 3420 : 255 - 0xff
      12'hD5D: dout <= 8'b11111111; // 3421 : 255 - 0xff
      12'hD5E: dout <= 8'b11111111; // 3422 : 255 - 0xff
      12'hD5F: dout <= 8'b01111111; // 3423 : 127 - 0x7f
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xd6
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout <= 8'b10000000; // 3427 : 128 - 0x80
      12'hD64: dout <= 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout <= 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout <= 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout <= 8'b10100000; // 3431 : 160 - 0xa0
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout <= 8'b11000000; // 3435 : 192 - 0xc0
      12'hD6C: dout <= 8'b11100000; // 3436 : 224 - 0xe0
      12'hD6D: dout <= 8'b11110000; // 3437 : 240 - 0xf0
      12'hD6E: dout <= 8'b11110000; // 3438 : 240 - 0xf0
      12'hD6F: dout <= 8'b11111000; // 3439 : 248 - 0xf8
      12'hD70: dout <= 8'b11100000; // 3440 : 224 - 0xe0 -- Background 0xd7
      12'hD71: dout <= 8'b11110000; // 3441 : 240 - 0xf0
      12'hD72: dout <= 8'b11100000; // 3442 : 224 - 0xe0
      12'hD73: dout <= 8'b11011101; // 3443 : 221 - 0xdd
      12'hD74: dout <= 8'b11111010; // 3444 : 250 - 0xfa
      12'hD75: dout <= 8'b11101011; // 3445 : 235 - 0xeb
      12'hD76: dout <= 8'b10000000; // 3446 : 128 - 0x80
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b11111100; // 3448 : 252 - 0xfc -- plane 1
      12'hD79: dout <= 8'b11111000; // 3449 : 248 - 0xf8
      12'hD7A: dout <= 8'b11110000; // 3450 : 240 - 0xf0
      12'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      12'hD7C: dout <= 8'b11111111; // 3452 : 255 - 0xff
      12'hD7D: dout <= 8'b11111111; // 3453 : 255 - 0xff
      12'hD7E: dout <= 8'b11111111; // 3454 : 255 - 0xff
      12'hD7F: dout <= 8'b11111111; // 3455 : 255 - 0xff
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xd8
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      12'hD83: dout <= 8'b00000011; // 3459 :   3 - 0x3
      12'hD84: dout <= 8'b00000110; // 3460 :   6 - 0x6
      12'hD85: dout <= 8'b00000000; // 3461 :   0 - 0x0
      12'hD86: dout <= 8'b00000001; // 3462 :   1 - 0x1
      12'hD87: dout <= 8'b00000001; // 3463 :   1 - 0x1
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- plane 1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b00000000; // 3466 :   0 - 0x0
      12'hD8B: dout <= 8'b00000000; // 3467 :   0 - 0x0
      12'hD8C: dout <= 8'b00000011; // 3468 :   3 - 0x3
      12'hD8D: dout <= 8'b00000111; // 3469 :   7 - 0x7
      12'hD8E: dout <= 8'b00001111; // 3470 :  15 - 0xf
      12'hD8F: dout <= 8'b00011111; // 3471 :  31 - 0x1f
      12'hD90: dout <= 8'b00001011; // 3472 :  11 - 0xb -- Background 0xd9
      12'hD91: dout <= 8'b00000111; // 3473 :   7 - 0x7
      12'hD92: dout <= 8'b00000011; // 3474 :   3 - 0x3
      12'hD93: dout <= 8'b01011101; // 3475 :  93 - 0x5d
      12'hD94: dout <= 8'b10101111; // 3476 : 175 - 0xaf
      12'hD95: dout <= 8'b01010011; // 3477 :  83 - 0x53
      12'hD96: dout <= 8'b00000000; // 3478 :   0 - 0x0
      12'hD97: dout <= 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout <= 8'b00111111; // 3480 :  63 - 0x3f -- plane 1
      12'hD99: dout <= 8'b00011111; // 3481 :  31 - 0x1f
      12'hD9A: dout <= 8'b00000111; // 3482 :   7 - 0x7
      12'hD9B: dout <= 8'b11111111; // 3483 : 255 - 0xff
      12'hD9C: dout <= 8'b11111111; // 3484 : 255 - 0xff
      12'hD9D: dout <= 8'b11111111; // 3485 : 255 - 0xff
      12'hD9E: dout <= 8'b11111111; // 3486 : 255 - 0xff
      12'hD9F: dout <= 8'b11111111; // 3487 : 255 - 0xff
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xda
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout <= 8'b10000000; // 3491 : 128 - 0x80
      12'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      12'hDA5: dout <= 8'b00000000; // 3493 :   0 - 0x0
      12'hDA6: dout <= 8'b01100000; // 3494 :  96 - 0x60
      12'hDA7: dout <= 8'b11110000; // 3495 : 240 - 0xf0
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b11000000; // 3499 : 192 - 0xc0
      12'hDAC: dout <= 8'b11000000; // 3500 : 192 - 0xc0
      12'hDAD: dout <= 8'b11000000; // 3501 : 192 - 0xc0
      12'hDAE: dout <= 8'b11100000; // 3502 : 224 - 0xe0
      12'hDAF: dout <= 8'b11111000; // 3503 : 248 - 0xf8
      12'hDB0: dout <= 8'b11111000; // 3504 : 248 - 0xf8 -- Background 0xdb
      12'hDB1: dout <= 8'b11111100; // 3505 : 252 - 0xfc
      12'hDB2: dout <= 8'b11111100; // 3506 : 252 - 0xfc
      12'hDB3: dout <= 8'b11111110; // 3507 : 254 - 0xfe
      12'hDB4: dout <= 8'b11111110; // 3508 : 254 - 0xfe
      12'hDB5: dout <= 8'b11111111; // 3509 : 255 - 0xff
      12'hDB6: dout <= 8'b11111111; // 3510 : 255 - 0xff
      12'hDB7: dout <= 8'b01111110; // 3511 : 126 - 0x7e
      12'hDB8: dout <= 8'b11111100; // 3512 : 252 - 0xfc -- plane 1
      12'hDB9: dout <= 8'b11111110; // 3513 : 254 - 0xfe
      12'hDBA: dout <= 8'b11111110; // 3514 : 254 - 0xfe
      12'hDBB: dout <= 8'b11111111; // 3515 : 255 - 0xff
      12'hDBC: dout <= 8'b11111111; // 3516 : 255 - 0xff
      12'hDBD: dout <= 8'b11111111; // 3517 : 255 - 0xff
      12'hDBE: dout <= 8'b11111111; // 3518 : 255 - 0xff
      12'hDBF: dout <= 8'b11111110; // 3519 : 254 - 0xfe
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xdc
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      12'hDC3: dout <= 8'b00000000; // 3523 :   0 - 0x0
      12'hDC4: dout <= 8'b00000000; // 3524 :   0 - 0x0
      12'hDC5: dout <= 8'b00000000; // 3525 :   0 - 0x0
      12'hDC6: dout <= 8'b00100001; // 3526 :  33 - 0x21
      12'hDC7: dout <= 8'b00111111; // 3527 :  63 - 0x3f
      12'hDC8: dout <= 8'b00110110; // 3528 :  54 - 0x36 -- plane 1
      12'hDC9: dout <= 8'b00110110; // 3529 :  54 - 0x36
      12'hDCA: dout <= 8'b01111110; // 3530 : 126 - 0x7e
      12'hDCB: dout <= 8'b01111111; // 3531 : 127 - 0x7f
      12'hDCC: dout <= 8'b01111111; // 3532 : 127 - 0x7f
      12'hDCD: dout <= 8'b01111111; // 3533 : 127 - 0x7f
      12'hDCE: dout <= 8'b00111111; // 3534 :  63 - 0x3f
      12'hDCF: dout <= 8'b00111111; // 3535 :  63 - 0x3f
      12'hDD0: dout <= 8'b00111111; // 3536 :  63 - 0x3f -- Background 0xdd
      12'hDD1: dout <= 8'b00011111; // 3537 :  31 - 0x1f
      12'hDD2: dout <= 8'b00011111; // 3538 :  31 - 0x1f
      12'hDD3: dout <= 8'b00001111; // 3539 :  15 - 0xf
      12'hDD4: dout <= 8'b00000111; // 3540 :   7 - 0x7
      12'hDD5: dout <= 8'b00000011; // 3541 :   3 - 0x3
      12'hDD6: dout <= 8'b00000000; // 3542 :   0 - 0x0
      12'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout <= 8'b00111111; // 3544 :  63 - 0x3f -- plane 1
      12'hDD9: dout <= 8'b00011111; // 3545 :  31 - 0x1f
      12'hDDA: dout <= 8'b00011111; // 3546 :  31 - 0x1f
      12'hDDB: dout <= 8'b00001111; // 3547 :  15 - 0xf
      12'hDDC: dout <= 8'b00000111; // 3548 :   7 - 0x7
      12'hDDD: dout <= 8'b00000011; // 3549 :   3 - 0x3
      12'hDDE: dout <= 8'b00000000; // 3550 :   0 - 0x0
      12'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout <= 8'b00111110; // 3552 :  62 - 0x3e -- Background 0xde
      12'hDE1: dout <= 8'b00011110; // 3553 :  30 - 0x1e
      12'hDE2: dout <= 8'b00011110; // 3554 :  30 - 0x1e
      12'hDE3: dout <= 8'b00001110; // 3555 :  14 - 0xe
      12'hDE4: dout <= 8'b00001111; // 3556 :  15 - 0xf
      12'hDE5: dout <= 8'b00011111; // 3557 :  31 - 0x1f
      12'hDE6: dout <= 8'b10011111; // 3558 : 159 - 0x9f
      12'hDE7: dout <= 8'b10011111; // 3559 : 159 - 0x9f
      12'hDE8: dout <= 8'b00111111; // 3560 :  63 - 0x3f -- plane 1
      12'hDE9: dout <= 8'b00011111; // 3561 :  31 - 0x1f
      12'hDEA: dout <= 8'b11011111; // 3562 : 223 - 0xdf
      12'hDEB: dout <= 8'b11001111; // 3563 : 207 - 0xcf
      12'hDEC: dout <= 8'b11001111; // 3564 : 207 - 0xcf
      12'hDED: dout <= 8'b10011111; // 3565 : 159 - 0x9f
      12'hDEE: dout <= 8'b11011111; // 3566 : 223 - 0xdf
      12'hDEF: dout <= 8'b11111111; // 3567 : 255 - 0xff
      12'hDF0: dout <= 8'b11011111; // 3568 : 223 - 0xdf -- Background 0xdf
      12'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout <= 8'b11111111; // 3570 : 255 - 0xff
      12'hDF3: dout <= 8'b11111111; // 3571 : 255 - 0xff
      12'hDF4: dout <= 8'b11111111; // 3572 : 255 - 0xff
      12'hDF5: dout <= 8'b11011111; // 3573 : 223 - 0xdf
      12'hDF6: dout <= 8'b11100111; // 3574 : 231 - 0xe7
      12'hDF7: dout <= 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout <= 8'b11111111; // 3576 : 255 - 0xff -- plane 1
      12'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      12'hDFA: dout <= 8'b11111111; // 3578 : 255 - 0xff
      12'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout <= 8'b11111111; // 3580 : 255 - 0xff
      12'hDFD: dout <= 8'b11111111; // 3581 : 255 - 0xff
      12'hDFE: dout <= 8'b11111111; // 3582 : 255 - 0xff
      12'hDFF: dout <= 8'b00001111; // 3583 :  15 - 0xf
      12'hE00: dout <= 8'b00100000; // 3584 :  32 - 0x20 -- Background 0xe0
      12'hE01: dout <= 8'b00001111; // 3585 :  15 - 0xf
      12'hE02: dout <= 8'b00110000; // 3586 :  48 - 0x30
      12'hE03: dout <= 8'b01000000; // 3587 :  64 - 0x40
      12'hE04: dout <= 8'b10011000; // 3588 : 152 - 0x98
      12'hE05: dout <= 8'b00111110; // 3589 :  62 - 0x3e
      12'hE06: dout <= 8'b00011111; // 3590 :  31 - 0x1f
      12'hE07: dout <= 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout <= 8'b11111111; // 3592 : 255 - 0xff -- plane 1
      12'hE09: dout <= 8'b11111111; // 3593 : 255 - 0xff
      12'hE0A: dout <= 8'b11111111; // 3594 : 255 - 0xff
      12'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      12'hE0C: dout <= 8'b11111111; // 3596 : 255 - 0xff
      12'hE0D: dout <= 8'b11111111; // 3597 : 255 - 0xff
      12'hE0E: dout <= 8'b11111111; // 3598 : 255 - 0xff
      12'hE0F: dout <= 8'b11111111; // 3599 : 255 - 0xff
      12'hE10: dout <= 8'b10000001; // 3600 : 129 - 0x81 -- Background 0xe1
      12'hE11: dout <= 8'b00110110; // 3601 :  54 - 0x36
      12'hE12: dout <= 8'b00101110; // 3602 :  46 - 0x2e
      12'hE13: dout <= 8'b10101111; // 3603 : 175 - 0xaf
      12'hE14: dout <= 8'b10101110; // 3604 : 174 - 0xae
      12'hE15: dout <= 8'b11010001; // 3605 : 209 - 0xd1
      12'hE16: dout <= 8'b11101111; // 3606 : 239 - 0xef
      12'hE17: dout <= 8'b10000111; // 3607 : 135 - 0x87
      12'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout <= 8'b11111001; // 3609 : 249 - 0xf9
      12'hE1A: dout <= 8'b11110000; // 3610 : 240 - 0xf0
      12'hE1B: dout <= 8'b11110000; // 3611 : 240 - 0xf0
      12'hE1C: dout <= 8'b10110001; // 3612 : 177 - 0xb1
      12'hE1D: dout <= 8'b11011111; // 3613 : 223 - 0xdf
      12'hE1E: dout <= 8'b11101111; // 3614 : 239 - 0xef
      12'hE1F: dout <= 8'b10000111; // 3615 : 135 - 0x87
      12'hE20: dout <= 8'b00000010; // 3616 :   2 - 0x2 -- Background 0xe2
      12'hE21: dout <= 8'b11111000; // 3617 : 248 - 0xf8
      12'hE22: dout <= 8'b00000110; // 3618 :   6 - 0x6
      12'hE23: dout <= 8'b00000001; // 3619 :   1 - 0x1
      12'hE24: dout <= 8'b00001100; // 3620 :  12 - 0xc
      12'hE25: dout <= 8'b00111110; // 3621 :  62 - 0x3e
      12'hE26: dout <= 8'b11111100; // 3622 : 252 - 0xfc
      12'hE27: dout <= 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout <= 8'b11111111; // 3624 : 255 - 0xff -- plane 1
      12'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout <= 8'b11111111; // 3626 : 255 - 0xff
      12'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout <= 8'b11111111; // 3628 : 255 - 0xff
      12'hE2D: dout <= 8'b11111111; // 3629 : 255 - 0xff
      12'hE2E: dout <= 8'b11111111; // 3630 : 255 - 0xff
      12'hE2F: dout <= 8'b11111111; // 3631 : 255 - 0xff
      12'hE30: dout <= 8'b11000000; // 3632 : 192 - 0xc0 -- Background 0xe3
      12'hE31: dout <= 8'b00110110; // 3633 :  54 - 0x36
      12'hE32: dout <= 8'b00111110; // 3634 :  62 - 0x3e
      12'hE33: dout <= 8'b01111010; // 3635 : 122 - 0x7a
      12'hE34: dout <= 8'b10110110; // 3636 : 182 - 0xb6
      12'hE35: dout <= 8'b11001101; // 3637 : 205 - 0xcd
      12'hE36: dout <= 8'b11111011; // 3638 : 251 - 0xfb
      12'hE37: dout <= 8'b11110000; // 3639 : 240 - 0xf0
      12'hE38: dout <= 8'b11111111; // 3640 : 255 - 0xff -- plane 1
      12'hE39: dout <= 8'b11001111; // 3641 : 207 - 0xcf
      12'hE3A: dout <= 8'b10000111; // 3642 : 135 - 0x87
      12'hE3B: dout <= 8'b10000111; // 3643 : 135 - 0x87
      12'hE3C: dout <= 8'b11001110; // 3644 : 206 - 0xce
      12'hE3D: dout <= 8'b11111101; // 3645 : 253 - 0xfd
      12'hE3E: dout <= 8'b11111011; // 3646 : 251 - 0xfb
      12'hE3F: dout <= 8'b11110000; // 3647 : 240 - 0xf0
      12'hE40: dout <= 8'b00111110; // 3648 :  62 - 0x3e -- Background 0xe4
      12'hE41: dout <= 8'b00111100; // 3649 :  60 - 0x3c
      12'hE42: dout <= 8'b00111100; // 3650 :  60 - 0x3c
      12'hE43: dout <= 8'b00111000; // 3651 :  56 - 0x38
      12'hE44: dout <= 8'b11111000; // 3652 : 248 - 0xf8
      12'hE45: dout <= 8'b01111100; // 3653 : 124 - 0x7c
      12'hE46: dout <= 8'b01111110; // 3654 : 126 - 0x7e
      12'hE47: dout <= 8'b01111000; // 3655 : 120 - 0x78
      12'hE48: dout <= 8'b11111110; // 3656 : 254 - 0xfe -- plane 1
      12'hE49: dout <= 8'b11111100; // 3657 : 252 - 0xfc
      12'hE4A: dout <= 8'b11111100; // 3658 : 252 - 0xfc
      12'hE4B: dout <= 8'b11111000; // 3659 : 248 - 0xf8
      12'hE4C: dout <= 8'b11111011; // 3660 : 251 - 0xfb
      12'hE4D: dout <= 8'b11111101; // 3661 : 253 - 0xfd
      12'hE4E: dout <= 8'b11111110; // 3662 : 254 - 0xfe
      12'hE4F: dout <= 8'b11111111; // 3663 : 255 - 0xff
      12'hE50: dout <= 8'b11111000; // 3664 : 248 - 0xf8 -- Background 0xe5
      12'hE51: dout <= 8'b01111111; // 3665 : 127 - 0x7f
      12'hE52: dout <= 8'b01111111; // 3666 : 127 - 0x7f
      12'hE53: dout <= 8'b11111110; // 3667 : 254 - 0xfe
      12'hE54: dout <= 8'b11111111; // 3668 : 255 - 0xff
      12'hE55: dout <= 8'b11111111; // 3669 : 255 - 0xff
      12'hE56: dout <= 8'b11110011; // 3670 : 243 - 0xf3
      12'hE57: dout <= 8'b10000001; // 3671 : 129 - 0x81
      12'hE58: dout <= 8'b11111111; // 3672 : 255 - 0xff -- plane 1
      12'hE59: dout <= 8'b11111111; // 3673 : 255 - 0xff
      12'hE5A: dout <= 8'b11111111; // 3674 : 255 - 0xff
      12'hE5B: dout <= 8'b11111111; // 3675 : 255 - 0xff
      12'hE5C: dout <= 8'b11111111; // 3676 : 255 - 0xff
      12'hE5D: dout <= 8'b11111111; // 3677 : 255 - 0xff
      12'hE5E: dout <= 8'b11111111; // 3678 : 255 - 0xff
      12'hE5F: dout <= 8'b11111001; // 3679 : 249 - 0xf9
      12'hE60: dout <= 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xe6
      12'hE61: dout <= 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout <= 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout <= 8'b00010000; // 3683 :  16 - 0x10
      12'hE64: dout <= 8'b01000000; // 3684 :  64 - 0x40
      12'hE65: dout <= 8'b00100000; // 3685 :  32 - 0x20
      12'hE66: dout <= 8'b00000000; // 3686 :   0 - 0x0
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- plane 1
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b01111000; // 3691 : 120 - 0x78
      12'hE6C: dout <= 8'b11111100; // 3692 : 252 - 0xfc
      12'hE6D: dout <= 8'b11111100; // 3693 : 252 - 0xfc
      12'hE6E: dout <= 8'b11111100; // 3694 : 252 - 0xfc
      12'hE6F: dout <= 8'b11111100; // 3695 : 252 - 0xfc
      12'hE70: dout <= 8'b00000110; // 3696 :   6 - 0x6 -- Background 0xe7
      12'hE71: dout <= 8'b00001110; // 3697 :  14 - 0xe
      12'hE72: dout <= 8'b01111110; // 3698 : 126 - 0x7e
      12'hE73: dout <= 8'b11111110; // 3699 : 254 - 0xfe
      12'hE74: dout <= 8'b11111110; // 3700 : 254 - 0xfe
      12'hE75: dout <= 8'b11111100; // 3701 : 252 - 0xfc
      12'hE76: dout <= 8'b11111000; // 3702 : 248 - 0xf8
      12'hE77: dout <= 8'b11110000; // 3703 : 240 - 0xf0
      12'hE78: dout <= 8'b11111110; // 3704 : 254 - 0xfe -- plane 1
      12'hE79: dout <= 8'b11111110; // 3705 : 254 - 0xfe
      12'hE7A: dout <= 8'b11111110; // 3706 : 254 - 0xfe
      12'hE7B: dout <= 8'b11111110; // 3707 : 254 - 0xfe
      12'hE7C: dout <= 8'b11111110; // 3708 : 254 - 0xfe
      12'hE7D: dout <= 8'b11111100; // 3709 : 252 - 0xfc
      12'hE7E: dout <= 8'b11111000; // 3710 : 248 - 0xf8
      12'hE7F: dout <= 8'b11110000; // 3711 : 240 - 0xf0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xe8
      12'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout <= 8'b00000000; // 3714 :   0 - 0x0
      12'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout <= 8'b00000000; // 3716 :   0 - 0x0
      12'hE85: dout <= 8'b00000000; // 3717 :   0 - 0x0
      12'hE86: dout <= 8'b00000000; // 3718 :   0 - 0x0
      12'hE87: dout <= 8'b00000001; // 3719 :   1 - 0x1
      12'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0 -- plane 1
      12'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout <= 8'b00000000; // 3722 :   0 - 0x0
      12'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout <= 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout <= 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b00000010; // 3728 :   2 - 0x2 -- Background 0xe9
      12'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      12'hE92: dout <= 8'b00001000; // 3730 :   8 - 0x8
      12'hE93: dout <= 8'b00000001; // 3731 :   1 - 0x1
      12'hE94: dout <= 8'b00010011; // 3732 :  19 - 0x13
      12'hE95: dout <= 8'b00000001; // 3733 :   1 - 0x1
      12'hE96: dout <= 8'b00000000; // 3734 :   0 - 0x0
      12'hE97: dout <= 8'b00000000; // 3735 :   0 - 0x0
      12'hE98: dout <= 8'b00000001; // 3736 :   1 - 0x1 -- plane 1
      12'hE99: dout <= 8'b00001111; // 3737 :  15 - 0xf
      12'hE9A: dout <= 8'b00011111; // 3738 :  31 - 0x1f
      12'hE9B: dout <= 8'b00011111; // 3739 :  31 - 0x1f
      12'hE9C: dout <= 8'b00111011; // 3740 :  59 - 0x3b
      12'hE9D: dout <= 8'b00110011; // 3741 :  51 - 0x33
      12'hE9E: dout <= 8'b00000001; // 3742 :   1 - 0x1
      12'hE9F: dout <= 8'b00000001; // 3743 :   1 - 0x1
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xea
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout <= 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout <= 8'b00000000; // 3750 :   0 - 0x0
      12'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0 -- plane 1
      12'hEA9: dout <= 8'b00000000; // 3753 :   0 - 0x0
      12'hEAA: dout <= 8'b00000000; // 3754 :   0 - 0x0
      12'hEAB: dout <= 8'b00110110; // 3755 :  54 - 0x36
      12'hEAC: dout <= 8'b01101100; // 3756 : 108 - 0x6c
      12'hEAD: dout <= 8'b11111101; // 3757 : 253 - 0xfd
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xeb
      12'hEB1: dout <= 8'b01000011; // 3761 :  67 - 0x43
      12'hEB2: dout <= 8'b01111111; // 3762 : 127 - 0x7f
      12'hEB3: dout <= 8'b01111111; // 3763 : 127 - 0x7f
      12'hEB4: dout <= 8'b01111111; // 3764 : 127 - 0x7f
      12'hEB5: dout <= 8'b00111111; // 3765 :  63 - 0x3f
      12'hEB6: dout <= 8'b00011111; // 3766 :  31 - 0x1f
      12'hEB7: dout <= 8'b00000111; // 3767 :   7 - 0x7
      12'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff -- plane 1
      12'hEB9: dout <= 8'b01111111; // 3769 : 127 - 0x7f
      12'hEBA: dout <= 8'b01111111; // 3770 : 127 - 0x7f
      12'hEBB: dout <= 8'b01111111; // 3771 : 127 - 0x7f
      12'hEBC: dout <= 8'b01111111; // 3772 : 127 - 0x7f
      12'hEBD: dout <= 8'b00111111; // 3773 :  63 - 0x3f
      12'hEBE: dout <= 8'b00011111; // 3774 :  31 - 0x1f
      12'hEBF: dout <= 8'b00000111; // 3775 :   7 - 0x7
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xec
      12'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout <= 8'b00000000; // 3779 :   0 - 0x0
      12'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout <= 8'b11000000; // 3782 : 192 - 0xc0
      12'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      12'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout <= 8'b11100000; // 3791 : 224 - 0xe0
      12'hED0: dout <= 8'b00010000; // 3792 :  16 - 0x10 -- Background 0xed
      12'hED1: dout <= 8'b00111000; // 3793 :  56 - 0x38
      12'hED2: dout <= 8'b10111111; // 3794 : 191 - 0xbf
      12'hED3: dout <= 8'b11111111; // 3795 : 255 - 0xff
      12'hED4: dout <= 8'b11111111; // 3796 : 255 - 0xff
      12'hED5: dout <= 8'b11111111; // 3797 : 255 - 0xff
      12'hED6: dout <= 8'b11111111; // 3798 : 255 - 0xff
      12'hED7: dout <= 8'b11111111; // 3799 : 255 - 0xff
      12'hED8: dout <= 8'b11111000; // 3800 : 248 - 0xf8 -- plane 1
      12'hED9: dout <= 8'b11111111; // 3801 : 255 - 0xff
      12'hEDA: dout <= 8'b11111111; // 3802 : 255 - 0xff
      12'hEDB: dout <= 8'b11111111; // 3803 : 255 - 0xff
      12'hEDC: dout <= 8'b11111111; // 3804 : 255 - 0xff
      12'hEDD: dout <= 8'b11111111; // 3805 : 255 - 0xff
      12'hEDE: dout <= 8'b11111111; // 3806 : 255 - 0xff
      12'hEDF: dout <= 8'b11111111; // 3807 : 255 - 0xff
      12'hEE0: dout <= 8'b01111110; // 3808 : 126 - 0x7e -- Background 0xee
      12'hEE1: dout <= 8'b00011110; // 3809 :  30 - 0x1e
      12'hEE2: dout <= 8'b00011110; // 3810 :  30 - 0x1e
      12'hEE3: dout <= 8'b00001110; // 3811 :  14 - 0xe
      12'hEE4: dout <= 8'b00001111; // 3812 :  15 - 0xf
      12'hEE5: dout <= 8'b00011110; // 3813 :  30 - 0x1e
      12'hEE6: dout <= 8'b00011110; // 3814 :  30 - 0x1e
      12'hEE7: dout <= 8'b00111110; // 3815 :  62 - 0x3e
      12'hEE8: dout <= 8'b11111111; // 3816 : 255 - 0xff -- plane 1
      12'hEE9: dout <= 8'b01111111; // 3817 : 127 - 0x7f
      12'hEEA: dout <= 8'b00011111; // 3818 :  31 - 0x1f
      12'hEEB: dout <= 8'b00001111; // 3819 :  15 - 0xf
      12'hEEC: dout <= 8'b00001111; // 3820 :  15 - 0xf
      12'hEED: dout <= 8'b10011111; // 3821 : 159 - 0x9f
      12'hEEE: dout <= 8'b10011111; // 3822 : 159 - 0x9f
      12'hEEF: dout <= 8'b10111111; // 3823 : 191 - 0xbf
      12'hEF0: dout <= 8'b01111111; // 3824 : 127 - 0x7f -- Background 0xef
      12'hEF1: dout <= 8'b01111111; // 3825 : 127 - 0x7f
      12'hEF2: dout <= 8'b10111111; // 3826 : 191 - 0xbf
      12'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout <= 8'b11111111; // 3828 : 255 - 0xff
      12'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout <= 8'b11100111; // 3830 : 231 - 0xe7
      12'hEF7: dout <= 8'b11000000; // 3831 : 192 - 0xc0
      12'hEF8: dout <= 8'b01111111; // 3832 : 127 - 0x7f -- plane 1
      12'hEF9: dout <= 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout <= 8'b11111111; // 3834 : 255 - 0xff
      12'hEFB: dout <= 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout <= 8'b11111111; // 3836 : 255 - 0xff
      12'hEFD: dout <= 8'b11111111; // 3837 : 255 - 0xff
      12'hEFE: dout <= 8'b11111111; // 3838 : 255 - 0xff
      12'hEFF: dout <= 8'b11001111; // 3839 : 207 - 0xcf
      12'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xf0
      12'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout <= 8'b00010000; // 3842 :  16 - 0x10
      12'hF03: dout <= 8'b11111101; // 3843 : 253 - 0xfd
      12'hF04: dout <= 8'b11111010; // 3844 : 250 - 0xfa
      12'hF05: dout <= 8'b11101011; // 3845 : 235 - 0xeb
      12'hF06: dout <= 8'b10000000; // 3846 : 128 - 0x80
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout <= 8'b11110000; // 3850 : 240 - 0xf0
      12'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      12'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      12'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      12'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout <= 8'b00100000; // 3856 :  32 - 0x20 -- Background 0xf1
      12'hF11: dout <= 8'b00011111; // 3857 :  31 - 0x1f
      12'hF12: dout <= 8'b01100000; // 3858 :  96 - 0x60
      12'hF13: dout <= 8'b10001110; // 3859 : 142 - 0x8e
      12'hF14: dout <= 8'b00111111; // 3860 :  63 - 0x3f
      12'hF15: dout <= 8'b01111111; // 3861 : 127 - 0x7f
      12'hF16: dout <= 8'b01111111; // 3862 : 127 - 0x7f
      12'hF17: dout <= 8'b01111100; // 3863 : 124 - 0x7c
      12'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff -- plane 1
      12'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      12'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      12'hF1B: dout <= 8'b11110001; // 3867 : 241 - 0xf1
      12'hF1C: dout <= 8'b11000100; // 3868 : 196 - 0xc4
      12'hF1D: dout <= 8'b11101110; // 3869 : 238 - 0xee
      12'hF1E: dout <= 8'b11000100; // 3870 : 196 - 0xc4
      12'hF1F: dout <= 8'b10000011; // 3871 : 131 - 0x83
      12'hF20: dout <= 8'b00111001; // 3872 :  57 - 0x39 -- Background 0xf2
      12'hF21: dout <= 8'b00110110; // 3873 :  54 - 0x36
      12'hF22: dout <= 8'b00101110; // 3874 :  46 - 0x2e
      12'hF23: dout <= 8'b10101111; // 3875 : 175 - 0xaf
      12'hF24: dout <= 8'b10101110; // 3876 : 174 - 0xae
      12'hF25: dout <= 8'b11010001; // 3877 : 209 - 0xd1
      12'hF26: dout <= 8'b11101111; // 3878 : 239 - 0xef
      12'hF27: dout <= 8'b10000111; // 3879 : 135 - 0x87
      12'hF28: dout <= 8'b11000111; // 3880 : 199 - 0xc7 -- plane 1
      12'hF29: dout <= 8'b11111001; // 3881 : 249 - 0xf9
      12'hF2A: dout <= 8'b11110000; // 3882 : 240 - 0xf0
      12'hF2B: dout <= 8'b11110000; // 3883 : 240 - 0xf0
      12'hF2C: dout <= 8'b10110001; // 3884 : 177 - 0xb1
      12'hF2D: dout <= 8'b11011111; // 3885 : 223 - 0xdf
      12'hF2E: dout <= 8'b11101111; // 3886 : 239 - 0xef
      12'hF2F: dout <= 8'b10000111; // 3887 : 135 - 0x87
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xf3
      12'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout <= 8'b00000100; // 3890 :   4 - 0x4
      12'hF33: dout <= 8'b01011111; // 3891 :  95 - 0x5f
      12'hF34: dout <= 8'b10101111; // 3892 : 175 - 0xaf
      12'hF35: dout <= 8'b01010011; // 3893 :  83 - 0x53
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b00000000; // 3896 :   0 - 0x0 -- plane 1
      12'hF39: dout <= 8'b00000000; // 3897 :   0 - 0x0
      12'hF3A: dout <= 8'b00000111; // 3898 :   7 - 0x7
      12'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      12'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      12'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      12'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      12'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      12'hF40: dout <= 8'b00000010; // 3904 :   2 - 0x2 -- Background 0xf4
      12'hF41: dout <= 8'b11111100; // 3905 : 252 - 0xfc
      12'hF42: dout <= 8'b00000011; // 3906 :   3 - 0x3
      12'hF43: dout <= 8'b00111000; // 3907 :  56 - 0x38
      12'hF44: dout <= 8'b11111110; // 3908 : 254 - 0xfe
      12'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout <= 8'b00011110; // 3911 :  30 - 0x1e
      12'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff -- plane 1
      12'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      12'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      12'hF4B: dout <= 8'b11000111; // 3915 : 199 - 0xc7
      12'hF4C: dout <= 8'b01000101; // 3916 :  69 - 0x45
      12'hF4D: dout <= 8'b11101110; // 3917 : 238 - 0xee
      12'hF4E: dout <= 8'b01000100; // 3918 :  68 - 0x44
      12'hF4F: dout <= 8'b11100001; // 3919 : 225 - 0xe1
      12'hF50: dout <= 8'b11000000; // 3920 : 192 - 0xc0 -- Background 0xf5
      12'hF51: dout <= 8'b00110110; // 3921 :  54 - 0x36
      12'hF52: dout <= 8'b00111110; // 3922 :  62 - 0x3e
      12'hF53: dout <= 8'b01111010; // 3923 : 122 - 0x7a
      12'hF54: dout <= 8'b10110110; // 3924 : 182 - 0xb6
      12'hF55: dout <= 8'b11001101; // 3925 : 205 - 0xcd
      12'hF56: dout <= 8'b11111011; // 3926 : 251 - 0xfb
      12'hF57: dout <= 8'b11110000; // 3927 : 240 - 0xf0
      12'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff -- plane 1
      12'hF59: dout <= 8'b11001111; // 3929 : 207 - 0xcf
      12'hF5A: dout <= 8'b10000111; // 3930 : 135 - 0x87
      12'hF5B: dout <= 8'b10000111; // 3931 : 135 - 0x87
      12'hF5C: dout <= 8'b11001110; // 3932 : 206 - 0xce
      12'hF5D: dout <= 8'b11111101; // 3933 : 253 - 0xfd
      12'hF5E: dout <= 8'b11111011; // 3934 : 251 - 0xfb
      12'hF5F: dout <= 8'b11110000; // 3935 : 240 - 0xf0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xf6
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00001110; // 3941 :  14 - 0xe
      12'hF66: dout <= 8'b00001000; // 3942 :   8 - 0x8
      12'hF67: dout <= 8'b00001000; // 3943 :   8 - 0x8
      12'hF68: dout <= 8'b00000000; // 3944 :   0 - 0x0 -- plane 1
      12'hF69: dout <= 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout <= 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00000001; // 3949 :   1 - 0x1
      12'hF6E: dout <= 8'b00000111; // 3950 :   7 - 0x7
      12'hF6F: dout <= 8'b00001111; // 3951 :  15 - 0xf
      12'hF70: dout <= 8'b00011111; // 3952 :  31 - 0x1f -- Background 0xf7
      12'hF71: dout <= 8'b00111111; // 3953 :  63 - 0x3f
      12'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      12'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      12'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      12'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      12'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      12'hF77: dout <= 8'b01111111; // 3959 : 127 - 0x7f
      12'hF78: dout <= 8'b00111111; // 3960 :  63 - 0x3f -- plane 1
      12'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      12'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      12'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      12'hF80: dout <= 8'b00111111; // 3968 :  63 - 0x3f -- Background 0xf8
      12'hF81: dout <= 8'b00111110; // 3969 :  62 - 0x3e
      12'hF82: dout <= 8'b00111100; // 3970 :  60 - 0x3c
      12'hF83: dout <= 8'b10111000; // 3971 : 184 - 0xb8
      12'hF84: dout <= 8'b01111000; // 3972 : 120 - 0x78
      12'hF85: dout <= 8'b01111000; // 3973 : 120 - 0x78
      12'hF86: dout <= 8'b01111110; // 3974 : 126 - 0x7e
      12'hF87: dout <= 8'b01111110; // 3975 : 126 - 0x7e
      12'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff -- plane 1
      12'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout <= 8'b11111101; // 3978 : 253 - 0xfd
      12'hF8B: dout <= 8'b11111000; // 3979 : 248 - 0xf8
      12'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      12'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      12'hF8E: dout <= 8'b11111110; // 3982 : 254 - 0xfe
      12'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      12'hF90: dout <= 8'b11111101; // 3984 : 253 - 0xfd -- Background 0xf9
      12'hF91: dout <= 8'b01111001; // 3985 : 121 - 0x79
      12'hF92: dout <= 8'b01111011; // 3986 : 123 - 0x7b
      12'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout <= 8'b11110011; // 3990 : 243 - 0xf3
      12'hF97: dout <= 8'b10000000; // 3991 : 128 - 0x80
      12'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff -- plane 1
      12'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout <= 8'b11111000; // 3999 : 248 - 0xf8
      12'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xfa
      12'hFA1: dout <= 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout <= 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout <= 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0 -- plane 1
      12'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b11000000; // 4014 : 192 - 0xc0
      12'hFAF: dout <= 8'b11110000; // 4015 : 240 - 0xf0
      12'hFB0: dout <= 8'b00010000; // 4016 :  16 - 0x10 -- Background 0xfb
      12'hFB1: dout <= 8'b10000100; // 4017 : 132 - 0x84
      12'hFB2: dout <= 8'b11100000; // 4018 : 224 - 0xe0
      12'hFB3: dout <= 8'b11000000; // 4019 : 192 - 0xc0
      12'hFB4: dout <= 8'b10000000; // 4020 : 128 - 0x80
      12'hFB5: dout <= 8'b10000000; // 4021 : 128 - 0x80
      12'hFB6: dout <= 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout <= 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout <= 8'b11111100; // 4024 : 252 - 0xfc -- plane 1
      12'hFB9: dout <= 8'b11111110; // 4025 : 254 - 0xfe
      12'hFBA: dout <= 8'b11101100; // 4026 : 236 - 0xec
      12'hFBB: dout <= 8'b11100000; // 4027 : 224 - 0xe0
      12'hFBC: dout <= 8'b11000000; // 4028 : 192 - 0xc0
      12'hFBD: dout <= 8'b11000000; // 4029 : 192 - 0xc0
      12'hFBE: dout <= 8'b10000000; // 4030 : 128 - 0x80
      12'hFBF: dout <= 8'b10000000; // 4031 : 128 - 0x80
      12'hFC0: dout <= 8'b00000000; // 4032 :   0 - 0x0 -- Background 0xfc
      12'hFC1: dout <= 8'b01001000; // 4033 :  72 - 0x48
      12'hFC2: dout <= 8'b00100000; // 4034 :  32 - 0x20
      12'hFC3: dout <= 8'b00000000; // 4035 :   0 - 0x0
      12'hFC4: dout <= 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout <= 8'b00000100; // 4037 :   4 - 0x4
      12'hFC6: dout <= 8'b00001110; // 4038 :  14 - 0xe
      12'hFC7: dout <= 8'b11111110; // 4039 : 254 - 0xfe
      12'hFC8: dout <= 8'b01110000; // 4040 : 112 - 0x70 -- plane 1
      12'hFC9: dout <= 8'b11111100; // 4041 : 252 - 0xfc
      12'hFCA: dout <= 8'b11111100; // 4042 : 252 - 0xfc
      12'hFCB: dout <= 8'b11111100; // 4043 : 252 - 0xfc
      12'hFCC: dout <= 8'b11111100; // 4044 : 252 - 0xfc
      12'hFCD: dout <= 8'b11111100; // 4045 : 252 - 0xfc
      12'hFCE: dout <= 8'b11111110; // 4046 : 254 - 0xfe
      12'hFCF: dout <= 8'b11111110; // 4047 : 254 - 0xfe
      12'hFD0: dout <= 8'b11111110; // 4048 : 254 - 0xfe -- Background 0xfd
      12'hFD1: dout <= 8'b11111100; // 4049 : 252 - 0xfc
      12'hFD2: dout <= 8'b11111100; // 4050 : 252 - 0xfc
      12'hFD3: dout <= 8'b11111000; // 4051 : 248 - 0xf8
      12'hFD4: dout <= 8'b11110000; // 4052 : 240 - 0xf0
      12'hFD5: dout <= 8'b11100000; // 4053 : 224 - 0xe0
      12'hFD6: dout <= 8'b10000000; // 4054 : 128 - 0x80
      12'hFD7: dout <= 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout <= 8'b11111110; // 4056 : 254 - 0xfe -- plane 1
      12'hFD9: dout <= 8'b11111100; // 4057 : 252 - 0xfc
      12'hFDA: dout <= 8'b11111100; // 4058 : 252 - 0xfc
      12'hFDB: dout <= 8'b11111000; // 4059 : 248 - 0xf8
      12'hFDC: dout <= 8'b11110000; // 4060 : 240 - 0xf0
      12'hFDD: dout <= 8'b11100000; // 4061 : 224 - 0xe0
      12'hFDE: dout <= 8'b10000000; // 4062 : 128 - 0x80
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b00001111; // 4064 :  15 - 0xf -- Background 0xfe
      12'hFE1: dout <= 8'b00000110; // 4065 :   6 - 0x6
      12'hFE2: dout <= 8'b00000110; // 4066 :   6 - 0x6
      12'hFE3: dout <= 8'b00000110; // 4067 :   6 - 0x6
      12'hFE4: dout <= 8'b00000110; // 4068 :   6 - 0x6
      12'hFE5: dout <= 8'b00000110; // 4069 :   6 - 0x6
      12'hFE6: dout <= 8'b00001111; // 4070 :  15 - 0xf
      12'hFE7: dout <= 8'b00000000; // 4071 :   0 - 0x0
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- plane 1
      12'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout <= 8'b00000000; // 4075 :   0 - 0x0
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b11110000; // 4080 : 240 - 0xf0 -- Background 0xff
      12'hFF1: dout <= 8'b01100000; // 4081 :  96 - 0x60
      12'hFF2: dout <= 8'b01100000; // 4082 :  96 - 0x60
      12'hFF3: dout <= 8'b01100110; // 4083 : 102 - 0x66
      12'hFF4: dout <= 8'b01100110; // 4084 : 102 - 0x66
      12'hFF5: dout <= 8'b01100000; // 4085 :  96 - 0x60
      12'hFF6: dout <= 8'b11110000; // 4086 : 240 - 0xf0
      12'hFF7: dout <= 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
