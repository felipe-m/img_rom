--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: smario_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_SMARIO_color0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_SMARIO_color0;

architecture BEHAVIORAL of ROM_PTABLE_SMARIO_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000011", --    0 -  0x0  :    3 - 0x3 -- Sprite 0x0
    "00001111", --    1 -  0x1  :   15 - 0xf
    "00011111", --    2 -  0x2  :   31 - 0x1f
    "00011111", --    3 -  0x3  :   31 - 0x1f
    "00011100", --    4 -  0x4  :   28 - 0x1c
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100110", --    6 -  0x6  :   38 - 0x26
    "01100110", --    7 -  0x7  :  102 - 0x66
    "11100000", --    8 -  0x8  :  224 - 0xe0 -- Sprite 0x1
    "11000000", --    9 -  0x9  :  192 - 0xc0
    "10000000", --   10 -  0xa  :  128 - 0x80
    "11111100", --   11 -  0xb  :  252 - 0xfc
    "10000000", --   12 -  0xc  :  128 - 0x80
    "11000000", --   13 -  0xd  :  192 - 0xc0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00100000", --   15 -  0xf  :   32 - 0x20
    "01100000", --   16 - 0x10  :   96 - 0x60 -- Sprite 0x2
    "01110000", --   17 - 0x11  :  112 - 0x70
    "00011000", --   18 - 0x12  :   24 - 0x18
    "00000111", --   19 - 0x13  :    7 - 0x7
    "00001111", --   20 - 0x14  :   15 - 0xf
    "00011111", --   21 - 0x15  :   31 - 0x1f
    "00111111", --   22 - 0x16  :   63 - 0x3f
    "01111111", --   23 - 0x17  :  127 - 0x7f
    "11111100", --   24 - 0x18  :  252 - 0xfc -- Sprite 0x3
    "01111100", --   25 - 0x19  :  124 - 0x7c
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "11100000", --   28 - 0x1c  :  224 - 0xe0
    "11110000", --   29 - 0x1d  :  240 - 0xf0
    "11111000", --   30 - 0x1e  :  248 - 0xf8
    "11111000", --   31 - 0x1f  :  248 - 0xf8
    "01111111", --   32 - 0x20  :  127 - 0x7f -- Sprite 0x4
    "01111111", --   33 - 0x21  :  127 - 0x7f
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "00000111", --   36 - 0x24  :    7 - 0x7
    "00000111", --   37 - 0x25  :    7 - 0x7
    "00001111", --   38 - 0x26  :   15 - 0xf
    "00001111", --   39 - 0x27  :   15 - 0xf
    "11111101", --   40 - 0x28  :  253 - 0xfd -- Sprite 0x5
    "11111110", --   41 - 0x29  :  254 - 0xfe
    "10110100", --   42 - 0x2a  :  180 - 0xb4
    "11111000", --   43 - 0x2b  :  248 - 0xf8
    "11111000", --   44 - 0x2c  :  248 - 0xf8
    "11111001", --   45 - 0x2d  :  249 - 0xf9
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111111", --   47 - 0x2f  :  255 - 0xff
    "00011111", --   48 - 0x30  :   31 - 0x1f -- Sprite 0x6
    "00111111", --   49 - 0x31  :   63 - 0x3f
    "11111111", --   50 - 0x32  :  255 - 0xff
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111100", --   52 - 0x34  :  252 - 0xfc
    "01110000", --   53 - 0x35  :  112 - 0x70
    "01110000", --   54 - 0x36  :  112 - 0x70
    "00111000", --   55 - 0x37  :   56 - 0x38
    "11111111", --   56 - 0x38  :  255 - 0xff -- Sprite 0x7
    "11111111", --   57 - 0x39  :  255 - 0xff
    "11111111", --   58 - 0x3a  :  255 - 0xff
    "00011111", --   59 - 0x3b  :   31 - 0x1f
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000001", --   66 - 0x42  :    1 - 0x1
    "00000111", --   67 - 0x43  :    7 - 0x7
    "00001111", --   68 - 0x44  :   15 - 0xf
    "00001111", --   69 - 0x45  :   15 - 0xf
    "00001110", --   70 - 0x46  :   14 - 0xe
    "00010010", --   71 - 0x47  :   18 - 0x12
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Sprite 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "11110000", --   74 - 0x4a  :  240 - 0xf0
    "11100000", --   75 - 0x4b  :  224 - 0xe0
    "11000000", --   76 - 0x4c  :  192 - 0xc0
    "11111110", --   77 - 0x4d  :  254 - 0xfe
    "01000000", --   78 - 0x4e  :   64 - 0x40
    "01100000", --   79 - 0x4f  :   96 - 0x60
    "00010011", --   80 - 0x50  :   19 - 0x13 -- Sprite 0xa
    "00110011", --   81 - 0x51  :   51 - 0x33
    "00110000", --   82 - 0x52  :   48 - 0x30
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00000100", --   84 - 0x54  :    4 - 0x4
    "00001111", --   85 - 0x55  :   15 - 0xf
    "00011111", --   86 - 0x56  :   31 - 0x1f
    "00011111", --   87 - 0x57  :   31 - 0x1f
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Sprite 0xb
    "00010000", --   89 - 0x59  :   16 - 0x10
    "01111110", --   90 - 0x5a  :  126 - 0x7e
    "00111110", --   91 - 0x5b  :   62 - 0x3e
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "11000000", --   94 - 0x5e  :  192 - 0xc0
    "11100000", --   95 - 0x5f  :  224 - 0xe0
    "00111111", --   96 - 0x60  :   63 - 0x3f -- Sprite 0xc
    "00111111", --   97 - 0x61  :   63 - 0x3f
    "00111111", --   98 - 0x62  :   63 - 0x3f
    "00011111", --   99 - 0x63  :   31 - 0x1f
    "00011111", --  100 - 0x64  :   31 - 0x1f
    "00011111", --  101 - 0x65  :   31 - 0x1f
    "00011111", --  102 - 0x66  :   31 - 0x1f
    "00011111", --  103 - 0x67  :   31 - 0x1f
    "11110000", --  104 - 0x68  :  240 - 0xf0 -- Sprite 0xd
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11110000", --  106 - 0x6a  :  240 - 0xf0
    "11111000", --  107 - 0x6b  :  248 - 0xf8
    "11111000", --  108 - 0x6c  :  248 - 0xf8
    "11111000", --  109 - 0x6d  :  248 - 0xf8
    "11111000", --  110 - 0x6e  :  248 - 0xf8
    "11111000", --  111 - 0x6f  :  248 - 0xf8
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0xe
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111111", --  114 - 0x72  :  255 - 0xff
    "11111110", --  115 - 0x73  :  254 - 0xfe
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "10000000", --  118 - 0x76  :  128 - 0x80
    "00000000", --  119 - 0x77  :    0 - 0x0
    "11111100", --  120 - 0x78  :  252 - 0xfc -- Sprite 0xf
    "11111100", --  121 - 0x79  :  252 - 0xfc
    "11111000", --  122 - 0x7a  :  248 - 0xf8
    "01111000", --  123 - 0x7b  :  120 - 0x78
    "01111000", --  124 - 0x7c  :  120 - 0x78
    "01111000", --  125 - 0x7d  :  120 - 0x78
    "01111110", --  126 - 0x7e  :  126 - 0x7e
    "01111110", --  127 - 0x7f  :  126 - 0x7e
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  129 - 0x81  :    3 - 0x3
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00011111", --  131 - 0x83  :   31 - 0x1f
    "00011111", --  132 - 0x84  :   31 - 0x1f
    "00011100", --  133 - 0x85  :   28 - 0x1c
    "00100100", --  134 - 0x86  :   36 - 0x24
    "00100110", --  135 - 0x87  :   38 - 0x26
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x11
    "11100000", --  137 - 0x89  :  224 - 0xe0
    "11000000", --  138 - 0x8a  :  192 - 0xc0
    "10000000", --  139 - 0x8b  :  128 - 0x80
    "11111100", --  140 - 0x8c  :  252 - 0xfc
    "10000000", --  141 - 0x8d  :  128 - 0x80
    "11000000", --  142 - 0x8e  :  192 - 0xc0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "01100110", --  144 - 0x90  :  102 - 0x66 -- Sprite 0x12
    "01100000", --  145 - 0x91  :   96 - 0x60
    "00110000", --  146 - 0x92  :   48 - 0x30
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00001111", --  148 - 0x94  :   15 - 0xf
    "00011111", --  149 - 0x95  :   31 - 0x1f
    "00111111", --  150 - 0x96  :   63 - 0x3f
    "00111111", --  151 - 0x97  :   63 - 0x3f
    "00100000", --  152 - 0x98  :   32 - 0x20 -- Sprite 0x13
    "11111100", --  153 - 0x99  :  252 - 0xfc
    "01111100", --  154 - 0x9a  :  124 - 0x7c
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "11100000", --  157 - 0x9d  :  224 - 0xe0
    "11100000", --  158 - 0x9e  :  224 - 0xe0
    "11110000", --  159 - 0x9f  :  240 - 0xf0
    "00111111", --  160 - 0xa0  :   63 - 0x3f -- Sprite 0x14
    "00111111", --  161 - 0xa1  :   63 - 0x3f
    "00111111", --  162 - 0xa2  :   63 - 0x3f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00111111", --  164 - 0xa4  :   63 - 0x3f
    "00111111", --  165 - 0xa5  :   63 - 0x3f
    "00111111", --  166 - 0xa6  :   63 - 0x3f
    "00011111", --  167 - 0xa7  :   31 - 0x1f
    "11110000", --  168 - 0xa8  :  240 - 0xf0 -- Sprite 0x15
    "10010000", --  169 - 0xa9  :  144 - 0x90
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00001000", --  171 - 0xab  :    8 - 0x8
    "00001100", --  172 - 0xac  :   12 - 0xc
    "00011100", --  173 - 0xad  :   28 - 0x1c
    "11111100", --  174 - 0xae  :  252 - 0xfc
    "11111000", --  175 - 0xaf  :  248 - 0xf8
    "00001111", --  176 - 0xb0  :   15 - 0xf -- Sprite 0x16
    "00001111", --  177 - 0xb1  :   15 - 0xf
    "00000111", --  178 - 0xb2  :    7 - 0x7
    "00000111", --  179 - 0xb3  :    7 - 0x7
    "00000111", --  180 - 0xb4  :    7 - 0x7
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00001111", --  182 - 0xb6  :   15 - 0xf
    "00000011", --  183 - 0xb7  :    3 - 0x3
    "11111000", --  184 - 0xb8  :  248 - 0xf8 -- Sprite 0x17
    "11110000", --  185 - 0xb9  :  240 - 0xf0
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "11110000", --  187 - 0xbb  :  240 - 0xf0
    "10110000", --  188 - 0xbc  :  176 - 0xb0
    "10000000", --  189 - 0xbd  :  128 - 0x80
    "11100000", --  190 - 0xbe  :  224 - 0xe0
    "11100000", --  191 - 0xbf  :  224 - 0xe0
    "00000011", --  192 - 0xc0  :    3 - 0x3 -- Sprite 0x18
    "00111111", --  193 - 0xc1  :   63 - 0x3f
    "01111111", --  194 - 0xc2  :  127 - 0x7f
    "00011001", --  195 - 0xc3  :   25 - 0x19
    "00001001", --  196 - 0xc4  :    9 - 0x9
    "00001001", --  197 - 0xc5  :    9 - 0x9
    "00101000", --  198 - 0xc6  :   40 - 0x28
    "01011100", --  199 - 0xc7  :   92 - 0x5c
    "11111000", --  200 - 0xc8  :  248 - 0xf8 -- Sprite 0x19
    "11100000", --  201 - 0xc9  :  224 - 0xe0
    "11100000", --  202 - 0xca  :  224 - 0xe0
    "11111100", --  203 - 0xcb  :  252 - 0xfc
    "00100110", --  204 - 0xcc  :   38 - 0x26
    "00110000", --  205 - 0xcd  :   48 - 0x30
    "10000000", --  206 - 0xce  :  128 - 0x80
    "00010000", --  207 - 0xcf  :   16 - 0x10
    "00111110", --  208 - 0xd0  :   62 - 0x3e -- Sprite 0x1a
    "00011110", --  209 - 0xd1  :   30 - 0x1e
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "00111000", --  211 - 0xd3  :   56 - 0x38
    "00110000", --  212 - 0xd4  :   48 - 0x30
    "00110000", --  213 - 0xd5  :   48 - 0x30
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00111010", --  215 - 0xd7  :   58 - 0x3a
    "01111000", --  216 - 0xd8  :  120 - 0x78 -- Sprite 0x1b
    "00011110", --  217 - 0xd9  :   30 - 0x1e
    "10000000", --  218 - 0xda  :  128 - 0x80
    "11111110", --  219 - 0xdb  :  254 - 0xfe
    "01111110", --  220 - 0xdc  :  126 - 0x7e
    "01111110", --  221 - 0xdd  :  126 - 0x7e
    "01111111", --  222 - 0xde  :  127 - 0x7f
    "01111111", --  223 - 0xdf  :  127 - 0x7f
    "00111100", --  224 - 0xe0  :   60 - 0x3c -- Sprite 0x1c
    "00111111", --  225 - 0xe1  :   63 - 0x3f
    "00011111", --  226 - 0xe2  :   31 - 0x1f
    "00001111", --  227 - 0xe3  :   15 - 0xf
    "00000111", --  228 - 0xe4  :    7 - 0x7
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00100001", --  230 - 0xe6  :   33 - 0x21
    "00100000", --  231 - 0xe7  :   32 - 0x20
    "11111111", --  232 - 0xe8  :  255 - 0xff -- Sprite 0x1d
    "11111111", --  233 - 0xe9  :  255 - 0xff
    "11111111", --  234 - 0xea  :  255 - 0xff
    "11111110", --  235 - 0xeb  :  254 - 0xfe
    "11111110", --  236 - 0xec  :  254 - 0xfe
    "11111110", --  237 - 0xed  :  254 - 0xfe
    "11111100", --  238 - 0xee  :  252 - 0xfc
    "01110000", --  239 - 0xef  :  112 - 0x70
    "00001111", --  240 - 0xf0  :   15 - 0xf -- Sprite 0x1e
    "10011111", --  241 - 0xf1  :  159 - 0x9f
    "11001111", --  242 - 0xf2  :  207 - 0xcf
    "11111111", --  243 - 0xf3  :  255 - 0xff
    "01111111", --  244 - 0xf4  :  127 - 0x7f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00011110", --  246 - 0xf6  :   30 - 0x1e
    "00001110", --  247 - 0xf7  :   14 - 0xe
    "00100000", --  248 - 0xf8  :   32 - 0x20 -- Sprite 0x1f
    "11000000", --  249 - 0xf9  :  192 - 0xc0
    "10000000", --  250 - 0xfa  :  128 - 0x80
    "10000000", --  251 - 0xfb  :  128 - 0x80
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000011", --  258 - 0x102  :    3 - 0x3
    "00001111", --  259 - 0x103  :   15 - 0xf
    "00011111", --  260 - 0x104  :   31 - 0x1f
    "00011111", --  261 - 0x105  :   31 - 0x1f
    "00011100", --  262 - 0x106  :   28 - 0x1c
    "00100100", --  263 - 0x107  :   36 - 0x24
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000100", --  265 - 0x109  :    4 - 0x4
    "11100110", --  266 - 0x10a  :  230 - 0xe6
    "11100000", --  267 - 0x10b  :  224 - 0xe0
    "11111111", --  268 - 0x10c  :  255 - 0xff
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "10001111", --  270 - 0x10e  :  143 - 0x8f
    "10000011", --  271 - 0x10f  :  131 - 0x83
    "00100110", --  272 - 0x110  :   38 - 0x26 -- Sprite 0x22
    "00100110", --  273 - 0x111  :   38 - 0x26
    "01100000", --  274 - 0x112  :   96 - 0x60
    "01111000", --  275 - 0x113  :  120 - 0x78
    "00011000", --  276 - 0x114  :   24 - 0x18
    "00001111", --  277 - 0x115  :   15 - 0xf
    "01111111", --  278 - 0x116  :  127 - 0x7f
    "11111111", --  279 - 0x117  :  255 - 0xff
    "00000001", --  280 - 0x118  :    1 - 0x1 -- Sprite 0x23
    "00100001", --  281 - 0x119  :   33 - 0x21
    "11111110", --  282 - 0x11a  :  254 - 0xfe
    "01111010", --  283 - 0x11b  :  122 - 0x7a
    "00000110", --  284 - 0x11c  :    6 - 0x6
    "11111110", --  285 - 0x11d  :  254 - 0xfe
    "11111100", --  286 - 0x11e  :  252 - 0xfc
    "11111100", --  287 - 0x11f  :  252 - 0xfc
    "11111111", --  288 - 0x120  :  255 - 0xff -- Sprite 0x24
    "11001111", --  289 - 0x121  :  207 - 0xcf
    "10000111", --  290 - 0x122  :  135 - 0x87
    "00000111", --  291 - 0x123  :    7 - 0x7
    "00000111", --  292 - 0x124  :    7 - 0x7
    "00001111", --  293 - 0x125  :   15 - 0xf
    "00011111", --  294 - 0x126  :   31 - 0x1f
    "00011111", --  295 - 0x127  :   31 - 0x1f
    "11111000", --  296 - 0x128  :  248 - 0xf8 -- Sprite 0x25
    "11111000", --  297 - 0x129  :  248 - 0xf8
    "11110000", --  298 - 0x12a  :  240 - 0xf0
    "10111000", --  299 - 0x12b  :  184 - 0xb8
    "11111000", --  300 - 0x12c  :  248 - 0xf8
    "11111001", --  301 - 0x12d  :  249 - 0xf9
    "11111011", --  302 - 0x12e  :  251 - 0xfb
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "00011111", --  304 - 0x130  :   31 - 0x1f -- Sprite 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111110", --  309 - 0x135  :  254 - 0xfe
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "10000000", --  311 - 0x137  :  128 - 0x80
    "11111111", --  312 - 0x138  :  255 - 0xff -- Sprite 0x27
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "00111111", --  315 - 0x13b  :   63 - 0x3f
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00010011", --  320 - 0x140  :   19 - 0x13 -- Sprite 0x28
    "00110011", --  321 - 0x141  :   51 - 0x33
    "00110000", --  322 - 0x142  :   48 - 0x30
    "00011000", --  323 - 0x143  :   24 - 0x18
    "00000100", --  324 - 0x144  :    4 - 0x4
    "00001111", --  325 - 0x145  :   15 - 0xf
    "00011111", --  326 - 0x146  :   31 - 0x1f
    "00011111", --  327 - 0x147  :   31 - 0x1f
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Sprite 0x29
    "00010000", --  329 - 0x149  :   16 - 0x10
    "01111110", --  330 - 0x14a  :  126 - 0x7e
    "00110000", --  331 - 0x14b  :   48 - 0x30
    "11100000", --  332 - 0x14c  :  224 - 0xe0
    "11110000", --  333 - 0x14d  :  240 - 0xf0
    "11110000", --  334 - 0x14e  :  240 - 0xf0
    "11100000", --  335 - 0x14f  :  224 - 0xe0
    "00011111", --  336 - 0x150  :   31 - 0x1f -- Sprite 0x2a
    "00011111", --  337 - 0x151  :   31 - 0x1f
    "00001111", --  338 - 0x152  :   15 - 0xf
    "00001111", --  339 - 0x153  :   15 - 0xf
    "00001111", --  340 - 0x154  :   15 - 0xf
    "00011111", --  341 - 0x155  :   31 - 0x1f
    "00011111", --  342 - 0x156  :   31 - 0x1f
    "00011111", --  343 - 0x157  :   31 - 0x1f
    "11110000", --  344 - 0x158  :  240 - 0xf0 -- Sprite 0x2b
    "11110000", --  345 - 0x159  :  240 - 0xf0
    "11111000", --  346 - 0x15a  :  248 - 0xf8
    "11111000", --  347 - 0x15b  :  248 - 0xf8
    "10111000", --  348 - 0x15c  :  184 - 0xb8
    "11111000", --  349 - 0x15d  :  248 - 0xf8
    "11111000", --  350 - 0x15e  :  248 - 0xf8
    "11111000", --  351 - 0x15f  :  248 - 0xf8
    "00111111", --  352 - 0x160  :   63 - 0x3f -- Sprite 0x2c
    "11111111", --  353 - 0x161  :  255 - 0xff
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111111", --  355 - 0x163  :  255 - 0xff
    "11110110", --  356 - 0x164  :  246 - 0xf6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "10000100", --  358 - 0x166  :  132 - 0x84
    "00000000", --  359 - 0x167  :    0 - 0x0
    "11110000", --  360 - 0x168  :  240 - 0xf0 -- Sprite 0x2d
    "11100000", --  361 - 0x169  :  224 - 0xe0
    "10000000", --  362 - 0x16a  :  128 - 0x80
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00011111", --  368 - 0x170  :   31 - 0x1f -- Sprite 0x2e
    "00011111", --  369 - 0x171  :   31 - 0x1f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111111", --  371 - 0x173  :   63 - 0x3f
    "00011111", --  372 - 0x174  :   31 - 0x1f
    "00001111", --  373 - 0x175  :   15 - 0xf
    "00001111", --  374 - 0x176  :   15 - 0xf
    "00011111", --  375 - 0x177  :   31 - 0x1f
    "11110000", --  376 - 0x178  :  240 - 0xf0 -- Sprite 0x2f
    "11110000", --  377 - 0x179  :  240 - 0xf0
    "11111000", --  378 - 0x17a  :  248 - 0xf8
    "11111000", --  379 - 0x17b  :  248 - 0xf8
    "10111000", --  380 - 0x17c  :  184 - 0xb8
    "11111000", --  381 - 0x17d  :  248 - 0xf8
    "11111000", --  382 - 0x17e  :  248 - 0xf8
    "11110000", --  383 - 0x17f  :  240 - 0xf0
    "11100000", --  384 - 0x180  :  224 - 0xe0 -- Sprite 0x30
    "11110000", --  385 - 0x181  :  240 - 0xf0
    "11110000", --  386 - 0x182  :  240 - 0xf0
    "11110000", --  387 - 0x183  :  240 - 0xf0
    "11110000", --  388 - 0x184  :  240 - 0xf0
    "11110000", --  389 - 0x185  :  240 - 0xf0
    "11111000", --  390 - 0x186  :  248 - 0xf8
    "11110000", --  391 - 0x187  :  240 - 0xf0
    "00011111", --  392 - 0x188  :   31 - 0x1f -- Sprite 0x31
    "00011111", --  393 - 0x189  :   31 - 0x1f
    "00011111", --  394 - 0x18a  :   31 - 0x1f
    "00111111", --  395 - 0x18b  :   63 - 0x3f
    "00111110", --  396 - 0x18c  :   62 - 0x3e
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00111000", --  398 - 0x18e  :   56 - 0x38
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "00000011", --  401 - 0x191  :    3 - 0x3
    "00000111", --  402 - 0x192  :    7 - 0x7
    "00000111", --  403 - 0x193  :    7 - 0x7
    "00001010", --  404 - 0x194  :   10 - 0xa
    "00001011", --  405 - 0x195  :   11 - 0xb
    "00001100", --  406 - 0x196  :   12 - 0xc
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Sprite 0x33
    "11100000", --  409 - 0x199  :  224 - 0xe0
    "11111100", --  410 - 0x19a  :  252 - 0xfc
    "00100000", --  411 - 0x19b  :   32 - 0x20
    "00100000", --  412 - 0x19c  :   32 - 0x20
    "00010000", --  413 - 0x19d  :   16 - 0x10
    "00111100", --  414 - 0x19e  :   60 - 0x3c
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000111", --  416 - 0x1a0  :    7 - 0x7 -- Sprite 0x34
    "00000111", --  417 - 0x1a1  :    7 - 0x7
    "00000111", --  418 - 0x1a2  :    7 - 0x7
    "00011111", --  419 - 0x1a3  :   31 - 0x1f
    "00011111", --  420 - 0x1a4  :   31 - 0x1f
    "00111110", --  421 - 0x1a5  :   62 - 0x3e
    "00100001", --  422 - 0x1a6  :   33 - 0x21
    "00000001", --  423 - 0x1a7  :    1 - 0x1
    "11100000", --  424 - 0x1a8  :  224 - 0xe0 -- Sprite 0x35
    "11100000", --  425 - 0x1a9  :  224 - 0xe0
    "11100000", --  426 - 0x1aa  :  224 - 0xe0
    "11110000", --  427 - 0x1ab  :  240 - 0xf0
    "11110000", --  428 - 0x1ac  :  240 - 0xf0
    "11100000", --  429 - 0x1ad  :  224 - 0xe0
    "11000000", --  430 - 0x1ae  :  192 - 0xc0
    "11100000", --  431 - 0x1af  :  224 - 0xe0
    "00000111", --  432 - 0x1b0  :    7 - 0x7 -- Sprite 0x36
    "00001111", --  433 - 0x1b1  :   15 - 0xf
    "00001110", --  434 - 0x1b2  :   14 - 0xe
    "00010100", --  435 - 0x1b3  :   20 - 0x14
    "00010110", --  436 - 0x1b4  :   22 - 0x16
    "00011000", --  437 - 0x1b5  :   24 - 0x18
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00111111", --  439 - 0x1b7  :   63 - 0x3f
    "11000000", --  440 - 0x1b8  :  192 - 0xc0 -- Sprite 0x37
    "11111000", --  441 - 0x1b9  :  248 - 0xf8
    "01000000", --  442 - 0x1ba  :   64 - 0x40
    "01000000", --  443 - 0x1bb  :   64 - 0x40
    "00100000", --  444 - 0x1bc  :   32 - 0x20
    "01111000", --  445 - 0x1bd  :  120 - 0x78
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "11000000", --  447 - 0x1bf  :  192 - 0xc0
    "00111111", --  448 - 0x1c0  :   63 - 0x3f -- Sprite 0x38
    "00001110", --  449 - 0x1c1  :   14 - 0xe
    "00001111", --  450 - 0x1c2  :   15 - 0xf
    "00011111", --  451 - 0x1c3  :   31 - 0x1f
    "00111111", --  452 - 0x1c4  :   63 - 0x3f
    "01111100", --  453 - 0x1c5  :  124 - 0x7c
    "01110000", --  454 - 0x1c6  :  112 - 0x70
    "00111000", --  455 - 0x1c7  :   56 - 0x38
    "11110000", --  456 - 0x1c8  :  240 - 0xf0 -- Sprite 0x39
    "11111000", --  457 - 0x1c9  :  248 - 0xf8
    "11100100", --  458 - 0x1ca  :  228 - 0xe4
    "11111100", --  459 - 0x1cb  :  252 - 0xfc
    "11111100", --  460 - 0x1cc  :  252 - 0xfc
    "01111100", --  461 - 0x1cd  :  124 - 0x7c
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000111", --  464 - 0x1d0  :    7 - 0x7 -- Sprite 0x3a
    "00001111", --  465 - 0x1d1  :   15 - 0xf
    "00001110", --  466 - 0x1d2  :   14 - 0xe
    "00010100", --  467 - 0x1d3  :   20 - 0x14
    "00010110", --  468 - 0x1d4  :   22 - 0x16
    "00011000", --  469 - 0x1d5  :   24 - 0x18
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00001111", --  471 - 0x1d7  :   15 - 0xf
    "00011111", --  472 - 0x1d8  :   31 - 0x1f -- Sprite 0x3b
    "00011111", --  473 - 0x1d9  :   31 - 0x1f
    "00011111", --  474 - 0x1da  :   31 - 0x1f
    "00011100", --  475 - 0x1db  :   28 - 0x1c
    "00001100", --  476 - 0x1dc  :   12 - 0xc
    "00000111", --  477 - 0x1dd  :    7 - 0x7
    "00000111", --  478 - 0x1de  :    7 - 0x7
    "00000111", --  479 - 0x1df  :    7 - 0x7
    "11100000", --  480 - 0x1e0  :  224 - 0xe0 -- Sprite 0x3c
    "01100000", --  481 - 0x1e1  :   96 - 0x60
    "11110000", --  482 - 0x1e2  :  240 - 0xf0
    "01110000", --  483 - 0x1e3  :  112 - 0x70
    "11100000", --  484 - 0x1e4  :  224 - 0xe0
    "11100000", --  485 - 0x1e5  :  224 - 0xe0
    "11110000", --  486 - 0x1e6  :  240 - 0xf0
    "10000000", --  487 - 0x1e7  :  128 - 0x80
    "00000111", --  488 - 0x1e8  :    7 - 0x7 -- Sprite 0x3d
    "00011111", --  489 - 0x1e9  :   31 - 0x1f
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "00010010", --  491 - 0x1eb  :   18 - 0x12
    "00010011", --  492 - 0x1ec  :   19 - 0x13
    "00001000", --  493 - 0x1ed  :    8 - 0x8
    "00011111", --  494 - 0x1ee  :   31 - 0x1f
    "00110001", --  495 - 0x1ef  :   49 - 0x31
    "11000000", --  496 - 0x1f0  :  192 - 0xc0 -- Sprite 0x3e
    "11110000", --  497 - 0x1f1  :  240 - 0xf0
    "01000000", --  498 - 0x1f2  :   64 - 0x40
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00110000", --  500 - 0x1f4  :   48 - 0x30
    "00011000", --  501 - 0x1f5  :   24 - 0x18
    "11000000", --  502 - 0x1f6  :  192 - 0xc0
    "11111000", --  503 - 0x1f7  :  248 - 0xf8
    "00110001", --  504 - 0x1f8  :   49 - 0x31 -- Sprite 0x3f
    "00111001", --  505 - 0x1f9  :   57 - 0x39
    "00011111", --  506 - 0x1fa  :   31 - 0x1f
    "00011111", --  507 - 0x1fb  :   31 - 0x1f
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "01011111", --  509 - 0x1fd  :   95 - 0x5f
    "01111110", --  510 - 0x1fe  :  126 - 0x7e
    "00111100", --  511 - 0x1ff  :   60 - 0x3c
    "11111000", --  512 - 0x200  :  248 - 0xf8 -- Sprite 0x40
    "11111000", --  513 - 0x201  :  248 - 0xf8
    "11110000", --  514 - 0x202  :  240 - 0xf0
    "11100000", --  515 - 0x203  :  224 - 0xe0
    "11100000", --  516 - 0x204  :  224 - 0xe0
    "11000000", --  517 - 0x205  :  192 - 0xc0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Sprite 0x41
    "11100000", --  521 - 0x209  :  224 - 0xe0
    "11111100", --  522 - 0x20a  :  252 - 0xfc
    "00100111", --  523 - 0x20b  :   39 - 0x27
    "00100111", --  524 - 0x20c  :   39 - 0x27
    "00010001", --  525 - 0x20d  :   17 - 0x11
    "00111110", --  526 - 0x20e  :   62 - 0x3e
    "00000100", --  527 - 0x20f  :    4 - 0x4
    "00111111", --  528 - 0x210  :   63 - 0x3f -- Sprite 0x42
    "01111111", --  529 - 0x211  :  127 - 0x7f
    "00111111", --  530 - 0x212  :   63 - 0x3f
    "00001111", --  531 - 0x213  :   15 - 0xf
    "00011111", --  532 - 0x214  :   31 - 0x1f
    "00111111", --  533 - 0x215  :   63 - 0x3f
    "01111111", --  534 - 0x216  :  127 - 0x7f
    "01001111", --  535 - 0x217  :   79 - 0x4f
    "11111000", --  536 - 0x218  :  248 - 0xf8 -- Sprite 0x43
    "11111001", --  537 - 0x219  :  249 - 0xf9
    "11111001", --  538 - 0x21a  :  249 - 0xf9
    "10110111", --  539 - 0x21b  :  183 - 0xb7
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11100000", --  542 - 0x21e  :  224 - 0xe0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000111", --  544 - 0x220  :    7 - 0x7 -- Sprite 0x44
    "00000111", --  545 - 0x221  :    7 - 0x7
    "00001111", --  546 - 0x222  :   15 - 0xf
    "00111111", --  547 - 0x223  :   63 - 0x3f
    "00111111", --  548 - 0x224  :   63 - 0x3f
    "00111111", --  549 - 0x225  :   63 - 0x3f
    "00100110", --  550 - 0x226  :   38 - 0x26
    "00000100", --  551 - 0x227  :    4 - 0x4
    "11110000", --  552 - 0x228  :  240 - 0xf0 -- Sprite 0x45
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11110000", --  554 - 0x22a  :  240 - 0xf0
    "11100000", --  555 - 0x22b  :  224 - 0xe0
    "11000000", --  556 - 0x22c  :  192 - 0xc0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000111", --  560 - 0x230  :    7 - 0x7 -- Sprite 0x46
    "00000111", --  561 - 0x231  :    7 - 0x7
    "00001111", --  562 - 0x232  :   15 - 0xf
    "00011111", --  563 - 0x233  :   31 - 0x1f
    "00111111", --  564 - 0x234  :   63 - 0x3f
    "00001111", --  565 - 0x235  :   15 - 0xf
    "00011100", --  566 - 0x236  :   28 - 0x1c
    "00011000", --  567 - 0x237  :   24 - 0x18
    "11100000", --  568 - 0x238  :  224 - 0xe0 -- Sprite 0x47
    "11100000", --  569 - 0x239  :  224 - 0xe0
    "11100000", --  570 - 0x23a  :  224 - 0xe0
    "11100000", --  571 - 0x23b  :  224 - 0xe0
    "11000000", --  572 - 0x23c  :  192 - 0xc0
    "10000000", --  573 - 0x23d  :  128 - 0x80
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000111", --  576 - 0x240  :    7 - 0x7 -- Sprite 0x48
    "00001111", --  577 - 0x241  :   15 - 0xf
    "00011111", --  578 - 0x242  :   31 - 0x1f
    "00001111", --  579 - 0x243  :   15 - 0xf
    "00111111", --  580 - 0x244  :   63 - 0x3f
    "00001111", --  581 - 0x245  :   15 - 0xf
    "00011100", --  582 - 0x246  :   28 - 0x1c
    "00011000", --  583 - 0x247  :   24 - 0x18
    "11100000", --  584 - 0x248  :  224 - 0xe0 -- Sprite 0x49
    "11100000", --  585 - 0x249  :  224 - 0xe0
    "11100000", --  586 - 0x24a  :  224 - 0xe0
    "01000000", --  587 - 0x24b  :   64 - 0x40
    "11000000", --  588 - 0x24c  :  192 - 0xc0
    "10000000", --  589 - 0x24d  :  128 - 0x80
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "01111111", --  592 - 0x250  :  127 - 0x7f -- Sprite 0x4a
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111011", --  595 - 0x253  :  251 - 0xfb
    "00001111", --  596 - 0x254  :   15 - 0xf
    "00001111", --  597 - 0x255  :   15 - 0xf
    "00001111", --  598 - 0x256  :   15 - 0xf
    "00011111", --  599 - 0x257  :   31 - 0x1f
    "00111111", --  600 - 0x258  :   63 - 0x3f -- Sprite 0x4b
    "01111110", --  601 - 0x259  :  126 - 0x7e
    "01111100", --  602 - 0x25a  :  124 - 0x7c
    "01111100", --  603 - 0x25b  :  124 - 0x7c
    "00111100", --  604 - 0x25c  :   60 - 0x3c
    "00111100", --  605 - 0x25d  :   60 - 0x3c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "01100000", --  608 - 0x260  :   96 - 0x60 -- Sprite 0x4c
    "01110000", --  609 - 0x261  :  112 - 0x70
    "00011000", --  610 - 0x262  :   24 - 0x18
    "00001000", --  611 - 0x263  :    8 - 0x8
    "00001111", --  612 - 0x264  :   15 - 0xf
    "00011111", --  613 - 0x265  :   31 - 0x1f
    "00111111", --  614 - 0x266  :   63 - 0x3f
    "01111111", --  615 - 0x267  :  127 - 0x7f
    "11111100", --  616 - 0x268  :  252 - 0xfc -- Sprite 0x4d
    "01111100", --  617 - 0x269  :  124 - 0x7c
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00100000", --  619 - 0x26b  :   32 - 0x20
    "11110000", --  620 - 0x26c  :  240 - 0xf0
    "11111000", --  621 - 0x26d  :  248 - 0xf8
    "11111100", --  622 - 0x26e  :  252 - 0xfc
    "11111110", --  623 - 0x26f  :  254 - 0xfe
    "00001011", --  624 - 0x270  :   11 - 0xb -- Sprite 0x4e
    "00001111", --  625 - 0x271  :   15 - 0xf
    "00011111", --  626 - 0x272  :   31 - 0x1f
    "00011110", --  627 - 0x273  :   30 - 0x1e
    "00111100", --  628 - 0x274  :   60 - 0x3c
    "00111100", --  629 - 0x275  :   60 - 0x3c
    "00111100", --  630 - 0x276  :   60 - 0x3c
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "00011111", --  632 - 0x278  :   31 - 0x1f -- Sprite 0x4f
    "00111111", --  633 - 0x279  :   63 - 0x3f
    "00001101", --  634 - 0x27a  :   13 - 0xd
    "00000111", --  635 - 0x27b  :    7 - 0x7
    "00001111", --  636 - 0x27c  :   15 - 0xf
    "00001110", --  637 - 0x27d  :   14 - 0xe
    "00011100", --  638 - 0x27e  :   28 - 0x1c
    "00111100", --  639 - 0x27f  :   60 - 0x3c
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00000111", --  649 - 0x289  :    7 - 0x7
    "00011111", --  650 - 0x28a  :   31 - 0x1f
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "00000111", --  652 - 0x28c  :    7 - 0x7
    "00011111", --  653 - 0x28d  :   31 - 0x1f
    "00001111", --  654 - 0x28e  :   15 - 0xf
    "00000110", --  655 - 0x28f  :    6 - 0x6
    "00111111", --  656 - 0x290  :   63 - 0x3f -- Sprite 0x52
    "11111111", --  657 - 0x291  :  255 - 0xff
    "11111111", --  658 - 0x292  :  255 - 0xff
    "11111111", --  659 - 0x293  :  255 - 0xff
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111111", --  661 - 0x295  :  255 - 0xff
    "11111011", --  662 - 0x296  :  251 - 0xfb
    "01110110", --  663 - 0x297  :  118 - 0x76
    "00100000", --  664 - 0x298  :   32 - 0x20 -- Sprite 0x53
    "11111000", --  665 - 0x299  :  248 - 0xf8
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11000011", --  667 - 0x29b  :  195 - 0xc3
    "11111101", --  668 - 0x29c  :  253 - 0xfd
    "11111110", --  669 - 0x29d  :  254 - 0xfe
    "11110000", --  670 - 0x29e  :  240 - 0xf0
    "01000000", --  671 - 0x29f  :   64 - 0x40
    "01000000", --  672 - 0x2a0  :   64 - 0x40 -- Sprite 0x54
    "11100000", --  673 - 0x2a1  :  224 - 0xe0
    "01000000", --  674 - 0x2a2  :   64 - 0x40
    "01000000", --  675 - 0x2a3  :   64 - 0x40
    "01000001", --  676 - 0x2a4  :   65 - 0x41
    "01000001", --  677 - 0x2a5  :   65 - 0x41
    "01001111", --  678 - 0x2a6  :   79 - 0x4f
    "01000111", --  679 - 0x2a7  :   71 - 0x47
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "11100000", --  686 - 0x2ae  :  224 - 0xe0
    "11000000", --  687 - 0x2af  :  192 - 0xc0
    "01000011", --  688 - 0x2b0  :   67 - 0x43 -- Sprite 0x56
    "01000110", --  689 - 0x2b1  :   70 - 0x46
    "01000100", --  690 - 0x2b2  :   68 - 0x44
    "01000000", --  691 - 0x2b3  :   64 - 0x40
    "01000000", --  692 - 0x2b4  :   64 - 0x40
    "01000000", --  693 - 0x2b5  :   64 - 0x40
    "01000000", --  694 - 0x2b6  :   64 - 0x40
    "01000000", --  695 - 0x2b7  :   64 - 0x40
    "10000000", --  696 - 0x2b8  :  128 - 0x80 -- Sprite 0x57
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "01000000", --  698 - 0x2ba  :   64 - 0x40
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00110001", --  704 - 0x2c0  :   49 - 0x31 -- Sprite 0x58
    "00110000", --  705 - 0x2c1  :   48 - 0x30
    "00111000", --  706 - 0x2c2  :   56 - 0x38
    "01111100", --  707 - 0x2c3  :  124 - 0x7c
    "01111111", --  708 - 0x2c4  :  127 - 0x7f
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11111111", --  710 - 0x2c6  :  255 - 0xff
    "11111011", --  711 - 0x2c7  :  251 - 0xfb
    "00010000", --  712 - 0x2c8  :   16 - 0x10 -- Sprite 0x59
    "01111110", --  713 - 0x2c9  :  126 - 0x7e
    "00111110", --  714 - 0x2ca  :   62 - 0x3e
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00011110", --  716 - 0x2cc  :   30 - 0x1e
    "11111110", --  717 - 0x2cd  :  254 - 0xfe
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "11111111", --  720 - 0x2d0  :  255 - 0xff -- Sprite 0x5a
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11100011", --  722 - 0x2d2  :  227 - 0xe3
    "11000011", --  723 - 0x2d3  :  195 - 0xc3
    "10000111", --  724 - 0x2d4  :  135 - 0x87
    "01001000", --  725 - 0x2d5  :   72 - 0x48
    "00111100", --  726 - 0x2d6  :   60 - 0x3c
    "11111100", --  727 - 0x2d7  :  252 - 0xfc
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11000011", --  730 - 0x2da  :  195 - 0xc3
    "10000011", --  731 - 0x2db  :  131 - 0x83
    "10000011", --  732 - 0x2dc  :  131 - 0x83
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00011111", --  736 - 0x2e0  :   31 - 0x1f -- Sprite 0x5c
    "00011111", --  737 - 0x2e1  :   31 - 0x1f
    "00001111", --  738 - 0x2e2  :   15 - 0xf
    "00000111", --  739 - 0x2e3  :    7 - 0x7
    "00000001", --  740 - 0x2e4  :    1 - 0x1
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "11110000", --  744 - 0x2e8  :  240 - 0xf0 -- Sprite 0x5d
    "11111011", --  745 - 0x2e9  :  251 - 0xfb
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11111110", --  748 - 0x2ec  :  254 - 0xfe
    "00111110", --  749 - 0x2ed  :   62 - 0x3e
    "00001100", --  750 - 0x2ee  :   12 - 0xc
    "00000100", --  751 - 0x2ef  :    4 - 0x4
    "00011111", --  752 - 0x2f0  :   31 - 0x1f -- Sprite 0x5e
    "00011111", --  753 - 0x2f1  :   31 - 0x1f
    "00001111", --  754 - 0x2f2  :   15 - 0xf
    "00001111", --  755 - 0x2f3  :   15 - 0xf
    "00000111", --  756 - 0x2f4  :    7 - 0x7
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "11111011", --  760 - 0x2f8  :  251 - 0xfb -- Sprite 0x5f
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111111", --  763 - 0x2fb  :  255 - 0xff
    "11111111", --  764 - 0x2fc  :  255 - 0xff
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00011000", --  769 - 0x301  :   24 - 0x18
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "01111110", --  771 - 0x303  :  126 - 0x7e
    "01101110", --  772 - 0x304  :  110 - 0x6e
    "11011111", --  773 - 0x305  :  223 - 0xdf
    "11011111", --  774 - 0x306  :  223 - 0xdf
    "11011111", --  775 - 0x307  :  223 - 0xdf
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "00011000", --  777 - 0x309  :   24 - 0x18
    "00011000", --  778 - 0x30a  :   24 - 0x18
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "00111100", --  780 - 0x30c  :   60 - 0x3c
    "00111100", --  781 - 0x30d  :   60 - 0x3c
    "00111100", --  782 - 0x30e  :   60 - 0x3c
    "00011100", --  783 - 0x30f  :   28 - 0x1c
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x62
    "00001000", --  785 - 0x311  :    8 - 0x8
    "00001000", --  786 - 0x312  :    8 - 0x8
    "00001000", --  787 - 0x313  :    8 - 0x8
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00001000", --  789 - 0x315  :    8 - 0x8
    "00001000", --  790 - 0x316  :    8 - 0x8
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Sprite 0x63
    "00001000", --  793 - 0x319  :    8 - 0x8
    "00001000", --  794 - 0x31a  :    8 - 0x8
    "00000100", --  795 - 0x31b  :    4 - 0x4
    "00000100", --  796 - 0x31c  :    4 - 0x4
    "00000100", --  797 - 0x31d  :    4 - 0x4
    "00000100", --  798 - 0x31e  :    4 - 0x4
    "00000100", --  799 - 0x31f  :    4 - 0x4
    "00111100", --  800 - 0x320  :   60 - 0x3c -- Sprite 0x64
    "01111110", --  801 - 0x321  :  126 - 0x7e
    "01110111", --  802 - 0x322  :  119 - 0x77
    "11111011", --  803 - 0x323  :  251 - 0xfb
    "10011111", --  804 - 0x324  :  159 - 0x9f
    "01011111", --  805 - 0x325  :   95 - 0x5f
    "10001110", --  806 - 0x326  :  142 - 0x8e
    "00100000", --  807 - 0x327  :   32 - 0x20
    "01011100", --  808 - 0x328  :   92 - 0x5c -- Sprite 0x65
    "00101110", --  809 - 0x329  :   46 - 0x2e
    "10001111", --  810 - 0x32a  :  143 - 0x8f
    "00111111", --  811 - 0x32b  :   63 - 0x3f
    "01111011", --  812 - 0x32c  :  123 - 0x7b
    "01110111", --  813 - 0x32d  :  119 - 0x77
    "01111110", --  814 - 0x32e  :  126 - 0x7e
    "00111100", --  815 - 0x32f  :   60 - 0x3c
    "00010011", --  816 - 0x330  :   19 - 0x13 -- Sprite 0x66
    "01001111", --  817 - 0x331  :   79 - 0x4f
    "00111111", --  818 - 0x332  :   63 - 0x3f
    "10111111", --  819 - 0x333  :  191 - 0xbf
    "00111111", --  820 - 0x334  :   63 - 0x3f
    "01111010", --  821 - 0x335  :  122 - 0x7a
    "11111000", --  822 - 0x336  :  248 - 0xf8
    "11111000", --  823 - 0x337  :  248 - 0xf8
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Sprite 0x67
    "00001000", --  825 - 0x339  :    8 - 0x8
    "00000101", --  826 - 0x33a  :    5 - 0x5
    "00001111", --  827 - 0x33b  :   15 - 0xf
    "00101111", --  828 - 0x33c  :   47 - 0x2f
    "00011101", --  829 - 0x33d  :   29 - 0x1d
    "00011100", --  830 - 0x33e  :   28 - 0x1c
    "00111100", --  831 - 0x33f  :   60 - 0x3c
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000010", --  836 - 0x344  :    2 - 0x2
    "00001011", --  837 - 0x345  :   11 - 0xb
    "00000111", --  838 - 0x346  :    7 - 0x7
    "00001111", --  839 - 0x347  :   15 - 0xf
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00001000", --  845 - 0x34d  :    8 - 0x8
    "00000100", --  846 - 0x34e  :    4 - 0x4
    "00000100", --  847 - 0x34f  :    4 - 0x4
    "00000010", --  848 - 0x350  :    2 - 0x2 -- Sprite 0x6a
    "00000010", --  849 - 0x351  :    2 - 0x2
    "00000010", --  850 - 0x352  :    2 - 0x2
    "00000101", --  851 - 0x353  :    5 - 0x5
    "01110001", --  852 - 0x354  :  113 - 0x71
    "01111111", --  853 - 0x355  :  127 - 0x7f
    "01111111", --  854 - 0x356  :  127 - 0x7f
    "01111111", --  855 - 0x357  :  127 - 0x7f
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000100", --  863 - 0x35f  :    4 - 0x4
    "00000010", --  864 - 0x360  :    2 - 0x2 -- Sprite 0x6c
    "00000010", --  865 - 0x361  :    2 - 0x2
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000001", --  867 - 0x363  :    1 - 0x1
    "00010011", --  868 - 0x364  :   19 - 0x13
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "01111111", --  870 - 0x366  :  127 - 0x7f
    "01111111", --  871 - 0x367  :  127 - 0x7f
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "01000000", --  873 - 0x369  :   64 - 0x40
    "01100000", --  874 - 0x36a  :   96 - 0x60
    "01110000", --  875 - 0x36b  :  112 - 0x70
    "01110011", --  876 - 0x36c  :  115 - 0x73
    "00100111", --  877 - 0x36d  :   39 - 0x27
    "00001111", --  878 - 0x36e  :   15 - 0xf
    "00011111", --  879 - 0x36f  :   31 - 0x1f
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000011", --  884 - 0x374  :    3 - 0x3
    "00000111", --  885 - 0x375  :    7 - 0x7
    "00001111", --  886 - 0x376  :   15 - 0xf
    "00011111", --  887 - 0x377  :   31 - 0x1f
    "01111111", --  888 - 0x378  :  127 - 0x7f -- Sprite 0x6f
    "01111111", --  889 - 0x379  :  127 - 0x7f
    "00111111", --  890 - 0x37a  :   63 - 0x3f
    "00111111", --  891 - 0x37b  :   63 - 0x3f
    "00011111", --  892 - 0x37c  :   31 - 0x1f
    "00011111", --  893 - 0x37d  :   31 - 0x1f
    "00001111", --  894 - 0x37e  :   15 - 0xf
    "00000111", --  895 - 0x37f  :    7 - 0x7
    "00000011", --  896 - 0x380  :    3 - 0x3 -- Sprite 0x70
    "00000111", --  897 - 0x381  :    7 - 0x7
    "00001111", --  898 - 0x382  :   15 - 0xf
    "00011111", --  899 - 0x383  :   31 - 0x1f
    "00111111", --  900 - 0x384  :   63 - 0x3f
    "01110111", --  901 - 0x385  :  119 - 0x77
    "01110111", --  902 - 0x386  :  119 - 0x77
    "11110101", --  903 - 0x387  :  245 - 0xf5
    "11000000", --  904 - 0x388  :  192 - 0xc0 -- Sprite 0x71
    "11100000", --  905 - 0x389  :  224 - 0xe0
    "11110000", --  906 - 0x38a  :  240 - 0xf0
    "11111000", --  907 - 0x38b  :  248 - 0xf8
    "11111100", --  908 - 0x38c  :  252 - 0xfc
    "11101110", --  909 - 0x38d  :  238 - 0xee
    "11101110", --  910 - 0x38e  :  238 - 0xee
    "10101111", --  911 - 0x38f  :  175 - 0xaf
    "11110001", --  912 - 0x390  :  241 - 0xf1 -- Sprite 0x72
    "11111111", --  913 - 0x391  :  255 - 0xff
    "01111000", --  914 - 0x392  :  120 - 0x78
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00011000", --  917 - 0x395  :   24 - 0x18
    "00011100", --  918 - 0x396  :   28 - 0x1c
    "00001110", --  919 - 0x397  :   14 - 0xe
    "10001111", --  920 - 0x398  :  143 - 0x8f -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "00011110", --  922 - 0x39a  :   30 - 0x1e
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00001100", --  924 - 0x39c  :   12 - 0xc
    "00111110", --  925 - 0x39d  :   62 - 0x3e
    "01111110", --  926 - 0x39e  :  126 - 0x7e
    "01111100", --  927 - 0x39f  :  124 - 0x7c
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Sprite 0x75
    "00000010", --  937 - 0x3a9  :    2 - 0x2
    "01000001", --  938 - 0x3aa  :   65 - 0x41
    "01000001", --  939 - 0x3ab  :   65 - 0x41
    "01100001", --  940 - 0x3ac  :   97 - 0x61
    "00110011", --  941 - 0x3ad  :   51 - 0x33
    "00000110", --  942 - 0x3ae  :    6 - 0x6
    "00111100", --  943 - 0x3af  :   60 - 0x3c
    "00000011", --  944 - 0x3b0  :    3 - 0x3 -- Sprite 0x76
    "00000111", --  945 - 0x3b1  :    7 - 0x7
    "00001111", --  946 - 0x3b2  :   15 - 0xf
    "00011111", --  947 - 0x3b3  :   31 - 0x1f
    "00111111", --  948 - 0x3b4  :   63 - 0x3f
    "01111111", --  949 - 0x3b5  :  127 - 0x7f
    "01111111", --  950 - 0x3b6  :  127 - 0x7f
    "11111111", --  951 - 0x3b7  :  255 - 0xff
    "11000000", --  952 - 0x3b8  :  192 - 0xc0 -- Sprite 0x77
    "11100000", --  953 - 0x3b9  :  224 - 0xe0
    "11110000", --  954 - 0x3ba  :  240 - 0xf0
    "11111000", --  955 - 0x3bb  :  248 - 0xf8
    "11111100", --  956 - 0x3bc  :  252 - 0xfc
    "11111110", --  957 - 0x3bd  :  254 - 0xfe
    "11111110", --  958 - 0x3be  :  254 - 0xfe
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Sprite 0x78
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "01111000", --  963 - 0x3c3  :  120 - 0x78
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Sprite 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "00011110", --  971 - 0x3cb  :   30 - 0x1e
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00100000", --  973 - 0x3cd  :   32 - 0x20
    "00100000", --  974 - 0x3ce  :   32 - 0x20
    "01000000", --  975 - 0x3cf  :   64 - 0x40
    "00010110", --  976 - 0x3d0  :   22 - 0x16 -- Sprite 0x7a
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00111111", --  978 - 0x3d2  :   63 - 0x3f
    "01111111", --  979 - 0x3d3  :  127 - 0x7f
    "00111101", --  980 - 0x3d4  :   61 - 0x3d
    "00011101", --  981 - 0x3d5  :   29 - 0x1d
    "00111111", --  982 - 0x3d6  :   63 - 0x3f
    "00011111", --  983 - 0x3d7  :   31 - 0x1f
    "10000000", --  984 - 0x3d8  :  128 - 0x80 -- Sprite 0x7b
    "10000000", --  985 - 0x3d9  :  128 - 0x80
    "11000000", --  986 - 0x3da  :  192 - 0xc0
    "11100000", --  987 - 0x3db  :  224 - 0xe0
    "11110000", --  988 - 0x3dc  :  240 - 0xf0
    "11110000", --  989 - 0x3dd  :  240 - 0xf0
    "11110000", --  990 - 0x3de  :  240 - 0xf0
    "11111000", --  991 - 0x3df  :  248 - 0xf8
    "00111100", --  992 - 0x3e0  :   60 - 0x3c -- Sprite 0x7c
    "11111010", --  993 - 0x3e1  :  250 - 0xfa
    "10110001", --  994 - 0x3e2  :  177 - 0xb1
    "01110010", --  995 - 0x3e3  :  114 - 0x72
    "11110010", --  996 - 0x3e4  :  242 - 0xf2
    "11011011", --  997 - 0x3e5  :  219 - 0xdb
    "11011111", --  998 - 0x3e6  :  223 - 0xdf
    "01011111", --  999 - 0x3e7  :   95 - 0x5f
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000001", -- 1003 - 0x3eb  :    1 - 0x1
    "00000001", -- 1004 - 0x3ec  :    1 - 0x1
    "00000001", -- 1005 - 0x3ed  :    1 - 0x1
    "00000110", -- 1006 - 0x3ee  :    6 - 0x6
    "00011110", -- 1007 - 0x3ef  :   30 - 0x1e
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- Sprite 0x7f
    "01111100", -- 1017 - 0x3f9  :  124 - 0x7c
    "11010110", -- 1018 - 0x3fa  :  214 - 0xd6
    "10010010", -- 1019 - 0x3fb  :  146 - 0x92
    "10111010", -- 1020 - 0x3fc  :  186 - 0xba
    "11101110", -- 1021 - 0x3fd  :  238 - 0xee
    "11111110", -- 1022 - 0x3fe  :  254 - 0xfe
    "00111000", -- 1023 - 0x3ff  :   56 - 0x38
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x80
    "00010101", -- 1025 - 0x401  :   21 - 0x15
    "00111111", -- 1026 - 0x402  :   63 - 0x3f
    "01100010", -- 1027 - 0x403  :   98 - 0x62
    "01011111", -- 1028 - 0x404  :   95 - 0x5f
    "11111111", -- 1029 - 0x405  :  255 - 0xff
    "10011111", -- 1030 - 0x406  :  159 - 0x9f
    "01111101", -- 1031 - 0x407  :  125 - 0x7d
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Sprite 0x81
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00101111", -- 1040 - 0x410  :   47 - 0x2f -- Sprite 0x82
    "00011110", -- 1041 - 0x411  :   30 - 0x1e
    "00101111", -- 1042 - 0x412  :   47 - 0x2f
    "00101111", -- 1043 - 0x413  :   47 - 0x2f
    "00101111", -- 1044 - 0x414  :   47 - 0x2f
    "00010101", -- 1045 - 0x415  :   21 - 0x15
    "00001101", -- 1046 - 0x416  :   13 - 0xd
    "00001110", -- 1047 - 0x417  :   14 - 0xe
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00011100", -- 1056 - 0x420  :   28 - 0x1c -- Sprite 0x84
    "00111110", -- 1057 - 0x421  :   62 - 0x3e
    "01111111", -- 1058 - 0x422  :  127 - 0x7f
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111110", -- 1061 - 0x425  :  254 - 0xfe
    "01111100", -- 1062 - 0x426  :  124 - 0x7c
    "00111000", -- 1063 - 0x427  :   56 - 0x38
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Sprite 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111111", -- 1067 - 0x42b  :  255 - 0xff
    "11111111", -- 1068 - 0x42c  :  255 - 0xff
    "11111111", -- 1069 - 0x42d  :  255 - 0xff
    "11111111", -- 1070 - 0x42e  :  255 - 0xff
    "11111111", -- 1071 - 0x42f  :  255 - 0xff
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11111111", -- 1078 - 0x436  :  255 - 0xff
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "01111111", -- 1080 - 0x438  :  127 - 0x7f -- Sprite 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "11111111", -- 1087 - 0x43f  :  255 - 0xff
    "01101000", -- 1088 - 0x440  :  104 - 0x68 -- Sprite 0x88
    "01001110", -- 1089 - 0x441  :   78 - 0x4e
    "11100000", -- 1090 - 0x442  :  224 - 0xe0
    "11100000", -- 1091 - 0x443  :  224 - 0xe0
    "11100000", -- 1092 - 0x444  :  224 - 0xe0
    "11110000", -- 1093 - 0x445  :  240 - 0xf0
    "11111000", -- 1094 - 0x446  :  248 - 0xf8
    "11111100", -- 1095 - 0x447  :  252 - 0xfc
    "00111111", -- 1096 - 0x448  :   63 - 0x3f -- Sprite 0x89
    "01011100", -- 1097 - 0x449  :   92 - 0x5c
    "00111001", -- 1098 - 0x44a  :   57 - 0x39
    "00111011", -- 1099 - 0x44b  :   59 - 0x3b
    "10111011", -- 1100 - 0x44c  :  187 - 0xbb
    "11111001", -- 1101 - 0x44d  :  249 - 0xf9
    "11111100", -- 1102 - 0x44e  :  252 - 0xfc
    "11111110", -- 1103 - 0x44f  :  254 - 0xfe
    "11000000", -- 1104 - 0x450  :  192 - 0xc0 -- Sprite 0x8a
    "11110000", -- 1105 - 0x451  :  240 - 0xf0
    "11110000", -- 1106 - 0x452  :  240 - 0xf0
    "11110000", -- 1107 - 0x453  :  240 - 0xf0
    "11110000", -- 1108 - 0x454  :  240 - 0xf0
    "11100000", -- 1109 - 0x455  :  224 - 0xe0
    "11000000", -- 1110 - 0x456  :  192 - 0xc0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "11111110", -- 1112 - 0x458  :  254 - 0xfe -- Sprite 0x8b
    "11111100", -- 1113 - 0x459  :  252 - 0xfc
    "01100001", -- 1114 - 0x45a  :   97 - 0x61
    "00001111", -- 1115 - 0x45b  :   15 - 0xf
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "11111110", -- 1117 - 0x45d  :  254 - 0xfe
    "11110000", -- 1118 - 0x45e  :  240 - 0xf0
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "01101110", -- 1120 - 0x460  :  110 - 0x6e -- Sprite 0x8c
    "01000000", -- 1121 - 0x461  :   64 - 0x40
    "11100000", -- 1122 - 0x462  :  224 - 0xe0
    "11100000", -- 1123 - 0x463  :  224 - 0xe0
    "11100000", -- 1124 - 0x464  :  224 - 0xe0
    "11100000", -- 1125 - 0x465  :  224 - 0xe0
    "11100000", -- 1126 - 0x466  :  224 - 0xe0
    "11000000", -- 1127 - 0x467  :  192 - 0xc0
    "00000001", -- 1128 - 0x468  :    1 - 0x1 -- Sprite 0x8d
    "00000001", -- 1129 - 0x469  :    1 - 0x1
    "00000011", -- 1130 - 0x46a  :    3 - 0x3
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000111", -- 1132 - 0x46c  :    7 - 0x7
    "01111111", -- 1133 - 0x46d  :  127 - 0x7f
    "01111111", -- 1134 - 0x46e  :  127 - 0x7f
    "00111111", -- 1135 - 0x46f  :   63 - 0x3f
    "00000110", -- 1136 - 0x470  :    6 - 0x6 -- Sprite 0x8e
    "00000111", -- 1137 - 0x471  :    7 - 0x7
    "00111111", -- 1138 - 0x472  :   63 - 0x3f
    "00111100", -- 1139 - 0x473  :   60 - 0x3c
    "00011001", -- 1140 - 0x474  :   25 - 0x19
    "01111011", -- 1141 - 0x475  :  123 - 0x7b
    "01111111", -- 1142 - 0x476  :  127 - 0x7f
    "00111111", -- 1143 - 0x477  :   63 - 0x3f
    "00111111", -- 1144 - 0x478  :   63 - 0x3f -- Sprite 0x8f
    "01111111", -- 1145 - 0x479  :  127 - 0x7f
    "01111111", -- 1146 - 0x47a  :  127 - 0x7f
    "00011111", -- 1147 - 0x47b  :   31 - 0x1f
    "00111111", -- 1148 - 0x47c  :   63 - 0x3f
    "00111111", -- 1149 - 0x47d  :   63 - 0x3f
    "00000111", -- 1150 - 0x47e  :    7 - 0x7
    "00000110", -- 1151 - 0x47f  :    6 - 0x6
    "00000011", -- 1152 - 0x480  :    3 - 0x3 -- Sprite 0x90
    "00000111", -- 1153 - 0x481  :    7 - 0x7
    "00001111", -- 1154 - 0x482  :   15 - 0xf
    "00001111", -- 1155 - 0x483  :   15 - 0xf
    "00001111", -- 1156 - 0x484  :   15 - 0xf
    "00001111", -- 1157 - 0x485  :   15 - 0xf
    "00000111", -- 1158 - 0x486  :    7 - 0x7
    "00000011", -- 1159 - 0x487  :    3 - 0x3
    "11111000", -- 1160 - 0x488  :  248 - 0xf8 -- Sprite 0x91
    "11111000", -- 1161 - 0x489  :  248 - 0xf8
    "11111000", -- 1162 - 0x48a  :  248 - 0xf8
    "10100000", -- 1163 - 0x48b  :  160 - 0xa0
    "11100001", -- 1164 - 0x48c  :  225 - 0xe1
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "00001111", -- 1168 - 0x490  :   15 - 0xf -- Sprite 0x92
    "00001111", -- 1169 - 0x491  :   15 - 0xf
    "00001111", -- 1170 - 0x492  :   15 - 0xf
    "00011111", -- 1171 - 0x493  :   31 - 0x1f
    "00011111", -- 1172 - 0x494  :   31 - 0x1f
    "00011111", -- 1173 - 0x495  :   31 - 0x1f
    "00001111", -- 1174 - 0x496  :   15 - 0xf
    "00000111", -- 1175 - 0x497  :    7 - 0x7
    "11100000", -- 1176 - 0x498  :  224 - 0xe0 -- Sprite 0x93
    "11111000", -- 1177 - 0x499  :  248 - 0xf8
    "11111000", -- 1178 - 0x49a  :  248 - 0xf8
    "11111000", -- 1179 - 0x49b  :  248 - 0xf8
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111110", -- 1181 - 0x49d  :  254 - 0xfe
    "11110000", -- 1182 - 0x49e  :  240 - 0xf0
    "11000000", -- 1183 - 0x49f  :  192 - 0xc0
    "00000001", -- 1184 - 0x4a0  :    1 - 0x1 -- Sprite 0x94
    "00001111", -- 1185 - 0x4a1  :   15 - 0xf
    "00001111", -- 1186 - 0x4a2  :   15 - 0xf
    "00011111", -- 1187 - 0x4a3  :   31 - 0x1f
    "00111001", -- 1188 - 0x4a4  :   57 - 0x39
    "00110011", -- 1189 - 0x4a5  :   51 - 0x33
    "00110111", -- 1190 - 0x4a6  :   55 - 0x37
    "01111111", -- 1191 - 0x4a7  :  127 - 0x7f
    "01111111", -- 1192 - 0x4a8  :  127 - 0x7f -- Sprite 0x95
    "00111111", -- 1193 - 0x4a9  :   63 - 0x3f
    "00111111", -- 1194 - 0x4aa  :   63 - 0x3f
    "00111111", -- 1195 - 0x4ab  :   63 - 0x3f
    "00011111", -- 1196 - 0x4ac  :   31 - 0x1f
    "00001111", -- 1197 - 0x4ad  :   15 - 0xf
    "00001111", -- 1198 - 0x4ae  :   15 - 0xf
    "00000001", -- 1199 - 0x4af  :    1 - 0x1
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000011", -- 1202 - 0x4b2  :    3 - 0x3
    "00000011", -- 1203 - 0x4b3  :    3 - 0x3
    "01000111", -- 1204 - 0x4b4  :   71 - 0x47
    "01100111", -- 1205 - 0x4b5  :  103 - 0x67
    "01110111", -- 1206 - 0x4b6  :  119 - 0x77
    "01110111", -- 1207 - 0x4b7  :  119 - 0x77
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- Sprite 0x97
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "10001000", -- 1212 - 0x4bc  :  136 - 0x88
    "10011000", -- 1213 - 0x4bd  :  152 - 0x98
    "11111000", -- 1214 - 0x4be  :  248 - 0xf8
    "11110000", -- 1215 - 0x4bf  :  240 - 0xf0
    "01111110", -- 1216 - 0x4c0  :  126 - 0x7e -- Sprite 0x98
    "01111111", -- 1217 - 0x4c1  :  127 - 0x7f
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "00011111", -- 1219 - 0x4c3  :   31 - 0x1f
    "00000111", -- 1220 - 0x4c4  :    7 - 0x7
    "00110000", -- 1221 - 0x4c5  :   48 - 0x30
    "00011100", -- 1222 - 0x4c6  :   28 - 0x1c
    "00001100", -- 1223 - 0x4c7  :   12 - 0xc
    "01111110", -- 1224 - 0x4c8  :  126 - 0x7e -- Sprite 0x99
    "00111000", -- 1225 - 0x4c9  :   56 - 0x38
    "11110110", -- 1226 - 0x4ca  :  246 - 0xf6
    "11101101", -- 1227 - 0x4cb  :  237 - 0xed
    "11011111", -- 1228 - 0x4cc  :  223 - 0xdf
    "00111000", -- 1229 - 0x4cd  :   56 - 0x38
    "01110000", -- 1230 - 0x4ce  :  112 - 0x70
    "01100000", -- 1231 - 0x4cf  :   96 - 0x60
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000011", -- 1235 - 0x4d3  :    3 - 0x3
    "00000011", -- 1236 - 0x4d4  :    3 - 0x3
    "01000111", -- 1237 - 0x4d5  :   71 - 0x47
    "01100111", -- 1238 - 0x4d6  :  103 - 0x67
    "01110111", -- 1239 - 0x4d7  :  119 - 0x77
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- Sprite 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "10001000", -- 1245 - 0x4dd  :  136 - 0x88
    "10011000", -- 1246 - 0x4de  :  152 - 0x98
    "11111000", -- 1247 - 0x4df  :  248 - 0xf8
    "01110111", -- 1248 - 0x4e0  :  119 - 0x77 -- Sprite 0x9c
    "01111110", -- 1249 - 0x4e1  :  126 - 0x7e
    "01111111", -- 1250 - 0x4e2  :  127 - 0x7f
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "00011111", -- 1252 - 0x4e4  :   31 - 0x1f
    "00000111", -- 1253 - 0x4e5  :    7 - 0x7
    "01110000", -- 1254 - 0x4e6  :  112 - 0x70
    "11110000", -- 1255 - 0x4e7  :  240 - 0xf0
    "11110000", -- 1256 - 0x4e8  :  240 - 0xf0 -- Sprite 0x9d
    "01111110", -- 1257 - 0x4e9  :  126 - 0x7e
    "00111000", -- 1258 - 0x4ea  :   56 - 0x38
    "11110110", -- 1259 - 0x4eb  :  246 - 0xf6
    "11101101", -- 1260 - 0x4ec  :  237 - 0xed
    "11011111", -- 1261 - 0x4ed  :  223 - 0xdf
    "00111000", -- 1262 - 0x4ee  :   56 - 0x38
    "00111100", -- 1263 - 0x4ef  :   60 - 0x3c
    "00000011", -- 1264 - 0x4f0  :    3 - 0x3 -- Sprite 0x9e
    "00000111", -- 1265 - 0x4f1  :    7 - 0x7
    "00001010", -- 1266 - 0x4f2  :   10 - 0xa
    "00011010", -- 1267 - 0x4f3  :   26 - 0x1a
    "00011100", -- 1268 - 0x4f4  :   28 - 0x1c
    "00011110", -- 1269 - 0x4f5  :   30 - 0x1e
    "00001011", -- 1270 - 0x4f6  :   11 - 0xb
    "00001000", -- 1271 - 0x4f7  :    8 - 0x8
    "00011100", -- 1272 - 0x4f8  :   28 - 0x1c -- Sprite 0x9f
    "00111111", -- 1273 - 0x4f9  :   63 - 0x3f
    "00111111", -- 1274 - 0x4fa  :   63 - 0x3f
    "00111101", -- 1275 - 0x4fb  :   61 - 0x3d
    "00111111", -- 1276 - 0x4fc  :   63 - 0x3f
    "00011111", -- 1277 - 0x4fd  :   31 - 0x1f
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0xa0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000100", -- 1282 - 0x502  :    4 - 0x4
    "01001100", -- 1283 - 0x503  :   76 - 0x4c
    "01001110", -- 1284 - 0x504  :   78 - 0x4e
    "01001110", -- 1285 - 0x505  :   78 - 0x4e
    "01000110", -- 1286 - 0x506  :   70 - 0x46
    "01101111", -- 1287 - 0x507  :  111 - 0x6f
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- Sprite 0xa1
    "00011111", -- 1289 - 0x509  :   31 - 0x1f
    "00111111", -- 1290 - 0x50a  :   63 - 0x3f
    "00111111", -- 1291 - 0x50b  :   63 - 0x3f
    "01001111", -- 1292 - 0x50c  :   79 - 0x4f
    "01011111", -- 1293 - 0x50d  :   95 - 0x5f
    "01111111", -- 1294 - 0x50e  :  127 - 0x7f
    "01111111", -- 1295 - 0x50f  :  127 - 0x7f
    "01111111", -- 1296 - 0x510  :  127 - 0x7f -- Sprite 0xa2
    "01100111", -- 1297 - 0x511  :  103 - 0x67
    "10100011", -- 1298 - 0x512  :  163 - 0xa3
    "10110000", -- 1299 - 0x513  :  176 - 0xb0
    "11011000", -- 1300 - 0x514  :  216 - 0xd8
    "11011110", -- 1301 - 0x515  :  222 - 0xde
    "11011100", -- 1302 - 0x516  :  220 - 0xdc
    "11001000", -- 1303 - 0x517  :  200 - 0xc8
    "01111111", -- 1304 - 0x518  :  127 - 0x7f -- Sprite 0xa3
    "01111111", -- 1305 - 0x519  :  127 - 0x7f
    "01111111", -- 1306 - 0x51a  :  127 - 0x7f
    "00011111", -- 1307 - 0x51b  :   31 - 0x1f
    "01000111", -- 1308 - 0x51c  :   71 - 0x47
    "01110000", -- 1309 - 0x51d  :  112 - 0x70
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "00111001", -- 1311 - 0x51f  :   57 - 0x39
    "11101000", -- 1312 - 0x520  :  232 - 0xe8 -- Sprite 0xa4
    "11101000", -- 1313 - 0x521  :  232 - 0xe8
    "11100000", -- 1314 - 0x522  :  224 - 0xe0
    "11000000", -- 1315 - 0x523  :  192 - 0xc0
    "00010000", -- 1316 - 0x524  :   16 - 0x10
    "01110000", -- 1317 - 0x525  :  112 - 0x70
    "11100000", -- 1318 - 0x526  :  224 - 0xe0
    "11000000", -- 1319 - 0x527  :  192 - 0xc0
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00100000", -- 1323 - 0x52b  :   32 - 0x20
    "01100110", -- 1324 - 0x52c  :  102 - 0x66
    "01100110", -- 1325 - 0x52d  :  102 - 0x66
    "01100110", -- 1326 - 0x52e  :  102 - 0x66
    "01100010", -- 1327 - 0x52f  :   98 - 0x62
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00011111", -- 1330 - 0x532  :   31 - 0x1f
    "00111111", -- 1331 - 0x533  :   63 - 0x3f
    "01111111", -- 1332 - 0x534  :  127 - 0x7f
    "01001111", -- 1333 - 0x535  :   79 - 0x4f
    "01011111", -- 1334 - 0x536  :   95 - 0x5f
    "01111111", -- 1335 - 0x537  :  127 - 0x7f
    "01110111", -- 1336 - 0x538  :  119 - 0x77 -- Sprite 0xa7
    "01111111", -- 1337 - 0x539  :  127 - 0x7f
    "00111111", -- 1338 - 0x53a  :   63 - 0x3f
    "10110111", -- 1339 - 0x53b  :  183 - 0xb7
    "10110011", -- 1340 - 0x53c  :  179 - 0xb3
    "11011011", -- 1341 - 0x53d  :  219 - 0xdb
    "11011010", -- 1342 - 0x53e  :  218 - 0xda
    "11011000", -- 1343 - 0x53f  :  216 - 0xd8
    "01111111", -- 1344 - 0x540  :  127 - 0x7f -- Sprite 0xa8
    "01111111", -- 1345 - 0x541  :  127 - 0x7f
    "01111111", -- 1346 - 0x542  :  127 - 0x7f
    "01111111", -- 1347 - 0x543  :  127 - 0x7f
    "00011111", -- 1348 - 0x544  :   31 - 0x1f
    "00000111", -- 1349 - 0x545  :    7 - 0x7
    "01110000", -- 1350 - 0x546  :  112 - 0x70
    "11110000", -- 1351 - 0x547  :  240 - 0xf0
    "11001100", -- 1352 - 0x548  :  204 - 0xcc -- Sprite 0xa9
    "11101000", -- 1353 - 0x549  :  232 - 0xe8
    "11101000", -- 1354 - 0x54a  :  232 - 0xe8
    "11100000", -- 1355 - 0x54b  :  224 - 0xe0
    "11000000", -- 1356 - 0x54c  :  192 - 0xc0
    "00011000", -- 1357 - 0x54d  :   24 - 0x18
    "01111100", -- 1358 - 0x54e  :  124 - 0x7c
    "00111110", -- 1359 - 0x54f  :   62 - 0x3e
    "00000011", -- 1360 - 0x550  :    3 - 0x3 -- Sprite 0xaa
    "00001111", -- 1361 - 0x551  :   15 - 0xf
    "00011111", -- 1362 - 0x552  :   31 - 0x1f
    "00111111", -- 1363 - 0x553  :   63 - 0x3f
    "00111011", -- 1364 - 0x554  :   59 - 0x3b
    "00111111", -- 1365 - 0x555  :   63 - 0x3f
    "01111111", -- 1366 - 0x556  :  127 - 0x7f
    "01111111", -- 1367 - 0x557  :  127 - 0x7f
    "10000000", -- 1368 - 0x558  :  128 - 0x80 -- Sprite 0xab
    "11110000", -- 1369 - 0x559  :  240 - 0xf0
    "11111000", -- 1370 - 0x55a  :  248 - 0xf8
    "11111100", -- 1371 - 0x55b  :  252 - 0xfc
    "11111110", -- 1372 - 0x55c  :  254 - 0xfe
    "11111110", -- 1373 - 0x55d  :  254 - 0xfe
    "11111111", -- 1374 - 0x55e  :  255 - 0xff
    "11111110", -- 1375 - 0x55f  :  254 - 0xfe
    "01111111", -- 1376 - 0x560  :  127 - 0x7f -- Sprite 0xac
    "01111111", -- 1377 - 0x561  :  127 - 0x7f
    "01111111", -- 1378 - 0x562  :  127 - 0x7f
    "01111111", -- 1379 - 0x563  :  127 - 0x7f
    "11111111", -- 1380 - 0x564  :  255 - 0xff
    "00001111", -- 1381 - 0x565  :   15 - 0xf
    "00000011", -- 1382 - 0x566  :    3 - 0x3
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "11111110", -- 1384 - 0x568  :  254 - 0xfe -- Sprite 0xad
    "11111011", -- 1385 - 0x569  :  251 - 0xfb
    "11111111", -- 1386 - 0x56a  :  255 - 0xff
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "11110110", -- 1388 - 0x56c  :  246 - 0xf6
    "11100000", -- 1389 - 0x56d  :  224 - 0xe0
    "11000000", -- 1390 - 0x56e  :  192 - 0xc0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00001111", -- 1394 - 0x572  :   15 - 0xf
    "00011111", -- 1395 - 0x573  :   31 - 0x1f
    "00111111", -- 1396 - 0x574  :   63 - 0x3f
    "00111011", -- 1397 - 0x575  :   59 - 0x3b
    "00111111", -- 1398 - 0x576  :   63 - 0x3f
    "01111111", -- 1399 - 0x577  :  127 - 0x7f
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "11000000", -- 1401 - 0x579  :  192 - 0xc0
    "11110000", -- 1402 - 0x57a  :  240 - 0xf0
    "11111000", -- 1403 - 0x57b  :  248 - 0xf8
    "11111100", -- 1404 - 0x57c  :  252 - 0xfc
    "11111110", -- 1405 - 0x57d  :  254 - 0xfe
    "11111110", -- 1406 - 0x57e  :  254 - 0xfe
    "11111111", -- 1407 - 0x57f  :  255 - 0xff
    "01111111", -- 1408 - 0x580  :  127 - 0x7f -- Sprite 0xb0
    "01111111", -- 1409 - 0x581  :  127 - 0x7f
    "01111111", -- 1410 - 0x582  :  127 - 0x7f
    "01111111", -- 1411 - 0x583  :  127 - 0x7f
    "01111111", -- 1412 - 0x584  :  127 - 0x7f
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "00001111", -- 1414 - 0x586  :   15 - 0xf
    "00000011", -- 1415 - 0x587  :    3 - 0x3
    "11111110", -- 1416 - 0x588  :  254 - 0xfe -- Sprite 0xb1
    "11111110", -- 1417 - 0x589  :  254 - 0xfe
    "11111011", -- 1418 - 0x58a  :  251 - 0xfb
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11110110", -- 1421 - 0x58d  :  246 - 0xf6
    "11100000", -- 1422 - 0x58e  :  224 - 0xe0
    "11000000", -- 1423 - 0x58f  :  192 - 0xc0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0xb2
    "00000001", -- 1425 - 0x591  :    1 - 0x1
    "00000001", -- 1426 - 0x592  :    1 - 0x1
    "00000001", -- 1427 - 0x593  :    1 - 0x1
    "00000001", -- 1428 - 0x594  :    1 - 0x1
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00001000", -- 1431 - 0x597  :    8 - 0x8
    "01111000", -- 1432 - 0x598  :  120 - 0x78 -- Sprite 0xb3
    "11110000", -- 1433 - 0x599  :  240 - 0xf0
    "11111000", -- 1434 - 0x59a  :  248 - 0xf8
    "11100100", -- 1435 - 0x59b  :  228 - 0xe4
    "11000000", -- 1436 - 0x59c  :  192 - 0xc0
    "11001010", -- 1437 - 0x59d  :  202 - 0xca
    "11001010", -- 1438 - 0x59e  :  202 - 0xca
    "11000000", -- 1439 - 0x59f  :  192 - 0xc0
    "00001111", -- 1440 - 0x5a0  :   15 - 0xf -- Sprite 0xb4
    "00011111", -- 1441 - 0x5a1  :   31 - 0x1f
    "10011111", -- 1442 - 0x5a2  :  159 - 0x9f
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "01111111", -- 1445 - 0x5a5  :  127 - 0x7f
    "01110100", -- 1446 - 0x5a6  :  116 - 0x74
    "00100000", -- 1447 - 0x5a7  :   32 - 0x20
    "11100100", -- 1448 - 0x5a8  :  228 - 0xe4 -- Sprite 0xb5
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111110", -- 1450 - 0x5aa  :  254 - 0xfe
    "11111100", -- 1451 - 0x5ab  :  252 - 0xfc
    "10011100", -- 1452 - 0x5ac  :  156 - 0x9c
    "00011110", -- 1453 - 0x5ad  :   30 - 0x1e
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "00000001", -- 1457 - 0x5b1  :    1 - 0x1
    "00000011", -- 1458 - 0x5b2  :    3 - 0x3
    "00000011", -- 1459 - 0x5b3  :    3 - 0x3
    "00000111", -- 1460 - 0x5b4  :    7 - 0x7
    "00000011", -- 1461 - 0x5b5  :    3 - 0x3
    "00000001", -- 1462 - 0x5b6  :    1 - 0x1
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- Sprite 0xb7
    "01011111", -- 1465 - 0x5b9  :   95 - 0x5f
    "01111111", -- 1466 - 0x5ba  :  127 - 0x7f
    "01111111", -- 1467 - 0x5bb  :  127 - 0x7f
    "00111111", -- 1468 - 0x5bc  :   63 - 0x3f
    "00111111", -- 1469 - 0x5bd  :   63 - 0x3f
    "00010100", -- 1470 - 0x5be  :   20 - 0x14
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0 -- Sprite 0xb8
    "11100000", -- 1473 - 0x5c1  :  224 - 0xe0
    "11110000", -- 1474 - 0x5c2  :  240 - 0xf0
    "00110000", -- 1475 - 0x5c3  :   48 - 0x30
    "00111000", -- 1476 - 0x5c4  :   56 - 0x38
    "00111100", -- 1477 - 0x5c5  :   60 - 0x3c
    "00111100", -- 1478 - 0x5c6  :   60 - 0x3c
    "11111100", -- 1479 - 0x5c7  :  252 - 0xfc
    "00000111", -- 1480 - 0x5c8  :    7 - 0x7 -- Sprite 0xb9
    "00001111", -- 1481 - 0x5c9  :   15 - 0xf
    "00011111", -- 1482 - 0x5ca  :   31 - 0x1f
    "00100010", -- 1483 - 0x5cb  :   34 - 0x22
    "00100000", -- 1484 - 0x5cc  :   32 - 0x20
    "00100101", -- 1485 - 0x5cd  :   37 - 0x25
    "00100101", -- 1486 - 0x5ce  :   37 - 0x25
    "00011111", -- 1487 - 0x5cf  :   31 - 0x1f
    "11111110", -- 1488 - 0x5d0  :  254 - 0xfe -- Sprite 0xba
    "11111110", -- 1489 - 0x5d1  :  254 - 0xfe
    "01111110", -- 1490 - 0x5d2  :  126 - 0x7e
    "00111010", -- 1491 - 0x5d3  :   58 - 0x3a
    "00000010", -- 1492 - 0x5d4  :    2 - 0x2
    "00000001", -- 1493 - 0x5d5  :    1 - 0x1
    "01000001", -- 1494 - 0x5d6  :   65 - 0x41
    "01000001", -- 1495 - 0x5d7  :   65 - 0x41
    "00011111", -- 1496 - 0x5d8  :   31 - 0x1f -- Sprite 0xbb
    "00111111", -- 1497 - 0x5d9  :   63 - 0x3f
    "01111110", -- 1498 - 0x5da  :  126 - 0x7e
    "01011100", -- 1499 - 0x5db  :   92 - 0x5c
    "01000000", -- 1500 - 0x5dc  :   64 - 0x40
    "10000000", -- 1501 - 0x5dd  :  128 - 0x80
    "10000010", -- 1502 - 0x5de  :  130 - 0x82
    "10000010", -- 1503 - 0x5df  :  130 - 0x82
    "10000010", -- 1504 - 0x5e0  :  130 - 0x82 -- Sprite 0xbc
    "10000000", -- 1505 - 0x5e1  :  128 - 0x80
    "10100000", -- 1506 - 0x5e2  :  160 - 0xa0
    "01000100", -- 1507 - 0x5e3  :   68 - 0x44
    "01000011", -- 1508 - 0x5e4  :   67 - 0x43
    "01000000", -- 1509 - 0x5e5  :   64 - 0x40
    "00100001", -- 1510 - 0x5e6  :   33 - 0x21
    "00011110", -- 1511 - 0x5e7  :   30 - 0x1e
    "00011100", -- 1512 - 0x5e8  :   28 - 0x1c -- Sprite 0xbd
    "00111111", -- 1513 - 0x5e9  :   63 - 0x3f
    "00111110", -- 1514 - 0x5ea  :   62 - 0x3e
    "00111100", -- 1515 - 0x5eb  :   60 - 0x3c
    "01000000", -- 1516 - 0x5ec  :   64 - 0x40
    "10000000", -- 1517 - 0x5ed  :  128 - 0x80
    "10000010", -- 1518 - 0x5ee  :  130 - 0x82
    "10000010", -- 1519 - 0x5ef  :  130 - 0x82
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "10000000", -- 1522 - 0x5f2  :  128 - 0x80
    "10000000", -- 1523 - 0x5f3  :  128 - 0x80
    "10010010", -- 1524 - 0x5f4  :  146 - 0x92
    "10011101", -- 1525 - 0x5f5  :  157 - 0x9d
    "11000111", -- 1526 - 0x5f6  :  199 - 0xc7
    "11101111", -- 1527 - 0x5f7  :  239 - 0xef
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00100011", -- 1529 - 0x5f9  :   35 - 0x23
    "00110011", -- 1530 - 0x5fa  :   51 - 0x33
    "00111111", -- 1531 - 0x5fb  :   63 - 0x3f
    "00111111", -- 1532 - 0x5fc  :   63 - 0x3f
    "01111111", -- 1533 - 0x5fd  :  127 - 0x7f
    "01111111", -- 1534 - 0x5fe  :  127 - 0x7f
    "01111111", -- 1535 - 0x5ff  :  127 - 0x7f
    "11111110", -- 1536 - 0x600  :  254 - 0xfe -- Sprite 0xc0
    "11111000", -- 1537 - 0x601  :  248 - 0xf8
    "10100000", -- 1538 - 0x602  :  160 - 0xa0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "10000000", -- 1542 - 0x606  :  128 - 0x80
    "10000000", -- 1543 - 0x607  :  128 - 0x80
    "01111110", -- 1544 - 0x608  :  126 - 0x7e -- Sprite 0xc1
    "01111111", -- 1545 - 0x609  :  127 - 0x7f
    "01111101", -- 1546 - 0x60a  :  125 - 0x7d
    "00111111", -- 1547 - 0x60b  :   63 - 0x3f
    "00011110", -- 1548 - 0x60c  :   30 - 0x1e
    "10001111", -- 1549 - 0x60d  :  143 - 0x8f
    "10001111", -- 1550 - 0x60e  :  143 - 0x8f
    "00011001", -- 1551 - 0x60f  :   25 - 0x19
    "11100000", -- 1552 - 0x610  :  224 - 0xe0 -- Sprite 0xc2
    "00001110", -- 1553 - 0x611  :   14 - 0xe
    "01110011", -- 1554 - 0x612  :  115 - 0x73
    "11110011", -- 1555 - 0x613  :  243 - 0xf3
    "11111001", -- 1556 - 0x614  :  249 - 0xf9
    "11111001", -- 1557 - 0x615  :  249 - 0xf9
    "11111000", -- 1558 - 0x616  :  248 - 0xf8
    "01110000", -- 1559 - 0x617  :  112 - 0x70
    "00001110", -- 1560 - 0x618  :   14 - 0xe -- Sprite 0xc3
    "01100110", -- 1561 - 0x619  :  102 - 0x66
    "11100010", -- 1562 - 0x61a  :  226 - 0xe2
    "11110110", -- 1563 - 0x61b  :  246 - 0xf6
    "11111111", -- 1564 - 0x61c  :  255 - 0xff
    "11111111", -- 1565 - 0x61d  :  255 - 0xff
    "00011111", -- 1566 - 0x61e  :   31 - 0x1f
    "10011000", -- 1567 - 0x61f  :  152 - 0x98
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000100", -- 1571 - 0x623  :    4 - 0x4
    "00001111", -- 1572 - 0x624  :   15 - 0xf
    "00001111", -- 1573 - 0x625  :   15 - 0xf
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000111", -- 1575 - 0x627  :    7 - 0x7
    "11110011", -- 1576 - 0x628  :  243 - 0xf3 -- Sprite 0xc5
    "11100111", -- 1577 - 0x629  :  231 - 0xe7
    "11101110", -- 1578 - 0x62a  :  238 - 0xee
    "11101100", -- 1579 - 0x62b  :  236 - 0xec
    "11001101", -- 1580 - 0x62c  :  205 - 0xcd
    "11001111", -- 1581 - 0x62d  :  207 - 0xcf
    "11001111", -- 1582 - 0x62e  :  207 - 0xcf
    "11011111", -- 1583 - 0x62f  :  223 - 0xdf
    "00100111", -- 1584 - 0x630  :   39 - 0x27 -- Sprite 0xc6
    "00111111", -- 1585 - 0x631  :   63 - 0x3f
    "00111111", -- 1586 - 0x632  :   63 - 0x3f
    "01111000", -- 1587 - 0x633  :  120 - 0x78
    "00111100", -- 1588 - 0x634  :   60 - 0x3c
    "00011111", -- 1589 - 0x635  :   31 - 0x1f
    "00011111", -- 1590 - 0x636  :   31 - 0x1f
    "01110011", -- 1591 - 0x637  :  115 - 0x73
    "10011111", -- 1592 - 0x638  :  159 - 0x9f -- Sprite 0xc7
    "00111110", -- 1593 - 0x639  :   62 - 0x3e
    "01111100", -- 1594 - 0x63a  :  124 - 0x7c
    "11111100", -- 1595 - 0x63b  :  252 - 0xfc
    "11111000", -- 1596 - 0x63c  :  248 - 0xf8
    "11111000", -- 1597 - 0x63d  :  248 - 0xf8
    "11000000", -- 1598 - 0x63e  :  192 - 0xc0
    "01000000", -- 1599 - 0x63f  :   64 - 0x40
    "01111111", -- 1600 - 0x640  :  127 - 0x7f -- Sprite 0xc8
    "01111110", -- 1601 - 0x641  :  126 - 0x7e
    "01111000", -- 1602 - 0x642  :  120 - 0x78
    "00000001", -- 1603 - 0x643  :    1 - 0x1
    "00000111", -- 1604 - 0x644  :    7 - 0x7
    "00011111", -- 1605 - 0x645  :   31 - 0x1f
    "00111100", -- 1606 - 0x646  :   60 - 0x3c
    "01111100", -- 1607 - 0x647  :  124 - 0x7c
    "11111100", -- 1608 - 0x648  :  252 - 0xfc -- Sprite 0xc9
    "11111000", -- 1609 - 0x649  :  248 - 0xf8
    "10100000", -- 1610 - 0x64a  :  160 - 0xa0
    "11111110", -- 1611 - 0x64b  :  254 - 0xfe
    "11111100", -- 1612 - 0x64c  :  252 - 0xfc
    "11110000", -- 1613 - 0x64d  :  240 - 0xf0
    "10000000", -- 1614 - 0x64e  :  128 - 0x80
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "01111110", -- 1616 - 0x650  :  126 - 0x7e -- Sprite 0xca
    "01111111", -- 1617 - 0x651  :  127 - 0x7f
    "01111111", -- 1618 - 0x652  :  127 - 0x7f
    "00111111", -- 1619 - 0x653  :   63 - 0x3f
    "00011111", -- 1620 - 0x654  :   31 - 0x1f
    "10001111", -- 1621 - 0x655  :  143 - 0x8f
    "10001111", -- 1622 - 0x656  :  143 - 0x8f
    "00011000", -- 1623 - 0x657  :   24 - 0x18
    "10011111", -- 1624 - 0x658  :  159 - 0x9f -- Sprite 0xcb
    "00111110", -- 1625 - 0x659  :   62 - 0x3e
    "01111100", -- 1626 - 0x65a  :  124 - 0x7c
    "11111000", -- 1627 - 0x65b  :  248 - 0xf8
    "11111000", -- 1628 - 0x65c  :  248 - 0xf8
    "00111100", -- 1629 - 0x65d  :   60 - 0x3c
    "00011000", -- 1630 - 0x65e  :   24 - 0x18
    "11111000", -- 1631 - 0x65f  :  248 - 0xf8
    "01111111", -- 1632 - 0x660  :  127 - 0x7f -- Sprite 0xcc
    "01111111", -- 1633 - 0x661  :  127 - 0x7f
    "01111000", -- 1634 - 0x662  :  120 - 0x78
    "00000001", -- 1635 - 0x663  :    1 - 0x1
    "00000111", -- 1636 - 0x664  :    7 - 0x7
    "00010011", -- 1637 - 0x665  :   19 - 0x13
    "11110001", -- 1638 - 0x666  :  241 - 0xf1
    "00000011", -- 1639 - 0x667  :    3 - 0x3
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00011100", -- 1642 - 0x66a  :   28 - 0x1c
    "00011101", -- 1643 - 0x66b  :   29 - 0x1d
    "00011011", -- 1644 - 0x66c  :   27 - 0x1b
    "11000011", -- 1645 - 0x66d  :  195 - 0xc3
    "11100011", -- 1646 - 0x66e  :  227 - 0xe3
    "11100001", -- 1647 - 0x66f  :  225 - 0xe1
    "11100000", -- 1648 - 0x670  :  224 - 0xe0 -- Sprite 0xce
    "11001101", -- 1649 - 0x671  :  205 - 0xcd
    "00011101", -- 1650 - 0x672  :   29 - 0x1d
    "01001111", -- 1651 - 0x673  :   79 - 0x4f
    "11101110", -- 1652 - 0x674  :  238 - 0xee
    "11111111", -- 1653 - 0x675  :  255 - 0xff
    "00111111", -- 1654 - 0x676  :   63 - 0x3f
    "00111111", -- 1655 - 0x677  :   63 - 0x3f
    "00111111", -- 1656 - 0x678  :   63 - 0x3f -- Sprite 0xcf
    "00111111", -- 1657 - 0x679  :   63 - 0x3f
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "01110000", -- 1660 - 0x67c  :  112 - 0x70
    "10111000", -- 1661 - 0x67d  :  184 - 0xb8
    "11111100", -- 1662 - 0x67e  :  252 - 0xfc
    "11111100", -- 1663 - 0x67f  :  252 - 0xfc
    "00000111", -- 1664 - 0x680  :    7 - 0x7 -- Sprite 0xd0
    "00001111", -- 1665 - 0x681  :   15 - 0xf
    "00011111", -- 1666 - 0x682  :   31 - 0x1f
    "00111111", -- 1667 - 0x683  :   63 - 0x3f
    "00111110", -- 1668 - 0x684  :   62 - 0x3e
    "01111100", -- 1669 - 0x685  :  124 - 0x7c
    "01111000", -- 1670 - 0x686  :  120 - 0x78
    "01111000", -- 1671 - 0x687  :  120 - 0x78
    "00111111", -- 1672 - 0x688  :   63 - 0x3f -- Sprite 0xd1
    "01011100", -- 1673 - 0x689  :   92 - 0x5c
    "00111001", -- 1674 - 0x68a  :   57 - 0x39
    "00111011", -- 1675 - 0x68b  :   59 - 0x3b
    "10111111", -- 1676 - 0x68c  :  191 - 0xbf
    "11111111", -- 1677 - 0x68d  :  255 - 0xff
    "11111110", -- 1678 - 0x68e  :  254 - 0xfe
    "11111110", -- 1679 - 0x68f  :  254 - 0xfe
    "11000000", -- 1680 - 0x690  :  192 - 0xc0 -- Sprite 0xd2
    "11000000", -- 1681 - 0x691  :  192 - 0xc0
    "10000000", -- 1682 - 0x692  :  128 - 0x80
    "10000000", -- 1683 - 0x693  :  128 - 0x80
    "10000000", -- 1684 - 0x694  :  128 - 0x80
    "10000000", -- 1685 - 0x695  :  128 - 0x80
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "11111110", -- 1688 - 0x698  :  254 - 0xfe -- Sprite 0xd3
    "11111100", -- 1689 - 0x699  :  252 - 0xfc
    "01100001", -- 1690 - 0x69a  :   97 - 0x61
    "00001111", -- 1691 - 0x69b  :   15 - 0xf
    "01111111", -- 1692 - 0x69c  :  127 - 0x7f
    "00111111", -- 1693 - 0x69d  :   63 - 0x3f
    "00011111", -- 1694 - 0x69e  :   31 - 0x1f
    "00011110", -- 1695 - 0x69f  :   30 - 0x1e
    "11110000", -- 1696 - 0x6a0  :  240 - 0xf0 -- Sprite 0xd4
    "01111000", -- 1697 - 0x6a1  :  120 - 0x78
    "11100100", -- 1698 - 0x6a2  :  228 - 0xe4
    "11001000", -- 1699 - 0x6a3  :  200 - 0xc8
    "11001100", -- 1700 - 0x6a4  :  204 - 0xcc
    "10111110", -- 1701 - 0x6a5  :  190 - 0xbe
    "10111110", -- 1702 - 0x6a6  :  190 - 0xbe
    "00111110", -- 1703 - 0x6a7  :   62 - 0x3e
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "00000001", -- 1705 - 0x6a9  :    1 - 0x1
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000111", -- 1707 - 0x6ab  :    7 - 0x7
    "00000111", -- 1708 - 0x6ac  :    7 - 0x7
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000111", -- 1710 - 0x6ae  :    7 - 0x7
    "00011111", -- 1711 - 0x6af  :   31 - 0x1f
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00001111", -- 1714 - 0x6b2  :   15 - 0xf
    "00111111", -- 1715 - 0x6b3  :   63 - 0x3f
    "00111111", -- 1716 - 0x6b4  :   63 - 0x3f
    "00001111", -- 1717 - 0x6b5  :   15 - 0xf
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "01111000", -- 1720 - 0x6b8  :  120 - 0x78 -- Sprite 0xd7
    "01111100", -- 1721 - 0x6b9  :  124 - 0x7c
    "01111110", -- 1722 - 0x6ba  :  126 - 0x7e
    "01111111", -- 1723 - 0x6bb  :  127 - 0x7f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00111111", -- 1725 - 0x6bd  :   63 - 0x3f
    "00011011", -- 1726 - 0x6be  :   27 - 0x1b
    "00001001", -- 1727 - 0x6bf  :    9 - 0x9
    "00001100", -- 1728 - 0x6c0  :   12 - 0xc -- Sprite 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000111", -- 1732 - 0x6c4  :    7 - 0x7
    "01111111", -- 1733 - 0x6c5  :  127 - 0x7f
    "01111100", -- 1734 - 0x6c6  :  124 - 0x7c
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000001", -- 1736 - 0x6c8  :    1 - 0x1 -- Sprite 0xd9
    "11100001", -- 1737 - 0x6c9  :  225 - 0xe1
    "01110001", -- 1738 - 0x6ca  :  113 - 0x71
    "01111001", -- 1739 - 0x6cb  :  121 - 0x79
    "00111101", -- 1740 - 0x6cc  :   61 - 0x3d
    "00111101", -- 1741 - 0x6cd  :   61 - 0x3d
    "00011111", -- 1742 - 0x6ce  :   31 - 0x1f
    "00000011", -- 1743 - 0x6cf  :    3 - 0x3
    "00111111", -- 1744 - 0x6d0  :   63 - 0x3f -- Sprite 0xda
    "00111111", -- 1745 - 0x6d1  :   63 - 0x3f
    "00011111", -- 1746 - 0x6d2  :   31 - 0x1f
    "00011011", -- 1747 - 0x6d3  :   27 - 0x1b
    "00110110", -- 1748 - 0x6d4  :   54 - 0x36
    "00110000", -- 1749 - 0x6d5  :   48 - 0x30
    "01111111", -- 1750 - 0x6d6  :  127 - 0x7f
    "00111111", -- 1751 - 0x6d7  :   63 - 0x3f
    "11111000", -- 1752 - 0x6d8  :  248 - 0xf8 -- Sprite 0xdb
    "11111000", -- 1753 - 0x6d9  :  248 - 0xf8
    "11111000", -- 1754 - 0x6da  :  248 - 0xf8
    "10111000", -- 1755 - 0x6db  :  184 - 0xb8
    "00011000", -- 1756 - 0x6dc  :   24 - 0x18
    "11011000", -- 1757 - 0x6dd  :  216 - 0xd8
    "11011000", -- 1758 - 0x6de  :  216 - 0xd8
    "10111000", -- 1759 - 0x6df  :  184 - 0xb8
    "00000001", -- 1760 - 0x6e0  :    1 - 0x1 -- Sprite 0xdc
    "00000010", -- 1761 - 0x6e1  :    2 - 0x2
    "00000100", -- 1762 - 0x6e2  :    4 - 0x4
    "00000100", -- 1763 - 0x6e3  :    4 - 0x4
    "00001000", -- 1764 - 0x6e4  :    8 - 0x8
    "00001000", -- 1765 - 0x6e5  :    8 - 0x8
    "00010000", -- 1766 - 0x6e6  :   16 - 0x10
    "00010000", -- 1767 - 0x6e7  :   16 - 0x10
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00001111", -- 1769 - 0x6e9  :   15 - 0xf
    "00010011", -- 1770 - 0x6ea  :   19 - 0x13
    "00001101", -- 1771 - 0x6eb  :   13 - 0xd
    "00001101", -- 1772 - 0x6ec  :   13 - 0xd
    "00010011", -- 1773 - 0x6ed  :   19 - 0x13
    "00001100", -- 1774 - 0x6ee  :   12 - 0xc
    "00100000", -- 1775 - 0x6ef  :   32 - 0x20
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0 -- Sprite 0xde
    "00100100", -- 1777 - 0x6f1  :   36 - 0x24
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00100100", -- 1779 - 0x6f3  :   36 - 0x24
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000100", -- 1781 - 0x6f5  :    4 - 0x4
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00001111", -- 1784 - 0x6f8  :   15 - 0xf -- Sprite 0xdf
    "01000001", -- 1785 - 0x6f9  :   65 - 0x41
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "10001000", -- 1787 - 0x6fb  :  136 - 0x88
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "01000100", -- 1789 - 0x6fd  :   68 - 0x44
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00111000", -- 1792 - 0x700  :   56 - 0x38 -- Sprite 0xe0
    "01111100", -- 1793 - 0x701  :  124 - 0x7c
    "11111110", -- 1794 - 0x702  :  254 - 0xfe
    "11111110", -- 1795 - 0x703  :  254 - 0xfe
    "00111011", -- 1796 - 0x704  :   59 - 0x3b
    "00000011", -- 1797 - 0x705  :    3 - 0x3
    "00000011", -- 1798 - 0x706  :    3 - 0x3
    "00000011", -- 1799 - 0x707  :    3 - 0x3
    "00000011", -- 1800 - 0x708  :    3 - 0x3 -- Sprite 0xe1
    "00110011", -- 1801 - 0x709  :   51 - 0x33
    "01111011", -- 1802 - 0x70a  :  123 - 0x7b
    "01111111", -- 1803 - 0x70b  :  127 - 0x7f
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111011", -- 1805 - 0x70d  :  251 - 0xfb
    "00000011", -- 1806 - 0x70e  :    3 - 0x3
    "00000011", -- 1807 - 0x70f  :    3 - 0x3
    "11011100", -- 1808 - 0x710  :  220 - 0xdc -- Sprite 0xe2
    "11000000", -- 1809 - 0x711  :  192 - 0xc0
    "11100000", -- 1810 - 0x712  :  224 - 0xe0
    "11100000", -- 1811 - 0x713  :  224 - 0xe0
    "11100000", -- 1812 - 0x714  :  224 - 0xe0
    "11100000", -- 1813 - 0x715  :  224 - 0xe0
    "11100000", -- 1814 - 0x716  :  224 - 0xe0
    "11000000", -- 1815 - 0x717  :  192 - 0xc0
    "00111111", -- 1816 - 0x718  :   63 - 0x3f -- Sprite 0xe3
    "01011111", -- 1817 - 0x719  :   95 - 0x5f
    "00111111", -- 1818 - 0x71a  :   63 - 0x3f
    "00111111", -- 1819 - 0x71b  :   63 - 0x3f
    "10111011", -- 1820 - 0x71c  :  187 - 0xbb
    "11111000", -- 1821 - 0x71d  :  248 - 0xf8
    "11111110", -- 1822 - 0x71e  :  254 - 0xfe
    "11111110", -- 1823 - 0x71f  :  254 - 0xfe
    "00011111", -- 1824 - 0x720  :   31 - 0x1f -- Sprite 0xe4
    "00001111", -- 1825 - 0x721  :   15 - 0xf
    "00001111", -- 1826 - 0x722  :   15 - 0xf
    "00011111", -- 1827 - 0x723  :   31 - 0x1f
    "00011111", -- 1828 - 0x724  :   31 - 0x1f
    "00011110", -- 1829 - 0x725  :   30 - 0x1e
    "00111000", -- 1830 - 0x726  :   56 - 0x38
    "00110000", -- 1831 - 0x727  :   48 - 0x30
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00100000", -- 1833 - 0x729  :   32 - 0x20
    "01100000", -- 1834 - 0x72a  :   96 - 0x60
    "01100000", -- 1835 - 0x72b  :   96 - 0x60
    "01110000", -- 1836 - 0x72c  :  112 - 0x70
    "11110000", -- 1837 - 0x72d  :  240 - 0xf0
    "11111000", -- 1838 - 0x72e  :  248 - 0xf8
    "11111000", -- 1839 - 0x72f  :  248 - 0xf8
    "11111000", -- 1840 - 0x730  :  248 - 0xf8 -- Sprite 0xe6
    "11111100", -- 1841 - 0x731  :  252 - 0xfc
    "11111100", -- 1842 - 0x732  :  252 - 0xfc
    "01111110", -- 1843 - 0x733  :  126 - 0x7e
    "01111110", -- 1844 - 0x734  :  126 - 0x7e
    "00111110", -- 1845 - 0x735  :   62 - 0x3e
    "00011111", -- 1846 - 0x736  :   31 - 0x1f
    "00000111", -- 1847 - 0x737  :    7 - 0x7
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "11000000", -- 1849 - 0x739  :  192 - 0xc0
    "01110000", -- 1850 - 0x73a  :  112 - 0x70
    "10111000", -- 1851 - 0x73b  :  184 - 0xb8
    "11110100", -- 1852 - 0x73c  :  244 - 0xf4
    "11110010", -- 1853 - 0x73d  :  242 - 0xf2
    "11110101", -- 1854 - 0x73e  :  245 - 0xf5
    "01111011", -- 1855 - 0x73f  :  123 - 0x7b
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "11011111", -- 1857 - 0x741  :  223 - 0xdf
    "00010000", -- 1858 - 0x742  :   16 - 0x10
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11011111", -- 1860 - 0x744  :  223 - 0xdf
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111001", -- 1863 - 0x747  :  249 - 0xf9
    "00011111", -- 1864 - 0x748  :   31 - 0x1f -- Sprite 0xe9
    "00011111", -- 1865 - 0x749  :   31 - 0x1f
    "00111110", -- 1866 - 0x74a  :   62 - 0x3e
    "11111100", -- 1867 - 0x74b  :  252 - 0xfc
    "11111000", -- 1868 - 0x74c  :  248 - 0xf8
    "11110000", -- 1869 - 0x74d  :  240 - 0xf0
    "11000000", -- 1870 - 0x74e  :  192 - 0xc0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "11111000", -- 1872 - 0x750  :  248 - 0xf8 -- Sprite 0xea
    "11111100", -- 1873 - 0x751  :  252 - 0xfc
    "11111110", -- 1874 - 0x752  :  254 - 0xfe
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11011111", -- 1877 - 0x755  :  223 - 0xdf
    "11011111", -- 1878 - 0x756  :  223 - 0xdf
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "11000001", -- 1880 - 0x758  :  193 - 0xc1 -- Sprite 0xeb
    "11110001", -- 1881 - 0x759  :  241 - 0xf1
    "01111001", -- 1882 - 0x75a  :  121 - 0x79
    "01111101", -- 1883 - 0x75b  :  125 - 0x7d
    "00111101", -- 1884 - 0x75c  :   61 - 0x3d
    "00111111", -- 1885 - 0x75d  :   63 - 0x3f
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000011", -- 1887 - 0x75f  :    3 - 0x3
    "00000010", -- 1888 - 0x760  :    2 - 0x2 -- Sprite 0xec
    "00000110", -- 1889 - 0x761  :    6 - 0x6
    "00001110", -- 1890 - 0x762  :   14 - 0xe
    "00001110", -- 1891 - 0x763  :   14 - 0xe
    "00011110", -- 1892 - 0x764  :   30 - 0x1e
    "00011110", -- 1893 - 0x765  :   30 - 0x1e
    "00111110", -- 1894 - 0x766  :   62 - 0x3e
    "00111110", -- 1895 - 0x767  :   62 - 0x3e
    "00111110", -- 1896 - 0x768  :   62 - 0x3e -- Sprite 0xed
    "00111110", -- 1897 - 0x769  :   62 - 0x3e
    "00111110", -- 1898 - 0x76a  :   62 - 0x3e
    "00111110", -- 1899 - 0x76b  :   62 - 0x3e
    "00011110", -- 1900 - 0x76c  :   30 - 0x1e
    "00011110", -- 1901 - 0x76d  :   30 - 0x1e
    "00001110", -- 1902 - 0x76e  :   14 - 0xe
    "00000010", -- 1903 - 0x76f  :    2 - 0x2
    "11000001", -- 1904 - 0x770  :  193 - 0xc1 -- Sprite 0xee
    "11110001", -- 1905 - 0x771  :  241 - 0xf1
    "01111001", -- 1906 - 0x772  :  121 - 0x79
    "01111101", -- 1907 - 0x773  :  125 - 0x7d
    "00111101", -- 1908 - 0x774  :   61 - 0x3d
    "00111111", -- 1909 - 0x775  :   63 - 0x3f
    "00011111", -- 1910 - 0x776  :   31 - 0x1f
    "00000011", -- 1911 - 0x777  :    3 - 0x3
    "01111100", -- 1912 - 0x778  :  124 - 0x7c -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11000011", -- 1916 - 0x77c  :  195 - 0xc3
    "01111111", -- 1917 - 0x77d  :  127 - 0x7f
    "00011111", -- 1918 - 0x77e  :   31 - 0x1f
    "00000011", -- 1919 - 0x77f  :    3 - 0x3
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "01111100", -- 1922 - 0x782  :  124 - 0x7c
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "01111100", -- 1925 - 0x785  :  124 - 0x7c
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000100", -- 1931 - 0x78b  :    4 - 0x4
    "00001100", -- 1932 - 0x78c  :   12 - 0xc
    "00011000", -- 1933 - 0x78d  :   24 - 0x18
    "00110000", -- 1934 - 0x78e  :   48 - 0x30
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000100", -- 1939 - 0x793  :    4 - 0x4
    "00000100", -- 1940 - 0x794  :    4 - 0x4
    "00000100", -- 1941 - 0x795  :    4 - 0x4
    "00001000", -- 1942 - 0x796  :    8 - 0x8
    "00001000", -- 1943 - 0x797  :    8 - 0x8
    "00001000", -- 1944 - 0x798  :    8 - 0x8 -- Sprite 0xf3
    "00010000", -- 1945 - 0x799  :   16 - 0x10
    "00010000", -- 1946 - 0x79a  :   16 - 0x10
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00010000", -- 1949 - 0x79d  :   16 - 0x10
    "00010000", -- 1950 - 0x79e  :   16 - 0x10
    "00001000", -- 1951 - 0x79f  :    8 - 0x8
    "01111111", -- 1952 - 0x7a0  :  127 - 0x7f -- Sprite 0xf4
    "00111111", -- 1953 - 0x7a1  :   63 - 0x3f
    "00111111", -- 1954 - 0x7a2  :   63 - 0x3f
    "00111110", -- 1955 - 0x7a3  :   62 - 0x3e
    "00011111", -- 1956 - 0x7a4  :   31 - 0x1f
    "00001111", -- 1957 - 0x7a5  :   15 - 0xf
    "00000011", -- 1958 - 0x7a6  :    3 - 0x3
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000011", -- 1960 - 0x7a8  :    3 - 0x3 -- Sprite 0xf5
    "00001111", -- 1961 - 0x7a9  :   15 - 0xf
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "01111111", -- 1963 - 0x7ab  :  127 - 0x7f
    "01111111", -- 1964 - 0x7ac  :  127 - 0x7f
    "01111111", -- 1965 - 0x7ad  :  127 - 0x7f
    "01111111", -- 1966 - 0x7ae  :  127 - 0x7f
    "01111111", -- 1967 - 0x7af  :  127 - 0x7f
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "01111100", -- 2045 - 0x7fd  :  124 - 0x7c
    "00111000", -- 2046 - 0x7fe  :   56 - 0x38
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
          -- Background pattern Table
    "00111000", -- 2048 - 0x800  :   56 - 0x38 -- Background 0x0
    "01001100", -- 2049 - 0x801  :   76 - 0x4c
    "11000110", -- 2050 - 0x802  :  198 - 0xc6
    "11000110", -- 2051 - 0x803  :  198 - 0xc6
    "11000110", -- 2052 - 0x804  :  198 - 0xc6
    "01100100", -- 2053 - 0x805  :  100 - 0x64
    "00111000", -- 2054 - 0x806  :   56 - 0x38
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00011000", -- 2056 - 0x808  :   24 - 0x18 -- Background 0x1
    "00111000", -- 2057 - 0x809  :   56 - 0x38
    "00011000", -- 2058 - 0x80a  :   24 - 0x18
    "00011000", -- 2059 - 0x80b  :   24 - 0x18
    "00011000", -- 2060 - 0x80c  :   24 - 0x18
    "00011000", -- 2061 - 0x80d  :   24 - 0x18
    "01111110", -- 2062 - 0x80e  :  126 - 0x7e
    "00000000", -- 2063 - 0x80f  :    0 - 0x0
    "01111100", -- 2064 - 0x810  :  124 - 0x7c -- Background 0x2
    "11000110", -- 2065 - 0x811  :  198 - 0xc6
    "00001110", -- 2066 - 0x812  :   14 - 0xe
    "00111100", -- 2067 - 0x813  :   60 - 0x3c
    "01111000", -- 2068 - 0x814  :  120 - 0x78
    "11100000", -- 2069 - 0x815  :  224 - 0xe0
    "11111110", -- 2070 - 0x816  :  254 - 0xfe
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "01111110", -- 2072 - 0x818  :  126 - 0x7e -- Background 0x3
    "00001100", -- 2073 - 0x819  :   12 - 0xc
    "00011000", -- 2074 - 0x81a  :   24 - 0x18
    "00111100", -- 2075 - 0x81b  :   60 - 0x3c
    "00000110", -- 2076 - 0x81c  :    6 - 0x6
    "11000110", -- 2077 - 0x81d  :  198 - 0xc6
    "01111100", -- 2078 - 0x81e  :  124 - 0x7c
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00011100", -- 2080 - 0x820  :   28 - 0x1c -- Background 0x4
    "00111100", -- 2081 - 0x821  :   60 - 0x3c
    "01101100", -- 2082 - 0x822  :  108 - 0x6c
    "11001100", -- 2083 - 0x823  :  204 - 0xcc
    "11111110", -- 2084 - 0x824  :  254 - 0xfe
    "00001100", -- 2085 - 0x825  :   12 - 0xc
    "00001100", -- 2086 - 0x826  :   12 - 0xc
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "11111100", -- 2088 - 0x828  :  252 - 0xfc -- Background 0x5
    "11000000", -- 2089 - 0x829  :  192 - 0xc0
    "11111100", -- 2090 - 0x82a  :  252 - 0xfc
    "00000110", -- 2091 - 0x82b  :    6 - 0x6
    "00000110", -- 2092 - 0x82c  :    6 - 0x6
    "11000110", -- 2093 - 0x82d  :  198 - 0xc6
    "01111100", -- 2094 - 0x82e  :  124 - 0x7c
    "00000000", -- 2095 - 0x82f  :    0 - 0x0
    "00111100", -- 2096 - 0x830  :   60 - 0x3c -- Background 0x6
    "01100000", -- 2097 - 0x831  :   96 - 0x60
    "11000000", -- 2098 - 0x832  :  192 - 0xc0
    "11111100", -- 2099 - 0x833  :  252 - 0xfc
    "11000110", -- 2100 - 0x834  :  198 - 0xc6
    "11000110", -- 2101 - 0x835  :  198 - 0xc6
    "01111100", -- 2102 - 0x836  :  124 - 0x7c
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "11111110", -- 2104 - 0x838  :  254 - 0xfe -- Background 0x7
    "11000110", -- 2105 - 0x839  :  198 - 0xc6
    "00001100", -- 2106 - 0x83a  :   12 - 0xc
    "00011000", -- 2107 - 0x83b  :   24 - 0x18
    "00110000", -- 2108 - 0x83c  :   48 - 0x30
    "00110000", -- 2109 - 0x83d  :   48 - 0x30
    "00110000", -- 2110 - 0x83e  :   48 - 0x30
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "01111100", -- 2112 - 0x840  :  124 - 0x7c -- Background 0x8
    "11000110", -- 2113 - 0x841  :  198 - 0xc6
    "11000110", -- 2114 - 0x842  :  198 - 0xc6
    "01111100", -- 2115 - 0x843  :  124 - 0x7c
    "11000110", -- 2116 - 0x844  :  198 - 0xc6
    "11000110", -- 2117 - 0x845  :  198 - 0xc6
    "01111100", -- 2118 - 0x846  :  124 - 0x7c
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "01111100", -- 2120 - 0x848  :  124 - 0x7c -- Background 0x9
    "11000110", -- 2121 - 0x849  :  198 - 0xc6
    "11000110", -- 2122 - 0x84a  :  198 - 0xc6
    "01111110", -- 2123 - 0x84b  :  126 - 0x7e
    "00000110", -- 2124 - 0x84c  :    6 - 0x6
    "00001100", -- 2125 - 0x84d  :   12 - 0xc
    "01111000", -- 2126 - 0x84e  :  120 - 0x78
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00111000", -- 2128 - 0x850  :   56 - 0x38 -- Background 0xa
    "01101100", -- 2129 - 0x851  :  108 - 0x6c
    "11000110", -- 2130 - 0x852  :  198 - 0xc6
    "11000110", -- 2131 - 0x853  :  198 - 0xc6
    "11111110", -- 2132 - 0x854  :  254 - 0xfe
    "11000110", -- 2133 - 0x855  :  198 - 0xc6
    "11000110", -- 2134 - 0x856  :  198 - 0xc6
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "11111100", -- 2136 - 0x858  :  252 - 0xfc -- Background 0xb
    "11000110", -- 2137 - 0x859  :  198 - 0xc6
    "11000110", -- 2138 - 0x85a  :  198 - 0xc6
    "11111100", -- 2139 - 0x85b  :  252 - 0xfc
    "11000110", -- 2140 - 0x85c  :  198 - 0xc6
    "11000110", -- 2141 - 0x85d  :  198 - 0xc6
    "11111100", -- 2142 - 0x85e  :  252 - 0xfc
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00111100", -- 2144 - 0x860  :   60 - 0x3c -- Background 0xc
    "01100110", -- 2145 - 0x861  :  102 - 0x66
    "11000000", -- 2146 - 0x862  :  192 - 0xc0
    "11000000", -- 2147 - 0x863  :  192 - 0xc0
    "11000000", -- 2148 - 0x864  :  192 - 0xc0
    "01100110", -- 2149 - 0x865  :  102 - 0x66
    "00111100", -- 2150 - 0x866  :   60 - 0x3c
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "11111000", -- 2152 - 0x868  :  248 - 0xf8 -- Background 0xd
    "11001100", -- 2153 - 0x869  :  204 - 0xcc
    "11000110", -- 2154 - 0x86a  :  198 - 0xc6
    "11000110", -- 2155 - 0x86b  :  198 - 0xc6
    "11000110", -- 2156 - 0x86c  :  198 - 0xc6
    "11001100", -- 2157 - 0x86d  :  204 - 0xcc
    "11111000", -- 2158 - 0x86e  :  248 - 0xf8
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "11111110", -- 2160 - 0x870  :  254 - 0xfe -- Background 0xe
    "11000000", -- 2161 - 0x871  :  192 - 0xc0
    "11000000", -- 2162 - 0x872  :  192 - 0xc0
    "11111100", -- 2163 - 0x873  :  252 - 0xfc
    "11000000", -- 2164 - 0x874  :  192 - 0xc0
    "11000000", -- 2165 - 0x875  :  192 - 0xc0
    "11111110", -- 2166 - 0x876  :  254 - 0xfe
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "11111110", -- 2168 - 0x878  :  254 - 0xfe -- Background 0xf
    "11000000", -- 2169 - 0x879  :  192 - 0xc0
    "11000000", -- 2170 - 0x87a  :  192 - 0xc0
    "11111100", -- 2171 - 0x87b  :  252 - 0xfc
    "11000000", -- 2172 - 0x87c  :  192 - 0xc0
    "11000000", -- 2173 - 0x87d  :  192 - 0xc0
    "11000000", -- 2174 - 0x87e  :  192 - 0xc0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00111110", -- 2176 - 0x880  :   62 - 0x3e -- Background 0x10
    "01100000", -- 2177 - 0x881  :   96 - 0x60
    "11000000", -- 2178 - 0x882  :  192 - 0xc0
    "11001110", -- 2179 - 0x883  :  206 - 0xce
    "11000110", -- 2180 - 0x884  :  198 - 0xc6
    "01100110", -- 2181 - 0x885  :  102 - 0x66
    "00111110", -- 2182 - 0x886  :   62 - 0x3e
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "11000110", -- 2184 - 0x888  :  198 - 0xc6 -- Background 0x11
    "11000110", -- 2185 - 0x889  :  198 - 0xc6
    "11000110", -- 2186 - 0x88a  :  198 - 0xc6
    "11111110", -- 2187 - 0x88b  :  254 - 0xfe
    "11000110", -- 2188 - 0x88c  :  198 - 0xc6
    "11000110", -- 2189 - 0x88d  :  198 - 0xc6
    "11000110", -- 2190 - 0x88e  :  198 - 0xc6
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "01111110", -- 2192 - 0x890  :  126 - 0x7e -- Background 0x12
    "00011000", -- 2193 - 0x891  :   24 - 0x18
    "00011000", -- 2194 - 0x892  :   24 - 0x18
    "00011000", -- 2195 - 0x893  :   24 - 0x18
    "00011000", -- 2196 - 0x894  :   24 - 0x18
    "00011000", -- 2197 - 0x895  :   24 - 0x18
    "01111110", -- 2198 - 0x896  :  126 - 0x7e
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00011110", -- 2200 - 0x898  :   30 - 0x1e -- Background 0x13
    "00000110", -- 2201 - 0x899  :    6 - 0x6
    "00000110", -- 2202 - 0x89a  :    6 - 0x6
    "00000110", -- 2203 - 0x89b  :    6 - 0x6
    "11000110", -- 2204 - 0x89c  :  198 - 0xc6
    "11000110", -- 2205 - 0x89d  :  198 - 0xc6
    "01111100", -- 2206 - 0x89e  :  124 - 0x7c
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "11000110", -- 2208 - 0x8a0  :  198 - 0xc6 -- Background 0x14
    "11001100", -- 2209 - 0x8a1  :  204 - 0xcc
    "11011000", -- 2210 - 0x8a2  :  216 - 0xd8
    "11110000", -- 2211 - 0x8a3  :  240 - 0xf0
    "11111000", -- 2212 - 0x8a4  :  248 - 0xf8
    "11011100", -- 2213 - 0x8a5  :  220 - 0xdc
    "11001110", -- 2214 - 0x8a6  :  206 - 0xce
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "01100000", -- 2216 - 0x8a8  :   96 - 0x60 -- Background 0x15
    "01100000", -- 2217 - 0x8a9  :   96 - 0x60
    "01100000", -- 2218 - 0x8aa  :   96 - 0x60
    "01100000", -- 2219 - 0x8ab  :   96 - 0x60
    "01100000", -- 2220 - 0x8ac  :   96 - 0x60
    "01100000", -- 2221 - 0x8ad  :   96 - 0x60
    "01111110", -- 2222 - 0x8ae  :  126 - 0x7e
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "11000110", -- 2224 - 0x8b0  :  198 - 0xc6 -- Background 0x16
    "11101110", -- 2225 - 0x8b1  :  238 - 0xee
    "11111110", -- 2226 - 0x8b2  :  254 - 0xfe
    "11111110", -- 2227 - 0x8b3  :  254 - 0xfe
    "11010110", -- 2228 - 0x8b4  :  214 - 0xd6
    "11000110", -- 2229 - 0x8b5  :  198 - 0xc6
    "11000110", -- 2230 - 0x8b6  :  198 - 0xc6
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "11000110", -- 2232 - 0x8b8  :  198 - 0xc6 -- Background 0x17
    "11100110", -- 2233 - 0x8b9  :  230 - 0xe6
    "11110110", -- 2234 - 0x8ba  :  246 - 0xf6
    "11111110", -- 2235 - 0x8bb  :  254 - 0xfe
    "11011110", -- 2236 - 0x8bc  :  222 - 0xde
    "11001110", -- 2237 - 0x8bd  :  206 - 0xce
    "11000110", -- 2238 - 0x8be  :  198 - 0xc6
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "01111100", -- 2240 - 0x8c0  :  124 - 0x7c -- Background 0x18
    "11000110", -- 2241 - 0x8c1  :  198 - 0xc6
    "11000110", -- 2242 - 0x8c2  :  198 - 0xc6
    "11000110", -- 2243 - 0x8c3  :  198 - 0xc6
    "11000110", -- 2244 - 0x8c4  :  198 - 0xc6
    "11000110", -- 2245 - 0x8c5  :  198 - 0xc6
    "01111100", -- 2246 - 0x8c6  :  124 - 0x7c
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "11111100", -- 2248 - 0x8c8  :  252 - 0xfc -- Background 0x19
    "11000110", -- 2249 - 0x8c9  :  198 - 0xc6
    "11000110", -- 2250 - 0x8ca  :  198 - 0xc6
    "11000110", -- 2251 - 0x8cb  :  198 - 0xc6
    "11111100", -- 2252 - 0x8cc  :  252 - 0xfc
    "11000000", -- 2253 - 0x8cd  :  192 - 0xc0
    "11000000", -- 2254 - 0x8ce  :  192 - 0xc0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "01111100", -- 2256 - 0x8d0  :  124 - 0x7c -- Background 0x1a
    "11000110", -- 2257 - 0x8d1  :  198 - 0xc6
    "11000110", -- 2258 - 0x8d2  :  198 - 0xc6
    "11000110", -- 2259 - 0x8d3  :  198 - 0xc6
    "11011110", -- 2260 - 0x8d4  :  222 - 0xde
    "11001100", -- 2261 - 0x8d5  :  204 - 0xcc
    "01111010", -- 2262 - 0x8d6  :  122 - 0x7a
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "11111100", -- 2264 - 0x8d8  :  252 - 0xfc -- Background 0x1b
    "11000110", -- 2265 - 0x8d9  :  198 - 0xc6
    "11000110", -- 2266 - 0x8da  :  198 - 0xc6
    "11001110", -- 2267 - 0x8db  :  206 - 0xce
    "11111000", -- 2268 - 0x8dc  :  248 - 0xf8
    "11011100", -- 2269 - 0x8dd  :  220 - 0xdc
    "11001110", -- 2270 - 0x8de  :  206 - 0xce
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "01111000", -- 2272 - 0x8e0  :  120 - 0x78 -- Background 0x1c
    "11001100", -- 2273 - 0x8e1  :  204 - 0xcc
    "11000000", -- 2274 - 0x8e2  :  192 - 0xc0
    "01111100", -- 2275 - 0x8e3  :  124 - 0x7c
    "00000110", -- 2276 - 0x8e4  :    6 - 0x6
    "11000110", -- 2277 - 0x8e5  :  198 - 0xc6
    "01111100", -- 2278 - 0x8e6  :  124 - 0x7c
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "01111110", -- 2280 - 0x8e8  :  126 - 0x7e -- Background 0x1d
    "00011000", -- 2281 - 0x8e9  :   24 - 0x18
    "00011000", -- 2282 - 0x8ea  :   24 - 0x18
    "00011000", -- 2283 - 0x8eb  :   24 - 0x18
    "00011000", -- 2284 - 0x8ec  :   24 - 0x18
    "00011000", -- 2285 - 0x8ed  :   24 - 0x18
    "00011000", -- 2286 - 0x8ee  :   24 - 0x18
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "11000110", -- 2288 - 0x8f0  :  198 - 0xc6 -- Background 0x1e
    "11000110", -- 2289 - 0x8f1  :  198 - 0xc6
    "11000110", -- 2290 - 0x8f2  :  198 - 0xc6
    "11000110", -- 2291 - 0x8f3  :  198 - 0xc6
    "11000110", -- 2292 - 0x8f4  :  198 - 0xc6
    "11000110", -- 2293 - 0x8f5  :  198 - 0xc6
    "01111100", -- 2294 - 0x8f6  :  124 - 0x7c
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "11000110", -- 2296 - 0x8f8  :  198 - 0xc6 -- Background 0x1f
    "11000110", -- 2297 - 0x8f9  :  198 - 0xc6
    "11000110", -- 2298 - 0x8fa  :  198 - 0xc6
    "11101110", -- 2299 - 0x8fb  :  238 - 0xee
    "01111100", -- 2300 - 0x8fc  :  124 - 0x7c
    "00111000", -- 2301 - 0x8fd  :   56 - 0x38
    "00010000", -- 2302 - 0x8fe  :   16 - 0x10
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "11000110", -- 2304 - 0x900  :  198 - 0xc6 -- Background 0x20
    "11000110", -- 2305 - 0x901  :  198 - 0xc6
    "11010110", -- 2306 - 0x902  :  214 - 0xd6
    "11111110", -- 2307 - 0x903  :  254 - 0xfe
    "11111110", -- 2308 - 0x904  :  254 - 0xfe
    "11101110", -- 2309 - 0x905  :  238 - 0xee
    "11000110", -- 2310 - 0x906  :  198 - 0xc6
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "11000110", -- 2312 - 0x908  :  198 - 0xc6 -- Background 0x21
    "11101110", -- 2313 - 0x909  :  238 - 0xee
    "01111100", -- 2314 - 0x90a  :  124 - 0x7c
    "00111000", -- 2315 - 0x90b  :   56 - 0x38
    "01111100", -- 2316 - 0x90c  :  124 - 0x7c
    "11101110", -- 2317 - 0x90d  :  238 - 0xee
    "11000110", -- 2318 - 0x90e  :  198 - 0xc6
    "00000000", -- 2319 - 0x90f  :    0 - 0x0
    "01100110", -- 2320 - 0x910  :  102 - 0x66 -- Background 0x22
    "01100110", -- 2321 - 0x911  :  102 - 0x66
    "01100110", -- 2322 - 0x912  :  102 - 0x66
    "00111100", -- 2323 - 0x913  :   60 - 0x3c
    "00011000", -- 2324 - 0x914  :   24 - 0x18
    "00011000", -- 2325 - 0x915  :   24 - 0x18
    "00011000", -- 2326 - 0x916  :   24 - 0x18
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "11111110", -- 2328 - 0x918  :  254 - 0xfe -- Background 0x23
    "00001110", -- 2329 - 0x919  :   14 - 0xe
    "00011100", -- 2330 - 0x91a  :   28 - 0x1c
    "00111000", -- 2331 - 0x91b  :   56 - 0x38
    "01110000", -- 2332 - 0x91c  :  112 - 0x70
    "11100000", -- 2333 - 0x91d  :  224 - 0xe0
    "11111110", -- 2334 - 0x91e  :  254 - 0xfe
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Background 0x24
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "00000000", -- 2339 - 0x923  :    0 - 0x0
    "00000000", -- 2340 - 0x924  :    0 - 0x0
    "00000000", -- 2341 - 0x925  :    0 - 0x0
    "00000000", -- 2342 - 0x926  :    0 - 0x0
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "11111111", -- 2344 - 0x928  :  255 - 0xff -- Background 0x25
    "11111111", -- 2345 - 0x929  :  255 - 0xff
    "11111111", -- 2346 - 0x92a  :  255 - 0xff
    "11111111", -- 2347 - 0x92b  :  255 - 0xff
    "11111111", -- 2348 - 0x92c  :  255 - 0xff
    "11111111", -- 2349 - 0x92d  :  255 - 0xff
    "11111111", -- 2350 - 0x92e  :  255 - 0xff
    "11111111", -- 2351 - 0x92f  :  255 - 0xff
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "00000000", -- 2353 - 0x931  :    0 - 0x0
    "00000000", -- 2354 - 0x932  :    0 - 0x0
    "00000000", -- 2355 - 0x933  :    0 - 0x0
    "00000000", -- 2356 - 0x934  :    0 - 0x0
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "11111111", -- 2360 - 0x938  :  255 - 0xff -- Background 0x27
    "11111111", -- 2361 - 0x939  :  255 - 0xff
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "11111111", -- 2363 - 0x93b  :  255 - 0xff
    "11111111", -- 2364 - 0x93c  :  255 - 0xff
    "11111111", -- 2365 - 0x93d  :  255 - 0xff
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "11111111", -- 2367 - 0x93f  :  255 - 0xff
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "01111110", -- 2371 - 0x943  :  126 - 0x7e
    "01111110", -- 2372 - 0x944  :  126 - 0x7e
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- Background 0x29
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "01000100", -- 2378 - 0x94a  :   68 - 0x44
    "00101000", -- 2379 - 0x94b  :   40 - 0x28
    "00010000", -- 2380 - 0x94c  :   16 - 0x10
    "00101000", -- 2381 - 0x94d  :   40 - 0x28
    "01000100", -- 2382 - 0x94e  :   68 - 0x44
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "11111111", -- 2384 - 0x950  :  255 - 0xff -- Background 0x2a
    "11111111", -- 2385 - 0x951  :  255 - 0xff
    "11111111", -- 2386 - 0x952  :  255 - 0xff
    "11111111", -- 2387 - 0x953  :  255 - 0xff
    "11111111", -- 2388 - 0x954  :  255 - 0xff
    "11111111", -- 2389 - 0x955  :  255 - 0xff
    "11111111", -- 2390 - 0x956  :  255 - 0xff
    "11111111", -- 2391 - 0x957  :  255 - 0xff
    "00011000", -- 2392 - 0x958  :   24 - 0x18 -- Background 0x2b
    "00111100", -- 2393 - 0x959  :   60 - 0x3c
    "00111100", -- 2394 - 0x95a  :   60 - 0x3c
    "00111100", -- 2395 - 0x95b  :   60 - 0x3c
    "00011000", -- 2396 - 0x95c  :   24 - 0x18
    "00011000", -- 2397 - 0x95d  :   24 - 0x18
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00011000", -- 2399 - 0x95f  :   24 - 0x18
    "11111111", -- 2400 - 0x960  :  255 - 0xff -- Background 0x2c
    "01111111", -- 2401 - 0x961  :  127 - 0x7f
    "01111111", -- 2402 - 0x962  :  127 - 0x7f
    "01111111", -- 2403 - 0x963  :  127 - 0x7f
    "01111111", -- 2404 - 0x964  :  127 - 0x7f
    "11111111", -- 2405 - 0x965  :  255 - 0xff
    "11100011", -- 2406 - 0x966  :  227 - 0xe3
    "11000001", -- 2407 - 0x967  :  193 - 0xc1
    "10000000", -- 2408 - 0x968  :  128 - 0x80 -- Background 0x2d
    "10000000", -- 2409 - 0x969  :  128 - 0x80
    "10000000", -- 2410 - 0x96a  :  128 - 0x80
    "11000001", -- 2411 - 0x96b  :  193 - 0xc1
    "11100011", -- 2412 - 0x96c  :  227 - 0xe3
    "11111111", -- 2413 - 0x96d  :  255 - 0xff
    "11111111", -- 2414 - 0x96e  :  255 - 0xff
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00111000", -- 2416 - 0x970  :   56 - 0x38 -- Background 0x2e
    "01111100", -- 2417 - 0x971  :  124 - 0x7c
    "01111100", -- 2418 - 0x972  :  124 - 0x7c
    "01111100", -- 2419 - 0x973  :  124 - 0x7c
    "01111100", -- 2420 - 0x974  :  124 - 0x7c
    "01111100", -- 2421 - 0x975  :  124 - 0x7c
    "00111000", -- 2422 - 0x976  :   56 - 0x38
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000011", -- 2424 - 0x978  :    3 - 0x3 -- Background 0x2f
    "00000110", -- 2425 - 0x979  :    6 - 0x6
    "00001100", -- 2426 - 0x97a  :   12 - 0xc
    "00001100", -- 2427 - 0x97b  :   12 - 0xc
    "00001000", -- 2428 - 0x97c  :    8 - 0x8
    "00001000", -- 2429 - 0x97d  :    8 - 0x8
    "00000100", -- 2430 - 0x97e  :    4 - 0x4
    "00000011", -- 2431 - 0x97f  :    3 - 0x3
    "00000001", -- 2432 - 0x980  :    1 - 0x1 -- Background 0x30
    "00000010", -- 2433 - 0x981  :    2 - 0x2
    "00000100", -- 2434 - 0x982  :    4 - 0x4
    "00001000", -- 2435 - 0x983  :    8 - 0x8
    "00010000", -- 2436 - 0x984  :   16 - 0x10
    "00100000", -- 2437 - 0x985  :   32 - 0x20
    "01000000", -- 2438 - 0x986  :   64 - 0x40
    "10000000", -- 2439 - 0x987  :  128 - 0x80
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- Background 0x31
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000111", -- 2445 - 0x98d  :    7 - 0x7
    "00111000", -- 2446 - 0x98e  :   56 - 0x38
    "11000000", -- 2447 - 0x98f  :  192 - 0xc0
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Background 0x32
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "11100000", -- 2453 - 0x995  :  224 - 0xe0
    "00011100", -- 2454 - 0x996  :   28 - 0x1c
    "00000011", -- 2455 - 0x997  :    3 - 0x3
    "10000000", -- 2456 - 0x998  :  128 - 0x80 -- Background 0x33
    "01000000", -- 2457 - 0x999  :   64 - 0x40
    "00100000", -- 2458 - 0x99a  :   32 - 0x20
    "00010000", -- 2459 - 0x99b  :   16 - 0x10
    "00001000", -- 2460 - 0x99c  :    8 - 0x8
    "00000100", -- 2461 - 0x99d  :    4 - 0x4
    "00000010", -- 2462 - 0x99e  :    2 - 0x2
    "00000001", -- 2463 - 0x99f  :    1 - 0x1
    "00000100", -- 2464 - 0x9a0  :    4 - 0x4 -- Background 0x34
    "00001110", -- 2465 - 0x9a1  :   14 - 0xe
    "00001110", -- 2466 - 0x9a2  :   14 - 0xe
    "00001110", -- 2467 - 0x9a3  :   14 - 0xe
    "01101110", -- 2468 - 0x9a4  :  110 - 0x6e
    "01100100", -- 2469 - 0x9a5  :  100 - 0x64
    "01100000", -- 2470 - 0x9a6  :   96 - 0x60
    "01100000", -- 2471 - 0x9a7  :   96 - 0x60
    "00000111", -- 2472 - 0x9a8  :    7 - 0x7 -- Background 0x35
    "00001111", -- 2473 - 0x9a9  :   15 - 0xf
    "00011111", -- 2474 - 0x9aa  :   31 - 0x1f
    "00011111", -- 2475 - 0x9ab  :   31 - 0x1f
    "01111111", -- 2476 - 0x9ac  :  127 - 0x7f
    "11111111", -- 2477 - 0x9ad  :  255 - 0xff
    "11111111", -- 2478 - 0x9ae  :  255 - 0xff
    "01111111", -- 2479 - 0x9af  :  127 - 0x7f
    "00000011", -- 2480 - 0x9b0  :    3 - 0x3 -- Background 0x36
    "00000111", -- 2481 - 0x9b1  :    7 - 0x7
    "00011111", -- 2482 - 0x9b2  :   31 - 0x1f
    "00111111", -- 2483 - 0x9b3  :   63 - 0x3f
    "00111111", -- 2484 - 0x9b4  :   63 - 0x3f
    "00111111", -- 2485 - 0x9b5  :   63 - 0x3f
    "01111001", -- 2486 - 0x9b6  :  121 - 0x79
    "11110111", -- 2487 - 0x9b7  :  247 - 0xf7
    "11000000", -- 2488 - 0x9b8  :  192 - 0xc0 -- Background 0x37
    "11100000", -- 2489 - 0x9b9  :  224 - 0xe0
    "11110000", -- 2490 - 0x9ba  :  240 - 0xf0
    "11110100", -- 2491 - 0x9bb  :  244 - 0xf4
    "11111110", -- 2492 - 0x9bc  :  254 - 0xfe
    "10111111", -- 2493 - 0x9bd  :  191 - 0xbf
    "11011111", -- 2494 - 0x9be  :  223 - 0xdf
    "11111111", -- 2495 - 0x9bf  :  255 - 0xff
    "10010000", -- 2496 - 0x9c0  :  144 - 0x90 -- Background 0x38
    "10111000", -- 2497 - 0x9c1  :  184 - 0xb8
    "11111000", -- 2498 - 0x9c2  :  248 - 0xf8
    "11111010", -- 2499 - 0x9c3  :  250 - 0xfa
    "11111111", -- 2500 - 0x9c4  :  255 - 0xff
    "11111111", -- 2501 - 0x9c5  :  255 - 0xff
    "11111111", -- 2502 - 0x9c6  :  255 - 0xff
    "11111110", -- 2503 - 0x9c7  :  254 - 0xfe
    "00111011", -- 2504 - 0x9c8  :   59 - 0x3b -- Background 0x39
    "00011101", -- 2505 - 0x9c9  :   29 - 0x1d
    "00001110", -- 2506 - 0x9ca  :   14 - 0xe
    "00001111", -- 2507 - 0x9cb  :   15 - 0xf
    "00000111", -- 2508 - 0x9cc  :    7 - 0x7
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "11111111", -- 2512 - 0x9d0  :  255 - 0xff -- Background 0x3a
    "10111111", -- 2513 - 0x9d1  :  191 - 0xbf
    "00011100", -- 2514 - 0x9d2  :   28 - 0x1c
    "11000000", -- 2515 - 0x9d3  :  192 - 0xc0
    "11110011", -- 2516 - 0x9d4  :  243 - 0xf3
    "11111111", -- 2517 - 0x9d5  :  255 - 0xff
    "01111110", -- 2518 - 0x9d6  :  126 - 0x7e
    "00011100", -- 2519 - 0x9d7  :   28 - 0x1c
    "10111111", -- 2520 - 0x9d8  :  191 - 0xbf -- Background 0x3b
    "01111111", -- 2521 - 0x9d9  :  127 - 0x7f
    "00111101", -- 2522 - 0x9da  :   61 - 0x3d
    "10000011", -- 2523 - 0x9db  :  131 - 0x83
    "11000111", -- 2524 - 0x9dc  :  199 - 0xc7
    "11111111", -- 2525 - 0x9dd  :  255 - 0xff
    "11111111", -- 2526 - 0x9de  :  255 - 0xff
    "00111100", -- 2527 - 0x9df  :   60 - 0x3c
    "11111100", -- 2528 - 0x9e0  :  252 - 0xfc -- Background 0x3c
    "11111110", -- 2529 - 0x9e1  :  254 - 0xfe
    "11111111", -- 2530 - 0x9e2  :  255 - 0xff
    "11111110", -- 2531 - 0x9e3  :  254 - 0xfe
    "11111110", -- 2532 - 0x9e4  :  254 - 0xfe
    "11111000", -- 2533 - 0x9e5  :  248 - 0xf8
    "01100000", -- 2534 - 0x9e6  :   96 - 0x60
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "11000000", -- 2536 - 0x9e8  :  192 - 0xc0 -- Background 0x3d
    "00100000", -- 2537 - 0x9e9  :   32 - 0x20
    "00010000", -- 2538 - 0x9ea  :   16 - 0x10
    "00010000", -- 2539 - 0x9eb  :   16 - 0x10
    "00010000", -- 2540 - 0x9ec  :   16 - 0x10
    "00010000", -- 2541 - 0x9ed  :   16 - 0x10
    "00100000", -- 2542 - 0x9ee  :   32 - 0x20
    "11000000", -- 2543 - 0x9ef  :  192 - 0xc0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00111111", -- 2548 - 0x9f4  :   63 - 0x3f
    "01111111", -- 2549 - 0x9f5  :  127 - 0x7f
    "11100000", -- 2550 - 0x9f6  :  224 - 0xe0
    "11000000", -- 2551 - 0x9f7  :  192 - 0xc0
    "10001000", -- 2552 - 0x9f8  :  136 - 0x88 -- Background 0x3f
    "10011100", -- 2553 - 0x9f9  :  156 - 0x9c
    "10001000", -- 2554 - 0x9fa  :  136 - 0x88
    "10000000", -- 2555 - 0x9fb  :  128 - 0x80
    "10000000", -- 2556 - 0x9fc  :  128 - 0x80
    "10000000", -- 2557 - 0x9fd  :  128 - 0x80
    "10000000", -- 2558 - 0x9fe  :  128 - 0x80
    "10000000", -- 2559 - 0x9ff  :  128 - 0x80
    "11111110", -- 2560 - 0xa00  :  254 - 0xfe -- Background 0x40
    "11111110", -- 2561 - 0xa01  :  254 - 0xfe
    "11111110", -- 2562 - 0xa02  :  254 - 0xfe
    "11111110", -- 2563 - 0xa03  :  254 - 0xfe
    "11111110", -- 2564 - 0xa04  :  254 - 0xfe
    "11111110", -- 2565 - 0xa05  :  254 - 0xfe
    "11111110", -- 2566 - 0xa06  :  254 - 0xfe
    "11111110", -- 2567 - 0xa07  :  254 - 0xfe
    "00001000", -- 2568 - 0xa08  :    8 - 0x8 -- Background 0x41
    "00010100", -- 2569 - 0xa09  :   20 - 0x14
    "00100100", -- 2570 - 0xa0a  :   36 - 0x24
    "11000100", -- 2571 - 0xa0b  :  196 - 0xc4
    "00000011", -- 2572 - 0xa0c  :    3 - 0x3
    "01000000", -- 2573 - 0xa0d  :   64 - 0x40
    "10100001", -- 2574 - 0xa0e  :  161 - 0xa1
    "00100110", -- 2575 - 0xa0f  :   38 - 0x26
    "11111111", -- 2576 - 0xa10  :  255 - 0xff -- Background 0x42
    "11111111", -- 2577 - 0xa11  :  255 - 0xff
    "11111111", -- 2578 - 0xa12  :  255 - 0xff
    "11111111", -- 2579 - 0xa13  :  255 - 0xff
    "01111111", -- 2580 - 0xa14  :  127 - 0x7f
    "01111111", -- 2581 - 0xa15  :  127 - 0x7f
    "01111111", -- 2582 - 0xa16  :  127 - 0x7f
    "01111111", -- 2583 - 0xa17  :  127 - 0x7f
    "11111111", -- 2584 - 0xa18  :  255 - 0xff -- Background 0x43
    "11111111", -- 2585 - 0xa19  :  255 - 0xff
    "11111111", -- 2586 - 0xa1a  :  255 - 0xff
    "11111111", -- 2587 - 0xa1b  :  255 - 0xff
    "11111111", -- 2588 - 0xa1c  :  255 - 0xff
    "11111111", -- 2589 - 0xa1d  :  255 - 0xff
    "11111111", -- 2590 - 0xa1e  :  255 - 0xff
    "11111111", -- 2591 - 0xa1f  :  255 - 0xff
    "01111111", -- 2592 - 0xa20  :  127 - 0x7f -- Background 0x44
    "10000000", -- 2593 - 0xa21  :  128 - 0x80
    "10000000", -- 2594 - 0xa22  :  128 - 0x80
    "10011000", -- 2595 - 0xa23  :  152 - 0x98
    "10011100", -- 2596 - 0xa24  :  156 - 0x9c
    "10001100", -- 2597 - 0xa25  :  140 - 0x8c
    "10000000", -- 2598 - 0xa26  :  128 - 0x80
    "10000000", -- 2599 - 0xa27  :  128 - 0x80
    "11111111", -- 2600 - 0xa28  :  255 - 0xff -- Background 0x45
    "00000001", -- 2601 - 0xa29  :    1 - 0x1
    "00000001", -- 2602 - 0xa2a  :    1 - 0x1
    "11111111", -- 2603 - 0xa2b  :  255 - 0xff
    "00010000", -- 2604 - 0xa2c  :   16 - 0x10
    "00010000", -- 2605 - 0xa2d  :   16 - 0x10
    "00010000", -- 2606 - 0xa2e  :   16 - 0x10
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "10000000", -- 2608 - 0xa30  :  128 - 0x80 -- Background 0x46
    "10000000", -- 2609 - 0xa31  :  128 - 0x80
    "10000000", -- 2610 - 0xa32  :  128 - 0x80
    "10000000", -- 2611 - 0xa33  :  128 - 0x80
    "10000000", -- 2612 - 0xa34  :  128 - 0x80
    "10000000", -- 2613 - 0xa35  :  128 - 0x80
    "10000000", -- 2614 - 0xa36  :  128 - 0x80
    "10000000", -- 2615 - 0xa37  :  128 - 0x80
    "00000001", -- 2616 - 0xa38  :    1 - 0x1 -- Background 0x47
    "00000001", -- 2617 - 0xa39  :    1 - 0x1
    "00000001", -- 2618 - 0xa3a  :    1 - 0x1
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "00010000", -- 2620 - 0xa3c  :   16 - 0x10
    "00010000", -- 2621 - 0xa3d  :   16 - 0x10
    "00010000", -- 2622 - 0xa3e  :   16 - 0x10
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "11111111", -- 2624 - 0xa40  :  255 - 0xff -- Background 0x48
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "11111110", -- 2632 - 0xa48  :  254 - 0xfe -- Background 0x49
    "00000001", -- 2633 - 0xa49  :    1 - 0x1
    "00000001", -- 2634 - 0xa4a  :    1 - 0x1
    "00011001", -- 2635 - 0xa4b  :   25 - 0x19
    "00011101", -- 2636 - 0xa4c  :   29 - 0x1d
    "00001101", -- 2637 - 0xa4d  :   13 - 0xd
    "00000001", -- 2638 - 0xa4e  :    1 - 0x1
    "00000001", -- 2639 - 0xa4f  :    1 - 0x1
    "00000001", -- 2640 - 0xa50  :    1 - 0x1 -- Background 0x4a
    "00000001", -- 2641 - 0xa51  :    1 - 0x1
    "00000001", -- 2642 - 0xa52  :    1 - 0x1
    "00000001", -- 2643 - 0xa53  :    1 - 0x1
    "00000001", -- 2644 - 0xa54  :    1 - 0x1
    "00000001", -- 2645 - 0xa55  :    1 - 0x1
    "00000001", -- 2646 - 0xa56  :    1 - 0x1
    "00000001", -- 2647 - 0xa57  :    1 - 0x1
    "00111111", -- 2648 - 0xa58  :   63 - 0x3f -- Background 0x4b
    "01111111", -- 2649 - 0xa59  :  127 - 0x7f
    "01111111", -- 2650 - 0xa5a  :  127 - 0x7f
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "11111111", -- 2652 - 0xa5c  :  255 - 0xff
    "11111111", -- 2653 - 0xa5d  :  255 - 0xff
    "11111111", -- 2654 - 0xa5e  :  255 - 0xff
    "11111111", -- 2655 - 0xa5f  :  255 - 0xff
    "11111111", -- 2656 - 0xa60  :  255 - 0xff -- Background 0x4c
    "11111111", -- 2657 - 0xa61  :  255 - 0xff
    "11111111", -- 2658 - 0xa62  :  255 - 0xff
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "11111111", -- 2660 - 0xa64  :  255 - 0xff
    "11111111", -- 2661 - 0xa65  :  255 - 0xff
    "01111110", -- 2662 - 0xa66  :  126 - 0x7e
    "00111100", -- 2663 - 0xa67  :   60 - 0x3c
    "11111111", -- 2664 - 0xa68  :  255 - 0xff -- Background 0x4d
    "11111111", -- 2665 - 0xa69  :  255 - 0xff
    "11111111", -- 2666 - 0xa6a  :  255 - 0xff
    "11111111", -- 2667 - 0xa6b  :  255 - 0xff
    "11111111", -- 2668 - 0xa6c  :  255 - 0xff
    "11111111", -- 2669 - 0xa6d  :  255 - 0xff
    "11111111", -- 2670 - 0xa6e  :  255 - 0xff
    "11111111", -- 2671 - 0xa6f  :  255 - 0xff
    "11111111", -- 2672 - 0xa70  :  255 - 0xff -- Background 0x4e
    "11111111", -- 2673 - 0xa71  :  255 - 0xff
    "11111111", -- 2674 - 0xa72  :  255 - 0xff
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111111", -- 2676 - 0xa74  :  255 - 0xff
    "11111111", -- 2677 - 0xa75  :  255 - 0xff
    "11111110", -- 2678 - 0xa76  :  254 - 0xfe
    "01111100", -- 2679 - 0xa77  :  124 - 0x7c
    "11111111", -- 2680 - 0xa78  :  255 - 0xff -- Background 0x4f
    "11111111", -- 2681 - 0xa79  :  255 - 0xff
    "11111111", -- 2682 - 0xa7a  :  255 - 0xff
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111111", -- 2684 - 0xa7c  :  255 - 0xff
    "11111111", -- 2685 - 0xa7d  :  255 - 0xff
    "11111110", -- 2686 - 0xa7e  :  254 - 0xfe
    "01111100", -- 2687 - 0xa7f  :  124 - 0x7c
    "11111000", -- 2688 - 0xa80  :  248 - 0xf8 -- Background 0x50
    "11111100", -- 2689 - 0xa81  :  252 - 0xfc
    "11111110", -- 2690 - 0xa82  :  254 - 0xfe
    "11111110", -- 2691 - 0xa83  :  254 - 0xfe
    "11111111", -- 2692 - 0xa84  :  255 - 0xff
    "11111111", -- 2693 - 0xa85  :  255 - 0xff
    "11111111", -- 2694 - 0xa86  :  255 - 0xff
    "11111111", -- 2695 - 0xa87  :  255 - 0xff
    "11111111", -- 2696 - 0xa88  :  255 - 0xff -- Background 0x51
    "11111111", -- 2697 - 0xa89  :  255 - 0xff
    "11111111", -- 2698 - 0xa8a  :  255 - 0xff
    "11111111", -- 2699 - 0xa8b  :  255 - 0xff
    "11111111", -- 2700 - 0xa8c  :  255 - 0xff
    "11111111", -- 2701 - 0xa8d  :  255 - 0xff
    "01111110", -- 2702 - 0xa8e  :  126 - 0x7e
    "00111100", -- 2703 - 0xa8f  :   60 - 0x3c
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00001000", -- 2705 - 0xa91  :    8 - 0x8
    "00001000", -- 2706 - 0xa92  :    8 - 0x8
    "00001000", -- 2707 - 0xa93  :    8 - 0x8
    "00010000", -- 2708 - 0xa94  :   16 - 0x10
    "00010000", -- 2709 - 0xa95  :   16 - 0x10
    "00010000", -- 2710 - 0xa96  :   16 - 0x10
    "00000000", -- 2711 - 0xa97  :    0 - 0x0
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- Background 0x53
    "01111111", -- 2713 - 0xa99  :  127 - 0x7f
    "01111111", -- 2714 - 0xa9a  :  127 - 0x7f
    "01111000", -- 2715 - 0xa9b  :  120 - 0x78
    "01110011", -- 2716 - 0xa9c  :  115 - 0x73
    "01110011", -- 2717 - 0xa9d  :  115 - 0x73
    "01110011", -- 2718 - 0xa9e  :  115 - 0x73
    "01111111", -- 2719 - 0xa9f  :  127 - 0x7f
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Background 0x54
    "11111111", -- 2721 - 0xaa1  :  255 - 0xff
    "11111111", -- 2722 - 0xaa2  :  255 - 0xff
    "00111111", -- 2723 - 0xaa3  :   63 - 0x3f
    "10011111", -- 2724 - 0xaa4  :  159 - 0x9f
    "10011111", -- 2725 - 0xaa5  :  159 - 0x9f
    "10011111", -- 2726 - 0xaa6  :  159 - 0x9f
    "00011111", -- 2727 - 0xaa7  :   31 - 0x1f
    "01111110", -- 2728 - 0xaa8  :  126 - 0x7e -- Background 0x55
    "01111110", -- 2729 - 0xaa9  :  126 - 0x7e
    "01111111", -- 2730 - 0xaaa  :  127 - 0x7f
    "01111110", -- 2731 - 0xaab  :  126 - 0x7e
    "01111110", -- 2732 - 0xaac  :  126 - 0x7e
    "01111111", -- 2733 - 0xaad  :  127 - 0x7f
    "01111111", -- 2734 - 0xaae  :  127 - 0x7f
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "01111111", -- 2736 - 0xab0  :  127 - 0x7f -- Background 0x56
    "01111111", -- 2737 - 0xab1  :  127 - 0x7f
    "11111111", -- 2738 - 0xab2  :  255 - 0xff
    "01111111", -- 2739 - 0xab3  :  127 - 0x7f
    "01111111", -- 2740 - 0xab4  :  127 - 0x7f
    "11111111", -- 2741 - 0xab5  :  255 - 0xff
    "11111111", -- 2742 - 0xab6  :  255 - 0xff
    "11111111", -- 2743 - 0xab7  :  255 - 0xff
    "01111111", -- 2744 - 0xab8  :  127 - 0x7f -- Background 0x57
    "10000000", -- 2745 - 0xab9  :  128 - 0x80
    "10100000", -- 2746 - 0xaba  :  160 - 0xa0
    "10000000", -- 2747 - 0xabb  :  128 - 0x80
    "10000000", -- 2748 - 0xabc  :  128 - 0x80
    "10000000", -- 2749 - 0xabd  :  128 - 0x80
    "10000000", -- 2750 - 0xabe  :  128 - 0x80
    "10000000", -- 2751 - 0xabf  :  128 - 0x80
    "11111110", -- 2752 - 0xac0  :  254 - 0xfe -- Background 0x58
    "00000001", -- 2753 - 0xac1  :    1 - 0x1
    "00000101", -- 2754 - 0xac2  :    5 - 0x5
    "00000001", -- 2755 - 0xac3  :    1 - 0x1
    "00000001", -- 2756 - 0xac4  :    1 - 0x1
    "00000001", -- 2757 - 0xac5  :    1 - 0x1
    "00000001", -- 2758 - 0xac6  :    1 - 0x1
    "00000001", -- 2759 - 0xac7  :    1 - 0x1
    "10000000", -- 2760 - 0xac8  :  128 - 0x80 -- Background 0x59
    "10000000", -- 2761 - 0xac9  :  128 - 0x80
    "10000000", -- 2762 - 0xaca  :  128 - 0x80
    "10000000", -- 2763 - 0xacb  :  128 - 0x80
    "10000000", -- 2764 - 0xacc  :  128 - 0x80
    "10100000", -- 2765 - 0xacd  :  160 - 0xa0
    "10000000", -- 2766 - 0xace  :  128 - 0x80
    "01111111", -- 2767 - 0xacf  :  127 - 0x7f
    "00000001", -- 2768 - 0xad0  :    1 - 0x1 -- Background 0x5a
    "00000001", -- 2769 - 0xad1  :    1 - 0x1
    "00000001", -- 2770 - 0xad2  :    1 - 0x1
    "00000001", -- 2771 - 0xad3  :    1 - 0x1
    "00000001", -- 2772 - 0xad4  :    1 - 0x1
    "00000101", -- 2773 - 0xad5  :    5 - 0x5
    "00000001", -- 2774 - 0xad6  :    1 - 0x1
    "11111110", -- 2775 - 0xad7  :  254 - 0xfe
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "11111100", -- 2780 - 0xadc  :  252 - 0xfc
    "11111110", -- 2781 - 0xadd  :  254 - 0xfe
    "00000111", -- 2782 - 0xade  :    7 - 0x7
    "00000011", -- 2783 - 0xadf  :    3 - 0x3
    "00010001", -- 2784 - 0xae0  :   17 - 0x11 -- Background 0x5c
    "00111001", -- 2785 - 0xae1  :   57 - 0x39
    "00010001", -- 2786 - 0xae2  :   17 - 0x11
    "00000001", -- 2787 - 0xae3  :    1 - 0x1
    "00000001", -- 2788 - 0xae4  :    1 - 0x1
    "00000001", -- 2789 - 0xae5  :    1 - 0x1
    "00000001", -- 2790 - 0xae6  :    1 - 0x1
    "00000001", -- 2791 - 0xae7  :    1 - 0x1
    "11101111", -- 2792 - 0xae8  :  239 - 0xef -- Background 0x5d
    "00101000", -- 2793 - 0xae9  :   40 - 0x28
    "00101000", -- 2794 - 0xaea  :   40 - 0x28
    "00101000", -- 2795 - 0xaeb  :   40 - 0x28
    "00101000", -- 2796 - 0xaec  :   40 - 0x28
    "00101000", -- 2797 - 0xaed  :   40 - 0x28
    "11101111", -- 2798 - 0xaee  :  239 - 0xef
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "11111110", -- 2800 - 0xaf0  :  254 - 0xfe -- Background 0x5e
    "10000010", -- 2801 - 0xaf1  :  130 - 0x82
    "10000010", -- 2802 - 0xaf2  :  130 - 0x82
    "10000010", -- 2803 - 0xaf3  :  130 - 0x82
    "10000010", -- 2804 - 0xaf4  :  130 - 0x82
    "10000010", -- 2805 - 0xaf5  :  130 - 0x82
    "11111110", -- 2806 - 0xaf6  :  254 - 0xfe
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "10000000", -- 2808 - 0xaf8  :  128 - 0x80 -- Background 0x5f
    "10000000", -- 2809 - 0xaf9  :  128 - 0x80
    "10000000", -- 2810 - 0xafa  :  128 - 0x80
    "10011000", -- 2811 - 0xafb  :  152 - 0x98
    "10011100", -- 2812 - 0xafc  :  156 - 0x9c
    "10001100", -- 2813 - 0xafd  :  140 - 0x8c
    "10000000", -- 2814 - 0xafe  :  128 - 0x80
    "01111111", -- 2815 - 0xaff  :  127 - 0x7f
    "11111111", -- 2816 - 0xb00  :  255 - 0xff -- Background 0x60
    "11111111", -- 2817 - 0xb01  :  255 - 0xff
    "10000011", -- 2818 - 0xb02  :  131 - 0x83
    "11110011", -- 2819 - 0xb03  :  243 - 0xf3
    "11110011", -- 2820 - 0xb04  :  243 - 0xf3
    "11110011", -- 2821 - 0xb05  :  243 - 0xf3
    "11110011", -- 2822 - 0xb06  :  243 - 0xf3
    "11110011", -- 2823 - 0xb07  :  243 - 0xf3
    "11111111", -- 2824 - 0xb08  :  255 - 0xff -- Background 0x61
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11110000", -- 2826 - 0xb0a  :  240 - 0xf0
    "11110110", -- 2827 - 0xb0b  :  246 - 0xf6
    "11110110", -- 2828 - 0xb0c  :  246 - 0xf6
    "11110110", -- 2829 - 0xb0d  :  246 - 0xf6
    "11110110", -- 2830 - 0xb0e  :  246 - 0xf6
    "11110110", -- 2831 - 0xb0f  :  246 - 0xf6
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Background 0x62
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "00000000", -- 2834 - 0xb12  :    0 - 0x0
    "00000000", -- 2835 - 0xb13  :    0 - 0x0
    "00000000", -- 2836 - 0xb14  :    0 - 0x0
    "00000000", -- 2837 - 0xb15  :    0 - 0x0
    "00000000", -- 2838 - 0xb16  :    0 - 0x0
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "11111111", -- 2840 - 0xb18  :  255 - 0xff -- Background 0x63
    "11111111", -- 2841 - 0xb19  :  255 - 0xff
    "00000001", -- 2842 - 0xb1a  :    1 - 0x1
    "01010111", -- 2843 - 0xb1b  :   87 - 0x57
    "00101111", -- 2844 - 0xb1c  :   47 - 0x2f
    "01010111", -- 2845 - 0xb1d  :   87 - 0x57
    "00101111", -- 2846 - 0xb1e  :   47 - 0x2f
    "01010111", -- 2847 - 0xb1f  :   87 - 0x57
    "11110011", -- 2848 - 0xb20  :  243 - 0xf3 -- Background 0x64
    "11110011", -- 2849 - 0xb21  :  243 - 0xf3
    "11110011", -- 2850 - 0xb22  :  243 - 0xf3
    "11110011", -- 2851 - 0xb23  :  243 - 0xf3
    "11110011", -- 2852 - 0xb24  :  243 - 0xf3
    "11110011", -- 2853 - 0xb25  :  243 - 0xf3
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "00111111", -- 2855 - 0xb27  :   63 - 0x3f
    "11110110", -- 2856 - 0xb28  :  246 - 0xf6 -- Background 0x65
    "11110110", -- 2857 - 0xb29  :  246 - 0xf6
    "11110110", -- 2858 - 0xb2a  :  246 - 0xf6
    "11110110", -- 2859 - 0xb2b  :  246 - 0xf6
    "11110110", -- 2860 - 0xb2c  :  246 - 0xf6
    "11110110", -- 2861 - 0xb2d  :  246 - 0xf6
    "11111111", -- 2862 - 0xb2e  :  255 - 0xff
    "11111111", -- 2863 - 0xb2f  :  255 - 0xff
    "00000000", -- 2864 - 0xb30  :    0 - 0x0 -- Background 0x66
    "00000000", -- 2865 - 0xb31  :    0 - 0x0
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "00000000", -- 2867 - 0xb33  :    0 - 0x0
    "00000000", -- 2868 - 0xb34  :    0 - 0x0
    "00000000", -- 2869 - 0xb35  :    0 - 0x0
    "11111111", -- 2870 - 0xb36  :  255 - 0xff
    "11111111", -- 2871 - 0xb37  :  255 - 0xff
    "00101111", -- 2872 - 0xb38  :   47 - 0x2f -- Background 0x67
    "01010111", -- 2873 - 0xb39  :   87 - 0x57
    "00101111", -- 2874 - 0xb3a  :   47 - 0x2f
    "01010111", -- 2875 - 0xb3b  :   87 - 0x57
    "00101111", -- 2876 - 0xb3c  :   47 - 0x2f
    "01010111", -- 2877 - 0xb3d  :   87 - 0x57
    "11111111", -- 2878 - 0xb3e  :  255 - 0xff
    "11111100", -- 2879 - 0xb3f  :  252 - 0xfc
    "00111100", -- 2880 - 0xb40  :   60 - 0x3c -- Background 0x68
    "00111100", -- 2881 - 0xb41  :   60 - 0x3c
    "00111100", -- 2882 - 0xb42  :   60 - 0x3c
    "00111100", -- 2883 - 0xb43  :   60 - 0x3c
    "00111100", -- 2884 - 0xb44  :   60 - 0x3c
    "00111100", -- 2885 - 0xb45  :   60 - 0x3c
    "00111100", -- 2886 - 0xb46  :   60 - 0x3c
    "00111100", -- 2887 - 0xb47  :   60 - 0x3c
    "11111011", -- 2888 - 0xb48  :  251 - 0xfb -- Background 0x69
    "11111011", -- 2889 - 0xb49  :  251 - 0xfb
    "11111011", -- 2890 - 0xb4a  :  251 - 0xfb
    "11111011", -- 2891 - 0xb4b  :  251 - 0xfb
    "11111011", -- 2892 - 0xb4c  :  251 - 0xfb
    "11111011", -- 2893 - 0xb4d  :  251 - 0xfb
    "11111011", -- 2894 - 0xb4e  :  251 - 0xfb
    "11111011", -- 2895 - 0xb4f  :  251 - 0xfb
    "10111100", -- 2896 - 0xb50  :  188 - 0xbc -- Background 0x6a
    "01011100", -- 2897 - 0xb51  :   92 - 0x5c
    "10111100", -- 2898 - 0xb52  :  188 - 0xbc
    "01011100", -- 2899 - 0xb53  :   92 - 0x5c
    "10111100", -- 2900 - 0xb54  :  188 - 0xbc
    "01011100", -- 2901 - 0xb55  :   92 - 0x5c
    "10111100", -- 2902 - 0xb56  :  188 - 0xbc
    "01011100", -- 2903 - 0xb57  :   92 - 0x5c
    "00011111", -- 2904 - 0xb58  :   31 - 0x1f -- Background 0x6b
    "00100000", -- 2905 - 0xb59  :   32 - 0x20
    "01000000", -- 2906 - 0xb5a  :   64 - 0x40
    "01000000", -- 2907 - 0xb5b  :   64 - 0x40
    "10000000", -- 2908 - 0xb5c  :  128 - 0x80
    "10000000", -- 2909 - 0xb5d  :  128 - 0x80
    "10000000", -- 2910 - 0xb5e  :  128 - 0x80
    "10000001", -- 2911 - 0xb5f  :  129 - 0x81
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Background 0x6c
    "10000000", -- 2913 - 0xb61  :  128 - 0x80
    "10000000", -- 2914 - 0xb62  :  128 - 0x80
    "11000000", -- 2915 - 0xb63  :  192 - 0xc0
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11111111", -- 2917 - 0xb65  :  255 - 0xff
    "11111110", -- 2918 - 0xb66  :  254 - 0xfe
    "11111110", -- 2919 - 0xb67  :  254 - 0xfe
    "11111111", -- 2920 - 0xb68  :  255 - 0xff -- Background 0x6d
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "01111111", -- 2922 - 0xb6a  :  127 - 0x7f
    "11111111", -- 2923 - 0xb6b  :  255 - 0xff
    "11111111", -- 2924 - 0xb6c  :  255 - 0xff
    "00000111", -- 2925 - 0xb6d  :    7 - 0x7
    "00000011", -- 2926 - 0xb6e  :    3 - 0x3
    "00000011", -- 2927 - 0xb6f  :    3 - 0x3
    "11111111", -- 2928 - 0xb70  :  255 - 0xff -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "10000001", -- 2933 - 0xb75  :  129 - 0x81
    "11000011", -- 2934 - 0xb76  :  195 - 0xc3
    "11111111", -- 2935 - 0xb77  :  255 - 0xff
    "11111000", -- 2936 - 0xb78  :  248 - 0xf8 -- Background 0x6f
    "11111100", -- 2937 - 0xb79  :  252 - 0xfc
    "11111110", -- 2938 - 0xb7a  :  254 - 0xfe
    "11111110", -- 2939 - 0xb7b  :  254 - 0xfe
    "11100011", -- 2940 - 0xb7c  :  227 - 0xe3
    "11000001", -- 2941 - 0xb7d  :  193 - 0xc1
    "10000001", -- 2942 - 0xb7e  :  129 - 0x81
    "10000001", -- 2943 - 0xb7f  :  129 - 0x81
    "10000011", -- 2944 - 0xb80  :  131 - 0x83 -- Background 0x70
    "11111111", -- 2945 - 0xb81  :  255 - 0xff
    "11111111", -- 2946 - 0xb82  :  255 - 0xff
    "11111111", -- 2947 - 0xb83  :  255 - 0xff
    "11111111", -- 2948 - 0xb84  :  255 - 0xff
    "11111111", -- 2949 - 0xb85  :  255 - 0xff
    "01111111", -- 2950 - 0xb86  :  127 - 0x7f
    "00011111", -- 2951 - 0xb87  :   31 - 0x1f
    "11111100", -- 2952 - 0xb88  :  252 - 0xfc -- Background 0x71
    "11111100", -- 2953 - 0xb89  :  252 - 0xfc
    "11111100", -- 2954 - 0xb8a  :  252 - 0xfc
    "11111100", -- 2955 - 0xb8b  :  252 - 0xfc
    "11111110", -- 2956 - 0xb8c  :  254 - 0xfe
    "11111110", -- 2957 - 0xb8d  :  254 - 0xfe
    "11111111", -- 2958 - 0xb8e  :  255 - 0xff
    "11111111", -- 2959 - 0xb8f  :  255 - 0xff
    "00000001", -- 2960 - 0xb90  :    1 - 0x1 -- Background 0x72
    "00000001", -- 2961 - 0xb91  :    1 - 0x1
    "00000001", -- 2962 - 0xb92  :    1 - 0x1
    "00000001", -- 2963 - 0xb93  :    1 - 0x1
    "00000011", -- 2964 - 0xb94  :    3 - 0x3
    "00000011", -- 2965 - 0xb95  :    3 - 0x3
    "00000111", -- 2966 - 0xb96  :    7 - 0x7
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "11111111", -- 2968 - 0xb98  :  255 - 0xff -- Background 0x73
    "11111111", -- 2969 - 0xb99  :  255 - 0xff
    "11111111", -- 2970 - 0xb9a  :  255 - 0xff
    "11111111", -- 2971 - 0xb9b  :  255 - 0xff
    "11111111", -- 2972 - 0xb9c  :  255 - 0xff
    "11111111", -- 2973 - 0xb9d  :  255 - 0xff
    "11111111", -- 2974 - 0xb9e  :  255 - 0xff
    "11111111", -- 2975 - 0xb9f  :  255 - 0xff
    "10000001", -- 2976 - 0xba0  :  129 - 0x81 -- Background 0x74
    "11000001", -- 2977 - 0xba1  :  193 - 0xc1
    "11100011", -- 2978 - 0xba2  :  227 - 0xe3
    "11111111", -- 2979 - 0xba3  :  255 - 0xff
    "11111111", -- 2980 - 0xba4  :  255 - 0xff
    "11111111", -- 2981 - 0xba5  :  255 - 0xff
    "11111111", -- 2982 - 0xba6  :  255 - 0xff
    "11111110", -- 2983 - 0xba7  :  254 - 0xfe
    "11111111", -- 2984 - 0xba8  :  255 - 0xff -- Background 0x75
    "11111111", -- 2985 - 0xba9  :  255 - 0xff
    "11111111", -- 2986 - 0xbaa  :  255 - 0xff
    "11111111", -- 2987 - 0xbab  :  255 - 0xff
    "11111111", -- 2988 - 0xbac  :  255 - 0xff
    "11111011", -- 2989 - 0xbad  :  251 - 0xfb
    "10110101", -- 2990 - 0xbae  :  181 - 0xb5
    "11001110", -- 2991 - 0xbaf  :  206 - 0xce
    "11111111", -- 2992 - 0xbb0  :  255 - 0xff -- Background 0x76
    "11111111", -- 2993 - 0xbb1  :  255 - 0xff
    "11111111", -- 2994 - 0xbb2  :  255 - 0xff
    "11111111", -- 2995 - 0xbb3  :  255 - 0xff
    "11111111", -- 2996 - 0xbb4  :  255 - 0xff
    "11011111", -- 2997 - 0xbb5  :  223 - 0xdf
    "10101101", -- 2998 - 0xbb6  :  173 - 0xad
    "01110011", -- 2999 - 0xbb7  :  115 - 0x73
    "01110111", -- 3000 - 0xbb8  :  119 - 0x77 -- Background 0x77
    "01110111", -- 3001 - 0xbb9  :  119 - 0x77
    "01110111", -- 3002 - 0xbba  :  119 - 0x77
    "01110111", -- 3003 - 0xbbb  :  119 - 0x77
    "01110111", -- 3004 - 0xbbc  :  119 - 0x77
    "01110111", -- 3005 - 0xbbd  :  119 - 0x77
    "01110111", -- 3006 - 0xbbe  :  119 - 0x77
    "01110111", -- 3007 - 0xbbf  :  119 - 0x77
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "11111111", -- 3015 - 0xbc7  :  255 - 0xff
    "01110111", -- 3016 - 0xbc8  :  119 - 0x77 -- Background 0x79
    "01110111", -- 3017 - 0xbc9  :  119 - 0x77
    "01110111", -- 3018 - 0xbca  :  119 - 0x77
    "01110111", -- 3019 - 0xbcb  :  119 - 0x77
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000001", -- 3024 - 0xbd0  :    1 - 0x1 -- Background 0x7a
    "00000001", -- 3025 - 0xbd1  :    1 - 0x1
    "00000001", -- 3026 - 0xbd2  :    1 - 0x1
    "00011001", -- 3027 - 0xbd3  :   25 - 0x19
    "00011101", -- 3028 - 0xbd4  :   29 - 0x1d
    "00001101", -- 3029 - 0xbd5  :   13 - 0xd
    "00000001", -- 3030 - 0xbd6  :    1 - 0x1
    "11111110", -- 3031 - 0xbd7  :  254 - 0xfe
    "00100000", -- 3032 - 0xbd8  :   32 - 0x20 -- Background 0x7b
    "01111000", -- 3033 - 0xbd9  :  120 - 0x78
    "01111111", -- 3034 - 0xbda  :  127 - 0x7f
    "11111110", -- 3035 - 0xbdb  :  254 - 0xfe
    "11111110", -- 3036 - 0xbdc  :  254 - 0xfe
    "11111110", -- 3037 - 0xbdd  :  254 - 0xfe
    "11111110", -- 3038 - 0xbde  :  254 - 0xfe
    "11111110", -- 3039 - 0xbdf  :  254 - 0xfe
    "00000100", -- 3040 - 0xbe0  :    4 - 0x4 -- Background 0x7c
    "10011010", -- 3041 - 0xbe1  :  154 - 0x9a
    "11111010", -- 3042 - 0xbe2  :  250 - 0xfa
    "11111101", -- 3043 - 0xbe3  :  253 - 0xfd
    "11111101", -- 3044 - 0xbe4  :  253 - 0xfd
    "11111101", -- 3045 - 0xbe5  :  253 - 0xfd
    "11111101", -- 3046 - 0xbe6  :  253 - 0xfd
    "11111101", -- 3047 - 0xbe7  :  253 - 0xfd
    "01111110", -- 3048 - 0xbe8  :  126 - 0x7e -- Background 0x7d
    "00111000", -- 3049 - 0xbe9  :   56 - 0x38
    "00100001", -- 3050 - 0xbea  :   33 - 0x21
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000001", -- 3052 - 0xbec  :    1 - 0x1
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000001", -- 3054 - 0xbee  :    1 - 0x1
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "11111010", -- 3056 - 0xbf0  :  250 - 0xfa -- Background 0x7e
    "10001010", -- 3057 - 0xbf1  :  138 - 0x8a
    "10000100", -- 3058 - 0xbf2  :  132 - 0x84
    "10000000", -- 3059 - 0xbf3  :  128 - 0x80
    "10000000", -- 3060 - 0xbf4  :  128 - 0x80
    "10000000", -- 3061 - 0xbf5  :  128 - 0x80
    "10000000", -- 3062 - 0xbf6  :  128 - 0x80
    "10000000", -- 3063 - 0xbf7  :  128 - 0x80
    "00000010", -- 3064 - 0xbf8  :    2 - 0x2 -- Background 0x7f
    "00000100", -- 3065 - 0xbf9  :    4 - 0x4
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00010000", -- 3067 - 0xbfb  :   16 - 0x10
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "01000000", -- 3069 - 0xbfd  :   64 - 0x40
    "10000000", -- 3070 - 0xbfe  :  128 - 0x80
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00001011", -- 3072 - 0xc00  :   11 - 0xb -- Background 0x80
    "00001011", -- 3073 - 0xc01  :   11 - 0xb
    "00111011", -- 3074 - 0xc02  :   59 - 0x3b
    "00001011", -- 3075 - 0xc03  :   11 - 0xb
    "11111011", -- 3076 - 0xc04  :  251 - 0xfb
    "00001011", -- 3077 - 0xc05  :   11 - 0xb
    "00001011", -- 3078 - 0xc06  :   11 - 0xb
    "00001010", -- 3079 - 0xc07  :   10 - 0xa
    "10010000", -- 3080 - 0xc08  :  144 - 0x90 -- Background 0x81
    "00010000", -- 3081 - 0xc09  :   16 - 0x10
    "00011111", -- 3082 - 0xc0a  :   31 - 0x1f
    "00010000", -- 3083 - 0xc0b  :   16 - 0x10
    "00011111", -- 3084 - 0xc0c  :   31 - 0x1f
    "00010000", -- 3085 - 0xc0d  :   16 - 0x10
    "00010000", -- 3086 - 0xc0e  :   16 - 0x10
    "10010000", -- 3087 - 0xc0f  :  144 - 0x90
    "00111111", -- 3088 - 0xc10  :   63 - 0x3f -- Background 0x82
    "01111000", -- 3089 - 0xc11  :  120 - 0x78
    "11100111", -- 3090 - 0xc12  :  231 - 0xe7
    "11001111", -- 3091 - 0xc13  :  207 - 0xcf
    "01011000", -- 3092 - 0xc14  :   88 - 0x58
    "01011000", -- 3093 - 0xc15  :   88 - 0x58
    "01010000", -- 3094 - 0xc16  :   80 - 0x50
    "10010000", -- 3095 - 0xc17  :  144 - 0x90
    "10110000", -- 3096 - 0xc18  :  176 - 0xb0 -- Background 0x83
    "11111100", -- 3097 - 0xc19  :  252 - 0xfc
    "11100010", -- 3098 - 0xc1a  :  226 - 0xe2
    "11000001", -- 3099 - 0xc1b  :  193 - 0xc1
    "11000001", -- 3100 - 0xc1c  :  193 - 0xc1
    "10000011", -- 3101 - 0xc1d  :  131 - 0x83
    "10001111", -- 3102 - 0xc1e  :  143 - 0x8f
    "01111110", -- 3103 - 0xc1f  :  126 - 0x7e
    "11111110", -- 3104 - 0xc20  :  254 - 0xfe -- Background 0x84
    "00000011", -- 3105 - 0xc21  :    3 - 0x3
    "00001111", -- 3106 - 0xc22  :   15 - 0xf
    "10010001", -- 3107 - 0xc23  :  145 - 0x91
    "01110000", -- 3108 - 0xc24  :  112 - 0x70
    "01100000", -- 3109 - 0xc25  :   96 - 0x60
    "00100000", -- 3110 - 0xc26  :   32 - 0x20
    "00110001", -- 3111 - 0xc27  :   49 - 0x31
    "00111111", -- 3112 - 0xc28  :   63 - 0x3f -- Background 0x85
    "00111111", -- 3113 - 0xc29  :   63 - 0x3f
    "00011101", -- 3114 - 0xc2a  :   29 - 0x1d
    "00111001", -- 3115 - 0xc2b  :   57 - 0x39
    "01111011", -- 3116 - 0xc2c  :  123 - 0x7b
    "11110011", -- 3117 - 0xc2d  :  243 - 0xf3
    "10000110", -- 3118 - 0xc2e  :  134 - 0x86
    "11111110", -- 3119 - 0xc2f  :  254 - 0xfe
    "11111111", -- 3120 - 0xc30  :  255 - 0xff -- Background 0x86
    "11111111", -- 3121 - 0xc31  :  255 - 0xff
    "11111111", -- 3122 - 0xc32  :  255 - 0xff
    "11111111", -- 3123 - 0xc33  :  255 - 0xff
    "11111111", -- 3124 - 0xc34  :  255 - 0xff
    "10000000", -- 3125 - 0xc35  :  128 - 0x80
    "10000000", -- 3126 - 0xc36  :  128 - 0x80
    "11111111", -- 3127 - 0xc37  :  255 - 0xff
    "11111110", -- 3128 - 0xc38  :  254 - 0xfe -- Background 0x87
    "11111111", -- 3129 - 0xc39  :  255 - 0xff
    "11111111", -- 3130 - 0xc3a  :  255 - 0xff
    "11111111", -- 3131 - 0xc3b  :  255 - 0xff
    "11111111", -- 3132 - 0xc3c  :  255 - 0xff
    "00000011", -- 3133 - 0xc3d  :    3 - 0x3
    "00000011", -- 3134 - 0xc3e  :    3 - 0x3
    "11111111", -- 3135 - 0xc3f  :  255 - 0xff
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0x88
    "11111111", -- 3137 - 0xc41  :  255 - 0xff
    "11111111", -- 3138 - 0xc42  :  255 - 0xff
    "11111111", -- 3139 - 0xc43  :  255 - 0xff
    "11111111", -- 3140 - 0xc44  :  255 - 0xff
    "11111111", -- 3141 - 0xc45  :  255 - 0xff
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00111100", -- 3144 - 0xc48  :   60 - 0x3c -- Background 0x89
    "11111100", -- 3145 - 0xc49  :  252 - 0xfc
    "11111100", -- 3146 - 0xc4a  :  252 - 0xfc
    "11111100", -- 3147 - 0xc4b  :  252 - 0xfc
    "11111100", -- 3148 - 0xc4c  :  252 - 0xfc
    "11111100", -- 3149 - 0xc4d  :  252 - 0xfc
    "00000100", -- 3150 - 0xc4e  :    4 - 0x4
    "00000100", -- 3151 - 0xc4f  :    4 - 0x4
    "11111111", -- 3152 - 0xc50  :  255 - 0xff -- Background 0x8a
    "11111111", -- 3153 - 0xc51  :  255 - 0xff
    "11111111", -- 3154 - 0xc52  :  255 - 0xff
    "11111111", -- 3155 - 0xc53  :  255 - 0xff
    "10000000", -- 3156 - 0xc54  :  128 - 0x80
    "11111111", -- 3157 - 0xc55  :  255 - 0xff
    "11111111", -- 3158 - 0xc56  :  255 - 0xff
    "11111111", -- 3159 - 0xc57  :  255 - 0xff
    "11111111", -- 3160 - 0xc58  :  255 - 0xff -- Background 0x8b
    "11111111", -- 3161 - 0xc59  :  255 - 0xff
    "11111111", -- 3162 - 0xc5a  :  255 - 0xff
    "11111111", -- 3163 - 0xc5b  :  255 - 0xff
    "00000011", -- 3164 - 0xc5c  :    3 - 0x3
    "11111111", -- 3165 - 0xc5d  :  255 - 0xff
    "11111111", -- 3166 - 0xc5e  :  255 - 0xff
    "11111111", -- 3167 - 0xc5f  :  255 - 0xff
    "11111111", -- 3168 - 0xc60  :  255 - 0xff -- Background 0x8c
    "11111111", -- 3169 - 0xc61  :  255 - 0xff
    "11111111", -- 3170 - 0xc62  :  255 - 0xff
    "11111111", -- 3171 - 0xc63  :  255 - 0xff
    "11111111", -- 3172 - 0xc64  :  255 - 0xff
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "11111111", -- 3174 - 0xc66  :  255 - 0xff
    "11111111", -- 3175 - 0xc67  :  255 - 0xff
    "11111100", -- 3176 - 0xc68  :  252 - 0xfc -- Background 0x8d
    "11111100", -- 3177 - 0xc69  :  252 - 0xfc
    "11111110", -- 3178 - 0xc6a  :  254 - 0xfe
    "11111110", -- 3179 - 0xc6b  :  254 - 0xfe
    "11111110", -- 3180 - 0xc6c  :  254 - 0xfe
    "00000010", -- 3181 - 0xc6d  :    2 - 0x2
    "11111110", -- 3182 - 0xc6e  :  254 - 0xfe
    "11111110", -- 3183 - 0xc6f  :  254 - 0xfe
    "11111111", -- 3184 - 0xc70  :  255 - 0xff -- Background 0x8e
    "10000000", -- 3185 - 0xc71  :  128 - 0x80
    "10000000", -- 3186 - 0xc72  :  128 - 0x80
    "10000000", -- 3187 - 0xc73  :  128 - 0x80
    "10000000", -- 3188 - 0xc74  :  128 - 0x80
    "10000000", -- 3189 - 0xc75  :  128 - 0x80
    "10000000", -- 3190 - 0xc76  :  128 - 0x80
    "10000000", -- 3191 - 0xc77  :  128 - 0x80
    "11111111", -- 3192 - 0xc78  :  255 - 0xff -- Background 0x8f
    "00000011", -- 3193 - 0xc79  :    3 - 0x3
    "00000011", -- 3194 - 0xc7a  :    3 - 0x3
    "00000011", -- 3195 - 0xc7b  :    3 - 0x3
    "00000011", -- 3196 - 0xc7c  :    3 - 0x3
    "00000011", -- 3197 - 0xc7d  :    3 - 0x3
    "00000011", -- 3198 - 0xc7e  :    3 - 0x3
    "00000011", -- 3199 - 0xc7f  :    3 - 0x3
    "00000010", -- 3200 - 0xc80  :    2 - 0x2 -- Background 0x90
    "00000010", -- 3201 - 0xc81  :    2 - 0x2
    "00000010", -- 3202 - 0xc82  :    2 - 0x2
    "00000010", -- 3203 - 0xc83  :    2 - 0x2
    "00000010", -- 3204 - 0xc84  :    2 - 0x2
    "00000010", -- 3205 - 0xc85  :    2 - 0x2
    "00000100", -- 3206 - 0xc86  :    4 - 0x4
    "00000100", -- 3207 - 0xc87  :    4 - 0x4
    "10000000", -- 3208 - 0xc88  :  128 - 0x80 -- Background 0x91
    "10000000", -- 3209 - 0xc89  :  128 - 0x80
    "10101010", -- 3210 - 0xc8a  :  170 - 0xaa
    "11010101", -- 3211 - 0xc8b  :  213 - 0xd5
    "10101010", -- 3212 - 0xc8c  :  170 - 0xaa
    "11111111", -- 3213 - 0xc8d  :  255 - 0xff
    "11111111", -- 3214 - 0xc8e  :  255 - 0xff
    "11111111", -- 3215 - 0xc8f  :  255 - 0xff
    "00000011", -- 3216 - 0xc90  :    3 - 0x3 -- Background 0x92
    "00000011", -- 3217 - 0xc91  :    3 - 0x3
    "10101011", -- 3218 - 0xc92  :  171 - 0xab
    "01010111", -- 3219 - 0xc93  :   87 - 0x57
    "10101011", -- 3220 - 0xc94  :  171 - 0xab
    "11111111", -- 3221 - 0xc95  :  255 - 0xff
    "11111111", -- 3222 - 0xc96  :  255 - 0xff
    "11111110", -- 3223 - 0xc97  :  254 - 0xfe
    "00000000", -- 3224 - 0xc98  :    0 - 0x0 -- Background 0x93
    "01010101", -- 3225 - 0xc99  :   85 - 0x55
    "10101010", -- 3226 - 0xc9a  :  170 - 0xaa
    "01010101", -- 3227 - 0xc9b  :   85 - 0x55
    "11111111", -- 3228 - 0xc9c  :  255 - 0xff
    "11111111", -- 3229 - 0xc9d  :  255 - 0xff
    "11111111", -- 3230 - 0xc9e  :  255 - 0xff
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000100", -- 3232 - 0xca0  :    4 - 0x4 -- Background 0x94
    "01010100", -- 3233 - 0xca1  :   84 - 0x54
    "10101100", -- 3234 - 0xca2  :  172 - 0xac
    "01011100", -- 3235 - 0xca3  :   92 - 0x5c
    "11111100", -- 3236 - 0xca4  :  252 - 0xfc
    "11111100", -- 3237 - 0xca5  :  252 - 0xfc
    "11111100", -- 3238 - 0xca6  :  252 - 0xfc
    "00111100", -- 3239 - 0xca7  :   60 - 0x3c
    "00111111", -- 3240 - 0xca8  :   63 - 0x3f -- Background 0x95
    "00111111", -- 3241 - 0xca9  :   63 - 0x3f
    "00111111", -- 3242 - 0xcaa  :   63 - 0x3f
    "00111111", -- 3243 - 0xcab  :   63 - 0x3f
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "11111111", -- 3247 - 0xcaf  :  255 - 0xff
    "01111110", -- 3248 - 0xcb0  :  126 - 0x7e -- Background 0x96
    "01111100", -- 3249 - 0xcb1  :  124 - 0x7c
    "01111100", -- 3250 - 0xcb2  :  124 - 0x7c
    "01111000", -- 3251 - 0xcb3  :  120 - 0x78
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "11111111", -- 3255 - 0xcb7  :  255 - 0xff
    "00011111", -- 3256 - 0xcb8  :   31 - 0x1f -- Background 0x97
    "00001111", -- 3257 - 0xcb9  :   15 - 0xf
    "00001111", -- 3258 - 0xcba  :   15 - 0xf
    "00000111", -- 3259 - 0xcbb  :    7 - 0x7
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00000000", -- 3261 - 0xcbd  :    0 - 0x0
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "11111111", -- 3263 - 0xcbf  :  255 - 0xff
    "11111110", -- 3264 - 0xcc0  :  254 - 0xfe -- Background 0x98
    "11111100", -- 3265 - 0xcc1  :  252 - 0xfc
    "11111100", -- 3266 - 0xcc2  :  252 - 0xfc
    "11111000", -- 3267 - 0xcc3  :  248 - 0xf8
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "11111111", -- 3277 - 0xccd  :  255 - 0xff
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00011000", -- 3280 - 0xcd0  :   24 - 0x18 -- Background 0x9a
    "00011000", -- 3281 - 0xcd1  :   24 - 0x18
    "00011000", -- 3282 - 0xcd2  :   24 - 0x18
    "00011000", -- 3283 - 0xcd3  :   24 - 0x18
    "00011000", -- 3284 - 0xcd4  :   24 - 0x18
    "00011000", -- 3285 - 0xcd5  :   24 - 0x18
    "00011000", -- 3286 - 0xcd6  :   24 - 0x18
    "00011000", -- 3287 - 0xcd7  :   24 - 0x18
    "00000111", -- 3288 - 0xcd8  :    7 - 0x7 -- Background 0x9b
    "00011111", -- 3289 - 0xcd9  :   31 - 0x1f
    "00111111", -- 3290 - 0xcda  :   63 - 0x3f
    "11111111", -- 3291 - 0xcdb  :  255 - 0xff
    "01111111", -- 3292 - 0xcdc  :  127 - 0x7f
    "01111111", -- 3293 - 0xcdd  :  127 - 0x7f
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "11100001", -- 3296 - 0xce0  :  225 - 0xe1 -- Background 0x9c
    "11111001", -- 3297 - 0xce1  :  249 - 0xf9
    "11111101", -- 3298 - 0xce2  :  253 - 0xfd
    "11111111", -- 3299 - 0xce3  :  255 - 0xff
    "11111110", -- 3300 - 0xce4  :  254 - 0xfe
    "11111110", -- 3301 - 0xce5  :  254 - 0xfe
    "11111111", -- 3302 - 0xce6  :  255 - 0xff
    "11111111", -- 3303 - 0xce7  :  255 - 0xff
    "11110000", -- 3304 - 0xce8  :  240 - 0xf0 -- Background 0x9d
    "00010000", -- 3305 - 0xce9  :   16 - 0x10
    "00010000", -- 3306 - 0xcea  :   16 - 0x10
    "00010000", -- 3307 - 0xceb  :   16 - 0x10
    "00010000", -- 3308 - 0xcec  :   16 - 0x10
    "00010000", -- 3309 - 0xced  :   16 - 0x10
    "00010000", -- 3310 - 0xcee  :   16 - 0x10
    "11111111", -- 3311 - 0xcef  :  255 - 0xff
    "00011111", -- 3312 - 0xcf0  :   31 - 0x1f -- Background 0x9e
    "00010000", -- 3313 - 0xcf1  :   16 - 0x10
    "00010000", -- 3314 - 0xcf2  :   16 - 0x10
    "00010000", -- 3315 - 0xcf3  :   16 - 0x10
    "00010000", -- 3316 - 0xcf4  :   16 - 0x10
    "00010000", -- 3317 - 0xcf5  :   16 - 0x10
    "00010000", -- 3318 - 0xcf6  :   16 - 0x10
    "11111111", -- 3319 - 0xcf7  :  255 - 0xff
    "10010010", -- 3320 - 0xcf8  :  146 - 0x92 -- Background 0x9f
    "10010010", -- 3321 - 0xcf9  :  146 - 0x92
    "10010010", -- 3322 - 0xcfa  :  146 - 0x92
    "11111110", -- 3323 - 0xcfb  :  254 - 0xfe
    "11111110", -- 3324 - 0xcfc  :  254 - 0xfe
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00001010", -- 3328 - 0xd00  :   10 - 0xa -- Background 0xa0
    "00001010", -- 3329 - 0xd01  :   10 - 0xa
    "00111010", -- 3330 - 0xd02  :   58 - 0x3a
    "00001010", -- 3331 - 0xd03  :   10 - 0xa
    "11111011", -- 3332 - 0xd04  :  251 - 0xfb
    "00001011", -- 3333 - 0xd05  :   11 - 0xb
    "00001011", -- 3334 - 0xd06  :   11 - 0xb
    "00001011", -- 3335 - 0xd07  :   11 - 0xb
    "10010000", -- 3336 - 0xd08  :  144 - 0x90 -- Background 0xa1
    "10010000", -- 3337 - 0xd09  :  144 - 0x90
    "10011111", -- 3338 - 0xd0a  :  159 - 0x9f
    "10010000", -- 3339 - 0xd0b  :  144 - 0x90
    "10011111", -- 3340 - 0xd0c  :  159 - 0x9f
    "10010000", -- 3341 - 0xd0d  :  144 - 0x90
    "10010000", -- 3342 - 0xd0e  :  144 - 0x90
    "10010000", -- 3343 - 0xd0f  :  144 - 0x90
    "00000001", -- 3344 - 0xd10  :    1 - 0x1 -- Background 0xa2
    "00000001", -- 3345 - 0xd11  :    1 - 0x1
    "00000001", -- 3346 - 0xd12  :    1 - 0x1
    "00000001", -- 3347 - 0xd13  :    1 - 0x1
    "00000001", -- 3348 - 0xd14  :    1 - 0x1
    "00000001", -- 3349 - 0xd15  :    1 - 0x1
    "00000001", -- 3350 - 0xd16  :    1 - 0x1
    "00000001", -- 3351 - 0xd17  :    1 - 0x1
    "10000000", -- 3352 - 0xd18  :  128 - 0x80 -- Background 0xa3
    "10000000", -- 3353 - 0xd19  :  128 - 0x80
    "10000000", -- 3354 - 0xd1a  :  128 - 0x80
    "10000000", -- 3355 - 0xd1b  :  128 - 0x80
    "10000000", -- 3356 - 0xd1c  :  128 - 0x80
    "10000000", -- 3357 - 0xd1d  :  128 - 0x80
    "10000000", -- 3358 - 0xd1e  :  128 - 0x80
    "10000000", -- 3359 - 0xd1f  :  128 - 0x80
    "00001000", -- 3360 - 0xd20  :    8 - 0x8 -- Background 0xa4
    "10001000", -- 3361 - 0xd21  :  136 - 0x88
    "10010001", -- 3362 - 0xd22  :  145 - 0x91
    "11010001", -- 3363 - 0xd23  :  209 - 0xd1
    "01010011", -- 3364 - 0xd24  :   83 - 0x53
    "01010011", -- 3365 - 0xd25  :   83 - 0x53
    "01110011", -- 3366 - 0xd26  :  115 - 0x73
    "00111111", -- 3367 - 0xd27  :   63 - 0x3f
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000111", -- 3370 - 0xd2a  :    7 - 0x7
    "00001111", -- 3371 - 0xd2b  :   15 - 0xf
    "00001100", -- 3372 - 0xd2c  :   12 - 0xc
    "00011011", -- 3373 - 0xd2d  :   27 - 0x1b
    "00011011", -- 3374 - 0xd2e  :   27 - 0x1b
    "00011011", -- 3375 - 0xd2f  :   27 - 0x1b
    "00000000", -- 3376 - 0xd30  :    0 - 0x0 -- Background 0xa6
    "00000000", -- 3377 - 0xd31  :    0 - 0x0
    "11100000", -- 3378 - 0xd32  :  224 - 0xe0
    "11110000", -- 3379 - 0xd33  :  240 - 0xf0
    "11110000", -- 3380 - 0xd34  :  240 - 0xf0
    "11111000", -- 3381 - 0xd35  :  248 - 0xf8
    "11111000", -- 3382 - 0xd36  :  248 - 0xf8
    "11111000", -- 3383 - 0xd37  :  248 - 0xf8
    "00011011", -- 3384 - 0xd38  :   27 - 0x1b -- Background 0xa7
    "00011011", -- 3385 - 0xd39  :   27 - 0x1b
    "00011011", -- 3386 - 0xd3a  :   27 - 0x1b
    "00011011", -- 3387 - 0xd3b  :   27 - 0x1b
    "00011011", -- 3388 - 0xd3c  :   27 - 0x1b
    "00001111", -- 3389 - 0xd3d  :   15 - 0xf
    "00001111", -- 3390 - 0xd3e  :   15 - 0xf
    "00000111", -- 3391 - 0xd3f  :    7 - 0x7
    "11111000", -- 3392 - 0xd40  :  248 - 0xf8 -- Background 0xa8
    "11111000", -- 3393 - 0xd41  :  248 - 0xf8
    "11111000", -- 3394 - 0xd42  :  248 - 0xf8
    "11111000", -- 3395 - 0xd43  :  248 - 0xf8
    "11111000", -- 3396 - 0xd44  :  248 - 0xf8
    "11110000", -- 3397 - 0xd45  :  240 - 0xf0
    "11110000", -- 3398 - 0xd46  :  240 - 0xf0
    "11100000", -- 3399 - 0xd47  :  224 - 0xe0
    "11110001", -- 3400 - 0xd48  :  241 - 0xf1 -- Background 0xa9
    "00010001", -- 3401 - 0xd49  :   17 - 0x11
    "00010001", -- 3402 - 0xd4a  :   17 - 0x11
    "00011111", -- 3403 - 0xd4b  :   31 - 0x1f
    "00010000", -- 3404 - 0xd4c  :   16 - 0x10
    "00010000", -- 3405 - 0xd4d  :   16 - 0x10
    "00010000", -- 3406 - 0xd4e  :   16 - 0x10
    "11111111", -- 3407 - 0xd4f  :  255 - 0xff
    "00011111", -- 3408 - 0xd50  :   31 - 0x1f -- Background 0xaa
    "00010000", -- 3409 - 0xd51  :   16 - 0x10
    "00010000", -- 3410 - 0xd52  :   16 - 0x10
    "11110000", -- 3411 - 0xd53  :  240 - 0xf0
    "00010000", -- 3412 - 0xd54  :   16 - 0x10
    "00010000", -- 3413 - 0xd55  :   16 - 0x10
    "00010000", -- 3414 - 0xd56  :   16 - 0x10
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "01111111", -- 3416 - 0xd58  :  127 - 0x7f -- Background 0xab
    "10111111", -- 3417 - 0xd59  :  191 - 0xbf
    "11011111", -- 3418 - 0xd5a  :  223 - 0xdf
    "11101111", -- 3419 - 0xd5b  :  239 - 0xef
    "11110000", -- 3420 - 0xd5c  :  240 - 0xf0
    "11110000", -- 3421 - 0xd5d  :  240 - 0xf0
    "11110000", -- 3422 - 0xd5e  :  240 - 0xf0
    "11110000", -- 3423 - 0xd5f  :  240 - 0xf0
    "11110000", -- 3424 - 0xd60  :  240 - 0xf0 -- Background 0xac
    "11110000", -- 3425 - 0xd61  :  240 - 0xf0
    "11110000", -- 3426 - 0xd62  :  240 - 0xf0
    "11110000", -- 3427 - 0xd63  :  240 - 0xf0
    "11111111", -- 3428 - 0xd64  :  255 - 0xff
    "11111111", -- 3429 - 0xd65  :  255 - 0xff
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "11111111", -- 3432 - 0xd68  :  255 - 0xff -- Background 0xad
    "11111111", -- 3433 - 0xd69  :  255 - 0xff
    "11111111", -- 3434 - 0xd6a  :  255 - 0xff
    "11111111", -- 3435 - 0xd6b  :  255 - 0xff
    "00001111", -- 3436 - 0xd6c  :   15 - 0xf
    "00001111", -- 3437 - 0xd6d  :   15 - 0xf
    "00001111", -- 3438 - 0xd6e  :   15 - 0xf
    "00001111", -- 3439 - 0xd6f  :   15 - 0xf
    "00001111", -- 3440 - 0xd70  :   15 - 0xf -- Background 0xae
    "00001111", -- 3441 - 0xd71  :   15 - 0xf
    "00001111", -- 3442 - 0xd72  :   15 - 0xf
    "00001111", -- 3443 - 0xd73  :   15 - 0xf
    "11110111", -- 3444 - 0xd74  :  247 - 0xf7
    "11111011", -- 3445 - 0xd75  :  251 - 0xfb
    "11111101", -- 3446 - 0xd76  :  253 - 0xfd
    "11111110", -- 3447 - 0xd77  :  254 - 0xfe
    "00000000", -- 3448 - 0xd78  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "00000000", -- 3451 - 0xd7b  :    0 - 0x0
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00011000", -- 3454 - 0xd7e  :   24 - 0x18
    "00011000", -- 3455 - 0xd7f  :   24 - 0x18
    "00011111", -- 3456 - 0xd80  :   31 - 0x1f -- Background 0xb0
    "00111111", -- 3457 - 0xd81  :   63 - 0x3f
    "01111111", -- 3458 - 0xd82  :  127 - 0x7f
    "01111111", -- 3459 - 0xd83  :  127 - 0x7f
    "01111111", -- 3460 - 0xd84  :  127 - 0x7f
    "11111111", -- 3461 - 0xd85  :  255 - 0xff
    "11111111", -- 3462 - 0xd86  :  255 - 0xff
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11111111", -- 3464 - 0xd88  :  255 - 0xff -- Background 0xb1
    "11111111", -- 3465 - 0xd89  :  255 - 0xff
    "11111111", -- 3466 - 0xd8a  :  255 - 0xff
    "01111111", -- 3467 - 0xd8b  :  127 - 0x7f
    "01111111", -- 3468 - 0xd8c  :  127 - 0x7f
    "01111111", -- 3469 - 0xd8d  :  127 - 0x7f
    "00111111", -- 3470 - 0xd8e  :   63 - 0x3f
    "00011110", -- 3471 - 0xd8f  :   30 - 0x1e
    "11111000", -- 3472 - 0xd90  :  248 - 0xf8 -- Background 0xb2
    "11111100", -- 3473 - 0xd91  :  252 - 0xfc
    "11111110", -- 3474 - 0xd92  :  254 - 0xfe
    "11111110", -- 3475 - 0xd93  :  254 - 0xfe
    "11111110", -- 3476 - 0xd94  :  254 - 0xfe
    "11111111", -- 3477 - 0xd95  :  255 - 0xff
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111111", -- 3479 - 0xd97  :  255 - 0xff
    "11111111", -- 3480 - 0xd98  :  255 - 0xff -- Background 0xb3
    "11111111", -- 3481 - 0xd99  :  255 - 0xff
    "11111111", -- 3482 - 0xd9a  :  255 - 0xff
    "11111110", -- 3483 - 0xd9b  :  254 - 0xfe
    "11111110", -- 3484 - 0xd9c  :  254 - 0xfe
    "11111110", -- 3485 - 0xd9d  :  254 - 0xfe
    "11111100", -- 3486 - 0xd9e  :  252 - 0xfc
    "01111000", -- 3487 - 0xd9f  :  120 - 0x78
    "01111111", -- 3488 - 0xda0  :  127 - 0x7f -- Background 0xb4
    "10000000", -- 3489 - 0xda1  :  128 - 0x80
    "10000000", -- 3490 - 0xda2  :  128 - 0x80
    "10000000", -- 3491 - 0xda3  :  128 - 0x80
    "10000000", -- 3492 - 0xda4  :  128 - 0x80
    "10000000", -- 3493 - 0xda5  :  128 - 0x80
    "10000000", -- 3494 - 0xda6  :  128 - 0x80
    "10000000", -- 3495 - 0xda7  :  128 - 0x80
    "11011110", -- 3496 - 0xda8  :  222 - 0xde -- Background 0xb5
    "01100001", -- 3497 - 0xda9  :   97 - 0x61
    "01100001", -- 3498 - 0xdaa  :   97 - 0x61
    "01100001", -- 3499 - 0xdab  :   97 - 0x61
    "01110001", -- 3500 - 0xdac  :  113 - 0x71
    "01011110", -- 3501 - 0xdad  :   94 - 0x5e
    "01111111", -- 3502 - 0xdae  :  127 - 0x7f
    "01100001", -- 3503 - 0xdaf  :   97 - 0x61
    "10000000", -- 3504 - 0xdb0  :  128 - 0x80 -- Background 0xb6
    "10000000", -- 3505 - 0xdb1  :  128 - 0x80
    "11000000", -- 3506 - 0xdb2  :  192 - 0xc0
    "11110000", -- 3507 - 0xdb3  :  240 - 0xf0
    "10111111", -- 3508 - 0xdb4  :  191 - 0xbf
    "10001111", -- 3509 - 0xdb5  :  143 - 0x8f
    "10000001", -- 3510 - 0xdb6  :  129 - 0x81
    "01111110", -- 3511 - 0xdb7  :  126 - 0x7e
    "01100001", -- 3512 - 0xdb8  :   97 - 0x61 -- Background 0xb7
    "01100001", -- 3513 - 0xdb9  :   97 - 0x61
    "11000001", -- 3514 - 0xdba  :  193 - 0xc1
    "11000001", -- 3515 - 0xdbb  :  193 - 0xc1
    "10000001", -- 3516 - 0xdbc  :  129 - 0x81
    "10000001", -- 3517 - 0xdbd  :  129 - 0x81
    "10000011", -- 3518 - 0xdbe  :  131 - 0x83
    "11111110", -- 3519 - 0xdbf  :  254 - 0xfe
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xb8
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000011", -- 3522 - 0xdc2  :    3 - 0x3
    "00001111", -- 3523 - 0xdc3  :   15 - 0xf
    "00011111", -- 3524 - 0xdc4  :   31 - 0x1f
    "00111111", -- 3525 - 0xdc5  :   63 - 0x3f
    "01111111", -- 3526 - 0xdc6  :  127 - 0x7f
    "01111111", -- 3527 - 0xdc7  :  127 - 0x7f
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0 -- Background 0xb9
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "11000000", -- 3530 - 0xdca  :  192 - 0xc0
    "11110000", -- 3531 - 0xdcb  :  240 - 0xf0
    "11111000", -- 3532 - 0xdcc  :  248 - 0xf8
    "11111100", -- 3533 - 0xdcd  :  252 - 0xfc
    "11111110", -- 3534 - 0xdce  :  254 - 0xfe
    "11111110", -- 3535 - 0xdcf  :  254 - 0xfe
    "11111111", -- 3536 - 0xdd0  :  255 - 0xff -- Background 0xba
    "11111111", -- 3537 - 0xdd1  :  255 - 0xff
    "11111111", -- 3538 - 0xdd2  :  255 - 0xff
    "11111111", -- 3539 - 0xdd3  :  255 - 0xff
    "11111111", -- 3540 - 0xdd4  :  255 - 0xff
    "11111111", -- 3541 - 0xdd5  :  255 - 0xff
    "11111111", -- 3542 - 0xdd6  :  255 - 0xff
    "11111111", -- 3543 - 0xdd7  :  255 - 0xff
    "11111111", -- 3544 - 0xdd8  :  255 - 0xff -- Background 0xbb
    "11111111", -- 3545 - 0xdd9  :  255 - 0xff
    "11111111", -- 3546 - 0xdda  :  255 - 0xff
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "11111111", -- 3548 - 0xddc  :  255 - 0xff
    "11111111", -- 3549 - 0xddd  :  255 - 0xff
    "11111111", -- 3550 - 0xdde  :  255 - 0xff
    "11111111", -- 3551 - 0xddf  :  255 - 0xff
    "01111111", -- 3552 - 0xde0  :  127 - 0x7f -- Background 0xbc
    "01111111", -- 3553 - 0xde1  :  127 - 0x7f
    "01111111", -- 3554 - 0xde2  :  127 - 0x7f
    "00111111", -- 3555 - 0xde3  :   63 - 0x3f
    "00111111", -- 3556 - 0xde4  :   63 - 0x3f
    "00011111", -- 3557 - 0xde5  :   31 - 0x1f
    "00001111", -- 3558 - 0xde6  :   15 - 0xf
    "00000111", -- 3559 - 0xde7  :    7 - 0x7
    "11111110", -- 3560 - 0xde8  :  254 - 0xfe -- Background 0xbd
    "11111110", -- 3561 - 0xde9  :  254 - 0xfe
    "11111110", -- 3562 - 0xdea  :  254 - 0xfe
    "11111100", -- 3563 - 0xdeb  :  252 - 0xfc
    "11111100", -- 3564 - 0xdec  :  252 - 0xfc
    "11111000", -- 3565 - 0xded  :  248 - 0xf8
    "11110000", -- 3566 - 0xdee  :  240 - 0xf0
    "11110000", -- 3567 - 0xdef  :  240 - 0xf0
    "00001111", -- 3568 - 0xdf0  :   15 - 0xf -- Background 0xbe
    "00001111", -- 3569 - 0xdf1  :   15 - 0xf
    "00001111", -- 3570 - 0xdf2  :   15 - 0xf
    "00001111", -- 3571 - 0xdf3  :   15 - 0xf
    "00001111", -- 3572 - 0xdf4  :   15 - 0xf
    "00001111", -- 3573 - 0xdf5  :   15 - 0xf
    "00000111", -- 3574 - 0xdf6  :    7 - 0x7
    "00001111", -- 3575 - 0xdf7  :   15 - 0xf
    "11110000", -- 3576 - 0xdf8  :  240 - 0xf0 -- Background 0xbf
    "11110000", -- 3577 - 0xdf9  :  240 - 0xf0
    "11110000", -- 3578 - 0xdfa  :  240 - 0xf0
    "11110000", -- 3579 - 0xdfb  :  240 - 0xf0
    "11110000", -- 3580 - 0xdfc  :  240 - 0xf0
    "11110000", -- 3581 - 0xdfd  :  240 - 0xf0
    "11100000", -- 3582 - 0xdfe  :  224 - 0xe0
    "11110000", -- 3583 - 0xdff  :  240 - 0xf0
    "10000001", -- 3584 - 0xe00  :  129 - 0x81 -- Background 0xc0
    "11000001", -- 3585 - 0xe01  :  193 - 0xc1
    "10100011", -- 3586 - 0xe02  :  163 - 0xa3
    "10100011", -- 3587 - 0xe03  :  163 - 0xa3
    "10011101", -- 3588 - 0xe04  :  157 - 0x9d
    "10000001", -- 3589 - 0xe05  :  129 - 0x81
    "10000001", -- 3590 - 0xe06  :  129 - 0x81
    "10000001", -- 3591 - 0xe07  :  129 - 0x81
    "11100011", -- 3592 - 0xe08  :  227 - 0xe3 -- Background 0xc1
    "11110111", -- 3593 - 0xe09  :  247 - 0xf7
    "11000001", -- 3594 - 0xe0a  :  193 - 0xc1
    "11000001", -- 3595 - 0xe0b  :  193 - 0xc1
    "11000001", -- 3596 - 0xe0c  :  193 - 0xc1
    "11000001", -- 3597 - 0xe0d  :  193 - 0xc1
    "11110111", -- 3598 - 0xe0e  :  247 - 0xf7
    "11100011", -- 3599 - 0xe0f  :  227 - 0xe3
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000111", -- 3602 - 0xe12  :    7 - 0x7
    "00001111", -- 3603 - 0xe13  :   15 - 0xf
    "00001100", -- 3604 - 0xe14  :   12 - 0xc
    "00011011", -- 3605 - 0xe15  :   27 - 0x1b
    "00011011", -- 3606 - 0xe16  :   27 - 0x1b
    "00011011", -- 3607 - 0xe17  :   27 - 0x1b
    "00000000", -- 3608 - 0xe18  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "11100000", -- 3610 - 0xe1a  :  224 - 0xe0
    "11110000", -- 3611 - 0xe1b  :  240 - 0xf0
    "11110000", -- 3612 - 0xe1c  :  240 - 0xf0
    "11111000", -- 3613 - 0xe1d  :  248 - 0xf8
    "11111000", -- 3614 - 0xe1e  :  248 - 0xf8
    "11111000", -- 3615 - 0xe1f  :  248 - 0xf8
    "00011011", -- 3616 - 0xe20  :   27 - 0x1b -- Background 0xc4
    "00011011", -- 3617 - 0xe21  :   27 - 0x1b
    "00011011", -- 3618 - 0xe22  :   27 - 0x1b
    "00011011", -- 3619 - 0xe23  :   27 - 0x1b
    "00011011", -- 3620 - 0xe24  :   27 - 0x1b
    "00001111", -- 3621 - 0xe25  :   15 - 0xf
    "00001111", -- 3622 - 0xe26  :   15 - 0xf
    "00000111", -- 3623 - 0xe27  :    7 - 0x7
    "11111000", -- 3624 - 0xe28  :  248 - 0xf8 -- Background 0xc5
    "11111000", -- 3625 - 0xe29  :  248 - 0xf8
    "11111000", -- 3626 - 0xe2a  :  248 - 0xf8
    "11111000", -- 3627 - 0xe2b  :  248 - 0xf8
    "11111000", -- 3628 - 0xe2c  :  248 - 0xf8
    "11110000", -- 3629 - 0xe2d  :  240 - 0xf0
    "11110000", -- 3630 - 0xe2e  :  240 - 0xf0
    "11100000", -- 3631 - 0xe2f  :  224 - 0xe0
    "11100000", -- 3632 - 0xe30  :  224 - 0xe0 -- Background 0xc6
    "11111111", -- 3633 - 0xe31  :  255 - 0xff
    "11111111", -- 3634 - 0xe32  :  255 - 0xff
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "11111111", -- 3636 - 0xe34  :  255 - 0xff
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "00000111", -- 3640 - 0xe38  :    7 - 0x7 -- Background 0xc7
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "11111111", -- 3642 - 0xe3a  :  255 - 0xff
    "11111111", -- 3643 - 0xe3b  :  255 - 0xff
    "11111111", -- 3644 - 0xe3c  :  255 - 0xff
    "11111111", -- 3645 - 0xe3d  :  255 - 0xff
    "11111111", -- 3646 - 0xe3e  :  255 - 0xff
    "11111111", -- 3647 - 0xe3f  :  255 - 0xff
    "11111111", -- 3648 - 0xe40  :  255 - 0xff -- Background 0xc8
    "11111111", -- 3649 - 0xe41  :  255 - 0xff
    "11111111", -- 3650 - 0xe42  :  255 - 0xff
    "11111111", -- 3651 - 0xe43  :  255 - 0xff
    "11111111", -- 3652 - 0xe44  :  255 - 0xff
    "11111110", -- 3653 - 0xe45  :  254 - 0xfe
    "11111111", -- 3654 - 0xe46  :  255 - 0xff
    "11101111", -- 3655 - 0xe47  :  239 - 0xef
    "11111111", -- 3656 - 0xe48  :  255 - 0xff -- Background 0xc9
    "11011111", -- 3657 - 0xe49  :  223 - 0xdf
    "11101111", -- 3658 - 0xe4a  :  239 - 0xef
    "10101111", -- 3659 - 0xe4b  :  175 - 0xaf
    "10101111", -- 3660 - 0xe4c  :  175 - 0xaf
    "01101111", -- 3661 - 0xe4d  :  111 - 0x6f
    "11101111", -- 3662 - 0xe4e  :  239 - 0xef
    "11100111", -- 3663 - 0xe4f  :  231 - 0xe7
    "00011111", -- 3664 - 0xe50  :   31 - 0x1f -- Background 0xca
    "00011111", -- 3665 - 0xe51  :   31 - 0x1f
    "00111111", -- 3666 - 0xe52  :   63 - 0x3f
    "00111111", -- 3667 - 0xe53  :   63 - 0x3f
    "01110000", -- 3668 - 0xe54  :  112 - 0x70
    "01100011", -- 3669 - 0xe55  :   99 - 0x63
    "11100111", -- 3670 - 0xe56  :  231 - 0xe7
    "11100101", -- 3671 - 0xe57  :  229 - 0xe5
    "11110000", -- 3672 - 0xe58  :  240 - 0xf0 -- Background 0xcb
    "11110000", -- 3673 - 0xe59  :  240 - 0xf0
    "11111000", -- 3674 - 0xe5a  :  248 - 0xf8
    "11111000", -- 3675 - 0xe5b  :  248 - 0xf8
    "00001100", -- 3676 - 0xe5c  :   12 - 0xc
    "11000100", -- 3677 - 0xe5d  :  196 - 0xc4
    "11100100", -- 3678 - 0xe5e  :  228 - 0xe4
    "10100110", -- 3679 - 0xe5f  :  166 - 0xa6
    "11101001", -- 3680 - 0xe60  :  233 - 0xe9 -- Background 0xcc
    "11101001", -- 3681 - 0xe61  :  233 - 0xe9
    "11101001", -- 3682 - 0xe62  :  233 - 0xe9
    "11101111", -- 3683 - 0xe63  :  239 - 0xef
    "11100010", -- 3684 - 0xe64  :  226 - 0xe2
    "11100011", -- 3685 - 0xe65  :  227 - 0xe3
    "11110000", -- 3686 - 0xe66  :  240 - 0xf0
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "10010110", -- 3688 - 0xe68  :  150 - 0x96 -- Background 0xcd
    "10010110", -- 3689 - 0xe69  :  150 - 0x96
    "10010110", -- 3690 - 0xe6a  :  150 - 0x96
    "11110110", -- 3691 - 0xe6b  :  246 - 0xf6
    "01000110", -- 3692 - 0xe6c  :   70 - 0x46
    "11000110", -- 3693 - 0xe6d  :  198 - 0xc6
    "00001110", -- 3694 - 0xe6e  :   14 - 0xe
    "11111110", -- 3695 - 0xe6f  :  254 - 0xfe
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "01111110", -- 3702 - 0xe76  :  126 - 0x7e
    "00111100", -- 3703 - 0xe77  :   60 - 0x3c
    "00111100", -- 3704 - 0xe78  :   60 - 0x3c -- Background 0xcf
    "01000010", -- 3705 - 0xe79  :   66 - 0x42
    "10011001", -- 3706 - 0xe7a  :  153 - 0x99
    "10100001", -- 3707 - 0xe7b  :  161 - 0xa1
    "10100001", -- 3708 - 0xe7c  :  161 - 0xa1
    "10011001", -- 3709 - 0xe7d  :  153 - 0x99
    "01000010", -- 3710 - 0xe7e  :   66 - 0x42
    "00111100", -- 3711 - 0xe7f  :   60 - 0x3c
    "00001111", -- 3712 - 0xe80  :   15 - 0xf -- Background 0xd0
    "00011111", -- 3713 - 0xe81  :   31 - 0x1f
    "00011111", -- 3714 - 0xe82  :   31 - 0x1f
    "00111111", -- 3715 - 0xe83  :   63 - 0x3f
    "00111111", -- 3716 - 0xe84  :   63 - 0x3f
    "01111111", -- 3717 - 0xe85  :  127 - 0x7f
    "01111111", -- 3718 - 0xe86  :  127 - 0x7f
    "01111111", -- 3719 - 0xe87  :  127 - 0x7f
    "11110000", -- 3720 - 0xe88  :  240 - 0xf0 -- Background 0xd1
    "11111000", -- 3721 - 0xe89  :  248 - 0xf8
    "11111000", -- 3722 - 0xe8a  :  248 - 0xf8
    "11111100", -- 3723 - 0xe8b  :  252 - 0xfc
    "11111100", -- 3724 - 0xe8c  :  252 - 0xfc
    "11111110", -- 3725 - 0xe8d  :  254 - 0xfe
    "11111110", -- 3726 - 0xe8e  :  254 - 0xfe
    "11111110", -- 3727 - 0xe8f  :  254 - 0xfe
    "01111111", -- 3728 - 0xe90  :  127 - 0x7f -- Background 0xd2
    "01111111", -- 3729 - 0xe91  :  127 - 0x7f
    "00111111", -- 3730 - 0xe92  :   63 - 0x3f
    "00111111", -- 3731 - 0xe93  :   63 - 0x3f
    "00111111", -- 3732 - 0xe94  :   63 - 0x3f
    "00111111", -- 3733 - 0xe95  :   63 - 0x3f
    "00011111", -- 3734 - 0xe96  :   31 - 0x1f
    "00011111", -- 3735 - 0xe97  :   31 - 0x1f
    "11111110", -- 3736 - 0xe98  :  254 - 0xfe -- Background 0xd3
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111100", -- 3740 - 0xe9c  :  252 - 0xfc
    "11111100", -- 3741 - 0xe9d  :  252 - 0xfc
    "11111110", -- 3742 - 0xe9e  :  254 - 0xfe
    "11111110", -- 3743 - 0xe9f  :  254 - 0xfe
    "01111111", -- 3744 - 0xea0  :  127 - 0x7f -- Background 0xd4
    "01111111", -- 3745 - 0xea1  :  127 - 0x7f
    "01111111", -- 3746 - 0xea2  :  127 - 0x7f
    "00111111", -- 3747 - 0xea3  :   63 - 0x3f
    "00111111", -- 3748 - 0xea4  :   63 - 0x3f
    "00111111", -- 3749 - 0xea5  :   63 - 0x3f
    "00111111", -- 3750 - 0xea6  :   63 - 0x3f
    "00011111", -- 3751 - 0xea7  :   31 - 0x1f
    "11111110", -- 3752 - 0xea8  :  254 - 0xfe -- Background 0xd5
    "11111110", -- 3753 - 0xea9  :  254 - 0xfe
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111110", -- 3759 - 0xeaf  :  254 - 0xfe
    "00011111", -- 3760 - 0xeb0  :   31 - 0x1f -- Background 0xd6
    "00001111", -- 3761 - 0xeb1  :   15 - 0xf
    "00001111", -- 3762 - 0xeb2  :   15 - 0xf
    "00000111", -- 3763 - 0xeb3  :    7 - 0x7
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "11111110", -- 3768 - 0xeb8  :  254 - 0xfe -- Background 0xd7
    "11111100", -- 3769 - 0xeb9  :  252 - 0xfc
    "11111100", -- 3770 - 0xeba  :  252 - 0xfc
    "11111000", -- 3771 - 0xebb  :  248 - 0xf8
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "01111110", -- 3776 - 0xec0  :  126 - 0x7e -- Background 0xd8
    "01111110", -- 3777 - 0xec1  :  126 - 0x7e
    "01111110", -- 3778 - 0xec2  :  126 - 0x7e
    "01111110", -- 3779 - 0xec3  :  126 - 0x7e
    "01111111", -- 3780 - 0xec4  :  127 - 0x7f
    "01111111", -- 3781 - 0xec5  :  127 - 0x7f
    "01111111", -- 3782 - 0xec6  :  127 - 0x7f
    "01111111", -- 3783 - 0xec7  :  127 - 0x7f
    "11111111", -- 3784 - 0xec8  :  255 - 0xff -- Background 0xd9
    "11111111", -- 3785 - 0xec9  :  255 - 0xff
    "11111111", -- 3786 - 0xeca  :  255 - 0xff
    "11111111", -- 3787 - 0xecb  :  255 - 0xff
    "11111111", -- 3788 - 0xecc  :  255 - 0xff
    "11111111", -- 3789 - 0xecd  :  255 - 0xff
    "11111111", -- 3790 - 0xece  :  255 - 0xff
    "11111110", -- 3791 - 0xecf  :  254 - 0xfe
    "11111110", -- 3792 - 0xed0  :  254 - 0xfe -- Background 0xda
    "11111110", -- 3793 - 0xed1  :  254 - 0xfe
    "11111110", -- 3794 - 0xed2  :  254 - 0xfe
    "11111110", -- 3795 - 0xed3  :  254 - 0xfe
    "11111111", -- 3796 - 0xed4  :  255 - 0xff
    "11111111", -- 3797 - 0xed5  :  255 - 0xff
    "11111111", -- 3798 - 0xed6  :  255 - 0xff
    "11111111", -- 3799 - 0xed7  :  255 - 0xff
    "01111111", -- 3800 - 0xed8  :  127 - 0x7f -- Background 0xdb
    "01111111", -- 3801 - 0xed9  :  127 - 0x7f
    "01111111", -- 3802 - 0xeda  :  127 - 0x7f
    "01111111", -- 3803 - 0xedb  :  127 - 0x7f
    "01111111", -- 3804 - 0xedc  :  127 - 0x7f
    "01111111", -- 3805 - 0xedd  :  127 - 0x7f
    "01111111", -- 3806 - 0xede  :  127 - 0x7f
    "01111111", -- 3807 - 0xedf  :  127 - 0x7f
    "11111111", -- 3808 - 0xee0  :  255 - 0xff -- Background 0xdc
    "11111111", -- 3809 - 0xee1  :  255 - 0xff
    "11111111", -- 3810 - 0xee2  :  255 - 0xff
    "11111111", -- 3811 - 0xee3  :  255 - 0xff
    "11111100", -- 3812 - 0xee4  :  252 - 0xfc
    "11111110", -- 3813 - 0xee5  :  254 - 0xfe
    "11111110", -- 3814 - 0xee6  :  254 - 0xfe
    "01111110", -- 3815 - 0xee7  :  126 - 0x7e
    "11111111", -- 3816 - 0xee8  :  255 - 0xff -- Background 0xdd
    "11111111", -- 3817 - 0xee9  :  255 - 0xff
    "11111111", -- 3818 - 0xeea  :  255 - 0xff
    "11111111", -- 3819 - 0xeeb  :  255 - 0xff
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "01111111", -- 3824 - 0xef0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 3825 - 0xef1  :  127 - 0x7f
    "01111111", -- 3826 - 0xef2  :  127 - 0x7f
    "01111111", -- 3827 - 0xef3  :  127 - 0x7f
    "01111111", -- 3828 - 0xef4  :  127 - 0x7f
    "01111111", -- 3829 - 0xef5  :  127 - 0x7f
    "01111111", -- 3830 - 0xef6  :  127 - 0x7f
    "01111111", -- 3831 - 0xef7  :  127 - 0x7f
    "11111111", -- 3832 - 0xef8  :  255 - 0xff -- Background 0xdf
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "11111111", -- 3834 - 0xefa  :  255 - 0xff
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111111", -- 3836 - 0xefc  :  255 - 0xff
    "11111111", -- 3837 - 0xefd  :  255 - 0xff
    "11111111", -- 3838 - 0xefe  :  255 - 0xff
    "11111110", -- 3839 - 0xeff  :  254 - 0xfe
    "01111110", -- 3840 - 0xf00  :  126 - 0x7e -- Background 0xe0
    "01111110", -- 3841 - 0xf01  :  126 - 0x7e
    "01111111", -- 3842 - 0xf02  :  127 - 0x7f
    "01111111", -- 3843 - 0xf03  :  127 - 0x7f
    "01111111", -- 3844 - 0xf04  :  127 - 0x7f
    "01111111", -- 3845 - 0xf05  :  127 - 0x7f
    "01111111", -- 3846 - 0xf06  :  127 - 0x7f
    "01111111", -- 3847 - 0xf07  :  127 - 0x7f
    "00111111", -- 3848 - 0xf08  :   63 - 0x3f -- Background 0xe1
    "00111111", -- 3849 - 0xf09  :   63 - 0x3f
    "00111111", -- 3850 - 0xf0a  :   63 - 0x3f
    "00111111", -- 3851 - 0xf0b  :   63 - 0x3f
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "01111110", -- 3856 - 0xf10  :  126 - 0x7e -- Background 0xe2
    "01111100", -- 3857 - 0xf11  :  124 - 0x7c
    "01111100", -- 3858 - 0xf12  :  124 - 0x7c
    "01111000", -- 3859 - 0xf13  :  120 - 0x78
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "11111110", -- 3864 - 0xf18  :  254 - 0xfe -- Background 0xe3
    "11111110", -- 3865 - 0xf19  :  254 - 0xfe
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11111111", -- 3867 - 0xf1b  :  255 - 0xff
    "01111111", -- 3868 - 0xf1c  :  127 - 0x7f
    "01111111", -- 3869 - 0xf1d  :  127 - 0x7f
    "01111111", -- 3870 - 0xf1e  :  127 - 0x7f
    "01111111", -- 3871 - 0xf1f  :  127 - 0x7f
    "01111111", -- 3872 - 0xf20  :  127 - 0x7f -- Background 0xe4
    "01111111", -- 3873 - 0xf21  :  127 - 0x7f
    "00111111", -- 3874 - 0xf22  :   63 - 0x3f
    "00111111", -- 3875 - 0xf23  :   63 - 0x3f
    "00111111", -- 3876 - 0xf24  :   63 - 0x3f
    "00111111", -- 3877 - 0xf25  :   63 - 0x3f
    "00011111", -- 3878 - 0xf26  :   31 - 0x1f
    "00011111", -- 3879 - 0xf27  :   31 - 0x1f
    "00111111", -- 3880 - 0xf28  :   63 - 0x3f -- Background 0xe5
    "10111111", -- 3881 - 0xf29  :  191 - 0xbf
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11111111", -- 3883 - 0xf2b  :  255 - 0xff
    "11111100", -- 3884 - 0xf2c  :  252 - 0xfc
    "11111100", -- 3885 - 0xf2d  :  252 - 0xfc
    "11111110", -- 3886 - 0xf2e  :  254 - 0xfe
    "11111110", -- 3887 - 0xf2f  :  254 - 0xfe
    "01111111", -- 3888 - 0xf30  :  127 - 0x7f -- Background 0xe6
    "01111111", -- 3889 - 0xf31  :  127 - 0x7f
    "01111110", -- 3890 - 0xf32  :  126 - 0x7e
    "01111110", -- 3891 - 0xf33  :  126 - 0x7e
    "01111111", -- 3892 - 0xf34  :  127 - 0x7f
    "01111111", -- 3893 - 0xf35  :  127 - 0x7f
    "01111111", -- 3894 - 0xf36  :  127 - 0x7f
    "01111111", -- 3895 - 0xf37  :  127 - 0x7f
    "01111110", -- 3896 - 0xf38  :  126 - 0x7e -- Background 0xe7
    "01111110", -- 3897 - 0xf39  :  126 - 0x7e
    "01111110", -- 3898 - 0xf3a  :  126 - 0x7e
    "01111110", -- 3899 - 0xf3b  :  126 - 0x7e
    "01111111", -- 3900 - 0xf3c  :  127 - 0x7f
    "01111111", -- 3901 - 0xf3d  :  127 - 0x7f
    "01111111", -- 3902 - 0xf3e  :  127 - 0x7f
    "01111111", -- 3903 - 0xf3f  :  127 - 0x7f
    "10000001", -- 3904 - 0xf40  :  129 - 0x81 -- Background 0xe8
    "11000011", -- 3905 - 0xf41  :  195 - 0xc3
    "11000011", -- 3906 - 0xf42  :  195 - 0xc3
    "11100111", -- 3907 - 0xf43  :  231 - 0xe7
    "11100111", -- 3908 - 0xf44  :  231 - 0xe7
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "00001111", -- 3912 - 0xf48  :   15 - 0xf -- Background 0xe9
    "01000011", -- 3913 - 0xf49  :   67 - 0x43
    "01011011", -- 3914 - 0xf4a  :   91 - 0x5b
    "01010011", -- 3915 - 0xf4b  :   83 - 0x53
    "00110001", -- 3916 - 0xf4c  :   49 - 0x31
    "00011001", -- 3917 - 0xf4d  :   25 - 0x19
    "00001111", -- 3918 - 0xf4e  :   15 - 0xf
    "00000111", -- 3919 - 0xf4f  :    7 - 0x7
    "11000001", -- 3920 - 0xf50  :  193 - 0xc1 -- Background 0xea
    "11000011", -- 3921 - 0xf51  :  195 - 0xc3
    "11000110", -- 3922 - 0xf52  :  198 - 0xc6
    "10000100", -- 3923 - 0xf53  :  132 - 0x84
    "11111100", -- 3924 - 0xf54  :  252 - 0xfc
    "11111100", -- 3925 - 0xf55  :  252 - 0xfc
    "00001110", -- 3926 - 0xf56  :   14 - 0xe
    "00000010", -- 3927 - 0xf57  :    2 - 0x2
    "00010000", -- 3928 - 0xf58  :   16 - 0x10 -- Background 0xeb
    "00100000", -- 3929 - 0xf59  :   32 - 0x20
    "00100010", -- 3930 - 0xf5a  :   34 - 0x22
    "10111010", -- 3931 - 0xf5b  :  186 - 0xba
    "11100110", -- 3932 - 0xf5c  :  230 - 0xe6
    "11100001", -- 3933 - 0xf5d  :  225 - 0xe1
    "11000000", -- 3934 - 0xf5e  :  192 - 0xc0
    "11000000", -- 3935 - 0xf5f  :  192 - 0xc0
    "00100000", -- 3936 - 0xf60  :   32 - 0x20 -- Background 0xec
    "10100110", -- 3937 - 0xf61  :  166 - 0xa6
    "01010100", -- 3938 - 0xf62  :   84 - 0x54
    "00100110", -- 3939 - 0xf63  :   38 - 0x26
    "00100000", -- 3940 - 0xf64  :   32 - 0x20
    "11000110", -- 3941 - 0xf65  :  198 - 0xc6
    "01010100", -- 3942 - 0xf66  :   84 - 0x54
    "00100110", -- 3943 - 0xf67  :   38 - 0x26
    "00100000", -- 3944 - 0xf68  :   32 - 0x20 -- Background 0xed
    "10000101", -- 3945 - 0xf69  :  133 - 0x85
    "00000001", -- 3946 - 0xf6a  :    1 - 0x1
    "01000100", -- 3947 - 0xf6b  :   68 - 0x44
    "00100000", -- 3948 - 0xf6c  :   32 - 0x20
    "10000110", -- 3949 - 0xf6d  :  134 - 0x86
    "01010100", -- 3950 - 0xf6e  :   84 - 0x54
    "01001000", -- 3951 - 0xf6f  :   72 - 0x48
    "00100000", -- 3952 - 0xf70  :   32 - 0x20 -- Background 0xee
    "10111010", -- 3953 - 0xf71  :  186 - 0xba
    "11001001", -- 3954 - 0xf72  :  201 - 0xc9
    "01001010", -- 3955 - 0xf73  :   74 - 0x4a
    "00100000", -- 3956 - 0xf74  :   32 - 0x20
    "10100110", -- 3957 - 0xf75  :  166 - 0xa6
    "00001010", -- 3958 - 0xf76  :   10 - 0xa
    "11010000", -- 3959 - 0xf77  :  208 - 0xd0
    "11010001", -- 3960 - 0xf78  :  209 - 0xd1 -- Background 0xef
    "00100000", -- 3961 - 0xf79  :   32 - 0x20
    "11000110", -- 3962 - 0xf7a  :  198 - 0xc6
    "00001010", -- 3963 - 0xf7b  :   10 - 0xa
    "11010010", -- 3964 - 0xf7c  :  210 - 0xd2
    "11010011", -- 3965 - 0xf7d  :  211 - 0xd3
    "11011011", -- 3966 - 0xf7e  :  219 - 0xdb
    "11011011", -- 3967 - 0xf7f  :  219 - 0xdb
    "00001010", -- 3968 - 0xf80  :   10 - 0xa -- Background 0xf0
    "11010100", -- 3969 - 0xf81  :  212 - 0xd4
    "11010101", -- 3970 - 0xf82  :  213 - 0xd5
    "11010100", -- 3971 - 0xf83  :  212 - 0xd4
    "11011001", -- 3972 - 0xf84  :  217 - 0xd9
    "11011011", -- 3973 - 0xf85  :  219 - 0xdb
    "11100010", -- 3974 - 0xf86  :  226 - 0xe2
    "11010100", -- 3975 - 0xf87  :  212 - 0xd4
    "11010110", -- 3976 - 0xf88  :  214 - 0xd6 -- Background 0xf1
    "11010111", -- 3977 - 0xf89  :  215 - 0xd7
    "11100001", -- 3978 - 0xf8a  :  225 - 0xe1
    "00100110", -- 3979 - 0xf8b  :   38 - 0x26
    "11010110", -- 3980 - 0xf8c  :  214 - 0xd6
    "11011101", -- 3981 - 0xf8d  :  221 - 0xdd
    "11100001", -- 3982 - 0xf8e  :  225 - 0xe1
    "11100001", -- 3983 - 0xf8f  :  225 - 0xe1
    "11011110", -- 3984 - 0xf90  :  222 - 0xde -- Background 0xf2
    "11010001", -- 3985 - 0xf91  :  209 - 0xd1
    "11011000", -- 3986 - 0xf92  :  216 - 0xd8
    "11010000", -- 3987 - 0xf93  :  208 - 0xd0
    "11010001", -- 3988 - 0xf94  :  209 - 0xd1
    "00100110", -- 3989 - 0xf95  :   38 - 0x26
    "11011110", -- 3990 - 0xf96  :  222 - 0xde
    "11010001", -- 3991 - 0xf97  :  209 - 0xd1
    "01000110", -- 3992 - 0xf98  :   70 - 0x46 -- Background 0xf3
    "00010100", -- 3993 - 0xf99  :   20 - 0x14
    "11011011", -- 3994 - 0xf9a  :  219 - 0xdb
    "01000010", -- 3995 - 0xf9b  :   66 - 0x42
    "01000010", -- 3996 - 0xf9c  :   66 - 0x42
    "11011011", -- 3997 - 0xf9d  :  219 - 0xdb
    "01000010", -- 3998 - 0xf9e  :   66 - 0x42
    "11011011", -- 3999 - 0xf9f  :  219 - 0xdb
    "01000010", -- 4000 - 0xfa0  :   66 - 0x42 -- Background 0xf4
    "11011011", -- 4001 - 0xfa1  :  219 - 0xdb
    "01000010", -- 4002 - 0xfa2  :   66 - 0x42
    "11011011", -- 4003 - 0xfa3  :  219 - 0xdb
    "01000010", -- 4004 - 0xfa4  :   66 - 0x42
    "00100110", -- 4005 - 0xfa5  :   38 - 0x26
    "00100001", -- 4006 - 0xfa6  :   33 - 0x21
    "01100110", -- 4007 - 0xfa7  :  102 - 0x66
    "11011011", -- 4008 - 0xfa8  :  219 - 0xdb -- Background 0xf5
    "00100110", -- 4009 - 0xfa9  :   38 - 0x26
    "11011011", -- 4010 - 0xfaa  :  219 - 0xdb
    "11011111", -- 4011 - 0xfab  :  223 - 0xdf
    "11011011", -- 4012 - 0xfac  :  219 - 0xdb
    "11011111", -- 4013 - 0xfad  :  223 - 0xdf
    "11011011", -- 4014 - 0xfae  :  219 - 0xdb
    "11011011", -- 4015 - 0xfaf  :  219 - 0xdb
    "11011011", -- 4016 - 0xfb0  :  219 - 0xdb -- Background 0xf6
    "11011110", -- 4017 - 0xfb1  :  222 - 0xde
    "01000011", -- 4018 - 0xfb2  :   67 - 0x43
    "11011011", -- 4019 - 0xfb3  :  219 - 0xdb
    "11100000", -- 4020 - 0xfb4  :  224 - 0xe0
    "11011011", -- 4021 - 0xfb5  :  219 - 0xdb
    "11011011", -- 4022 - 0xfb6  :  219 - 0xdb
    "11011011", -- 4023 - 0xfb7  :  219 - 0xdb
    "11100011", -- 4024 - 0xfb8  :  227 - 0xe3 -- Background 0xf7
    "00100110", -- 4025 - 0xfb9  :   38 - 0x26
    "00100001", -- 4026 - 0xfba  :   33 - 0x21
    "10100110", -- 4027 - 0xfbb  :  166 - 0xa6
    "00010100", -- 4028 - 0xfbc  :   20 - 0x14
    "11011011", -- 4029 - 0xfbd  :  219 - 0xdb
    "11011011", -- 4030 - 0xfbe  :  219 - 0xdb
    "11011011", -- 4031 - 0xfbf  :  219 - 0xdb
    "11011011", -- 4032 - 0xfc0  :  219 - 0xdb -- Background 0xf8
    "11011001", -- 4033 - 0xfc1  :  217 - 0xd9
    "11011011", -- 4034 - 0xfc2  :  219 - 0xdb
    "11011011", -- 4035 - 0xfc3  :  219 - 0xdb
    "11010100", -- 4036 - 0xfc4  :  212 - 0xd4
    "11011001", -- 4037 - 0xfc5  :  217 - 0xd9
    "11010100", -- 4038 - 0xfc6  :  212 - 0xd4
    "11011001", -- 4039 - 0xfc7  :  217 - 0xd9
    "10010101", -- 4040 - 0xfc8  :  149 - 0x95 -- Background 0xf9
    "10010101", -- 4041 - 0xfc9  :  149 - 0x95
    "10010101", -- 4042 - 0xfca  :  149 - 0x95
    "10010101", -- 4043 - 0xfcb  :  149 - 0x95
    "10010101", -- 4044 - 0xfcc  :  149 - 0x95
    "10010111", -- 4045 - 0xfcd  :  151 - 0x97
    "10011000", -- 4046 - 0xfce  :  152 - 0x98
    "01111000", -- 4047 - 0xfcf  :  120 - 0x78
    "10010101", -- 4048 - 0xfd0  :  149 - 0x95 -- Background 0xfa
    "01111010", -- 4049 - 0xfd1  :  122 - 0x7a
    "00100001", -- 4050 - 0xfd2  :   33 - 0x21
    "11101101", -- 4051 - 0xfd3  :  237 - 0xed
    "00001110", -- 4052 - 0xfd4  :   14 - 0xe
    "11001111", -- 4053 - 0xfd5  :  207 - 0xcf
    "00000001", -- 4054 - 0xfd6  :    1 - 0x1
    "00001001", -- 4055 - 0xfd7  :    9 - 0x9
    "00010111", -- 4056 - 0xfd8  :   23 - 0x17 -- Background 0xfb
    "00001101", -- 4057 - 0xfd9  :   13 - 0xd
    "00011000", -- 4058 - 0xfda  :   24 - 0x18
    "00100010", -- 4059 - 0xfdb  :   34 - 0x22
    "01001011", -- 4060 - 0xfdc  :   75 - 0x4b
    "00001101", -- 4061 - 0xfdd  :   13 - 0xd
    "00000001", -- 4062 - 0xfde  :    1 - 0x1
    "00100100", -- 4063 - 0xfdf  :   36 - 0x24
    "00001010", -- 4064 - 0xfe0  :   10 - 0xa -- Background 0xfc
    "00010110", -- 4065 - 0xfe1  :   22 - 0x16
    "00001110", -- 4066 - 0xfe2  :   14 - 0xe
    "00100010", -- 4067 - 0xfe3  :   34 - 0x22
    "10001011", -- 4068 - 0xfe4  :  139 - 0x8b
    "00001101", -- 4069 - 0xfe5  :   13 - 0xd
    "00000010", -- 4070 - 0xfe6  :    2 - 0x2
    "00100100", -- 4071 - 0xfe7  :   36 - 0x24
    "00001010", -- 4072 - 0xfe8  :   10 - 0xa -- Background 0xfd
    "00010110", -- 4073 - 0xfe9  :   22 - 0x16
    "00001110", -- 4074 - 0xfea  :   14 - 0xe
    "00100010", -- 4075 - 0xfeb  :   34 - 0x22
    "11101100", -- 4076 - 0xfec  :  236 - 0xec
    "00000100", -- 4077 - 0xfed  :    4 - 0x4
    "00011101", -- 4078 - 0xfee  :   29 - 0x1d
    "00011000", -- 4079 - 0xfef  :   24 - 0x18
    "01010110", -- 4080 - 0xff0  :   86 - 0x56 -- Background 0xfe
    "01010101", -- 4081 - 0xff1  :   85 - 0x55
    "00100011", -- 4082 - 0xff2  :   35 - 0x23
    "11100010", -- 4083 - 0xff3  :  226 - 0xe2
    "00000100", -- 4084 - 0xff4  :    4 - 0x4
    "10011001", -- 4085 - 0xff5  :  153 - 0x99
    "10101010", -- 4086 - 0xff6  :  170 - 0xaa
    "10101010", -- 4087 - 0xff7  :  170 - 0xaa
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- Background 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
