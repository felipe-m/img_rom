//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables


//-  Original memory dump file name: pacman_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE_PACMAN_00
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      11'h0: dout <= 8'b00100000; //    0 :  32 - 0x20 -- line 0x0
      11'h1: dout <= 8'b00100000; //    1 :  32 - 0x20
      11'h2: dout <= 8'b00100000; //    2 :  32 - 0x20
      11'h3: dout <= 8'b00100000; //    3 :  32 - 0x20
      11'h4: dout <= 8'b00100000; //    4 :  32 - 0x20
      11'h5: dout <= 8'b00100000; //    5 :  32 - 0x20
      11'h6: dout <= 8'b00100000; //    6 :  32 - 0x20
      11'h7: dout <= 8'b00100000; //    7 :  32 - 0x20
      11'h8: dout <= 8'b00100000; //    8 :  32 - 0x20
      11'h9: dout <= 8'b00100000; //    9 :  32 - 0x20
      11'hA: dout <= 8'b00100000; //   10 :  32 - 0x20
      11'hB: dout <= 8'b00100000; //   11 :  32 - 0x20
      11'hC: dout <= 8'b00100000; //   12 :  32 - 0x20
      11'hD: dout <= 8'b00100000; //   13 :  32 - 0x20
      11'hE: dout <= 8'b00100000; //   14 :  32 - 0x20
      11'hF: dout <= 8'b00100000; //   15 :  32 - 0x20
      11'h10: dout <= 8'b00100000; //   16 :  32 - 0x20
      11'h11: dout <= 8'b00100000; //   17 :  32 - 0x20
      11'h12: dout <= 8'b00100000; //   18 :  32 - 0x20
      11'h13: dout <= 8'b00100000; //   19 :  32 - 0x20
      11'h14: dout <= 8'b00100000; //   20 :  32 - 0x20
      11'h15: dout <= 8'b00100000; //   21 :  32 - 0x20
      11'h16: dout <= 8'b00100000; //   22 :  32 - 0x20
      11'h17: dout <= 8'b00100000; //   23 :  32 - 0x20
      11'h18: dout <= 8'b00100000; //   24 :  32 - 0x20
      11'h19: dout <= 8'b00100000; //   25 :  32 - 0x20
      11'h1A: dout <= 8'b00100000; //   26 :  32 - 0x20
      11'h1B: dout <= 8'b00100000; //   27 :  32 - 0x20
      11'h1C: dout <= 8'b00100000; //   28 :  32 - 0x20
      11'h1D: dout <= 8'b00100000; //   29 :  32 - 0x20
      11'h1E: dout <= 8'b00100000; //   30 :  32 - 0x20
      11'h1F: dout <= 8'b00100000; //   31 :  32 - 0x20
      11'h20: dout <= 8'b00100000; //   32 :  32 - 0x20 -- line 0x1
      11'h21: dout <= 8'b00100000; //   33 :  32 - 0x20
      11'h22: dout <= 8'b00100000; //   34 :  32 - 0x20
      11'h23: dout <= 8'b00100000; //   35 :  32 - 0x20
      11'h24: dout <= 8'b00100000; //   36 :  32 - 0x20
      11'h25: dout <= 8'b00100000; //   37 :  32 - 0x20
      11'h26: dout <= 8'b00100000; //   38 :  32 - 0x20
      11'h27: dout <= 8'b00100000; //   39 :  32 - 0x20
      11'h28: dout <= 8'b00100000; //   40 :  32 - 0x20
      11'h29: dout <= 8'b00100000; //   41 :  32 - 0x20
      11'h2A: dout <= 8'b00100000; //   42 :  32 - 0x20
      11'h2B: dout <= 8'b00100000; //   43 :  32 - 0x20
      11'h2C: dout <= 8'b00100000; //   44 :  32 - 0x20
      11'h2D: dout <= 8'b00100000; //   45 :  32 - 0x20
      11'h2E: dout <= 8'b00100000; //   46 :  32 - 0x20
      11'h2F: dout <= 8'b00100000; //   47 :  32 - 0x20
      11'h30: dout <= 8'b00100000; //   48 :  32 - 0x20
      11'h31: dout <= 8'b00100000; //   49 :  32 - 0x20
      11'h32: dout <= 8'b00100000; //   50 :  32 - 0x20
      11'h33: dout <= 8'b00100000; //   51 :  32 - 0x20
      11'h34: dout <= 8'b00100000; //   52 :  32 - 0x20
      11'h35: dout <= 8'b00100000; //   53 :  32 - 0x20
      11'h36: dout <= 8'b00100000; //   54 :  32 - 0x20
      11'h37: dout <= 8'b00100000; //   55 :  32 - 0x20
      11'h38: dout <= 8'b00100000; //   56 :  32 - 0x20
      11'h39: dout <= 8'b00100000; //   57 :  32 - 0x20
      11'h3A: dout <= 8'b00100000; //   58 :  32 - 0x20
      11'h3B: dout <= 8'b00100000; //   59 :  32 - 0x20
      11'h3C: dout <= 8'b00100000; //   60 :  32 - 0x20
      11'h3D: dout <= 8'b00100000; //   61 :  32 - 0x20
      11'h3E: dout <= 8'b00100000; //   62 :  32 - 0x20
      11'h3F: dout <= 8'b00100000; //   63 :  32 - 0x20
      11'h40: dout <= 8'b00101101; //   64 :  45 - 0x2d -- line 0x2
      11'h41: dout <= 8'b00011111; //   65 :  31 - 0x1f
      11'h42: dout <= 8'b00010000; //   66 :  16 - 0x10
      11'h43: dout <= 8'b00010000; //   67 :  16 - 0x10
      11'h44: dout <= 8'b00010000; //   68 :  16 - 0x10
      11'h45: dout <= 8'b00010000; //   69 :  16 - 0x10
      11'h46: dout <= 8'b00010000; //   70 :  16 - 0x10
      11'h47: dout <= 8'b00010000; //   71 :  16 - 0x10
      11'h48: dout <= 8'b00010000; //   72 :  16 - 0x10
      11'h49: dout <= 8'b00010000; //   73 :  16 - 0x10
      11'h4A: dout <= 8'b00010000; //   74 :  16 - 0x10
      11'h4B: dout <= 8'b00010011; //   75 :  19 - 0x13
      11'h4C: dout <= 8'b00010000; //   76 :  16 - 0x10
      11'h4D: dout <= 8'b00010000; //   77 :  16 - 0x10
      11'h4E: dout <= 8'b00010000; //   78 :  16 - 0x10
      11'h4F: dout <= 8'b00010000; //   79 :  16 - 0x10
      11'h50: dout <= 8'b00010000; //   80 :  16 - 0x10
      11'h51: dout <= 8'b00010000; //   81 :  16 - 0x10
      11'h52: dout <= 8'b00010000; //   82 :  16 - 0x10
      11'h53: dout <= 8'b00010000; //   83 :  16 - 0x10
      11'h54: dout <= 8'b00010000; //   84 :  16 - 0x10
      11'h55: dout <= 8'b00011101; //   85 :  29 - 0x1d
      11'h56: dout <= 8'b00100000; //   86 :  32 - 0x20
      11'h57: dout <= 8'b00100000; //   87 :  32 - 0x20
      11'h58: dout <= 8'b00100000; //   88 :  32 - 0x20
      11'h59: dout <= 8'b00100000; //   89 :  32 - 0x20
      11'h5A: dout <= 8'b00100000; //   90 :  32 - 0x20
      11'h5B: dout <= 8'b00100000; //   91 :  32 - 0x20
      11'h5C: dout <= 8'b00100000; //   92 :  32 - 0x20
      11'h5D: dout <= 8'b00100000; //   93 :  32 - 0x20
      11'h5E: dout <= 8'b00100000; //   94 :  32 - 0x20
      11'h5F: dout <= 8'b00100000; //   95 :  32 - 0x20
      11'h60: dout <= 8'b00101101; //   96 :  45 - 0x2d -- line 0x3
      11'h61: dout <= 8'b00010001; //   97 :  17 - 0x11
      11'h62: dout <= 8'b00000011; //   98 :   3 - 0x3
      11'h63: dout <= 8'b00000011; //   99 :   3 - 0x3
      11'h64: dout <= 8'b00000011; //  100 :   3 - 0x3
      11'h65: dout <= 8'b00000011; //  101 :   3 - 0x3
      11'h66: dout <= 8'b00000011; //  102 :   3 - 0x3
      11'h67: dout <= 8'b00000011; //  103 :   3 - 0x3
      11'h68: dout <= 8'b00000011; //  104 :   3 - 0x3
      11'h69: dout <= 8'b00000011; //  105 :   3 - 0x3
      11'h6A: dout <= 8'b00000011; //  106 :   3 - 0x3
      11'h6B: dout <= 8'b00010001; //  107 :  17 - 0x11
      11'h6C: dout <= 8'b00000011; //  108 :   3 - 0x3
      11'h6D: dout <= 8'b00000011; //  109 :   3 - 0x3
      11'h6E: dout <= 8'b00000011; //  110 :   3 - 0x3
      11'h6F: dout <= 8'b00000011; //  111 :   3 - 0x3
      11'h70: dout <= 8'b00000011; //  112 :   3 - 0x3
      11'h71: dout <= 8'b00000011; //  113 :   3 - 0x3
      11'h72: dout <= 8'b00000011; //  114 :   3 - 0x3
      11'h73: dout <= 8'b00000011; //  115 :   3 - 0x3
      11'h74: dout <= 8'b00000011; //  116 :   3 - 0x3
      11'h75: dout <= 8'b00010001; //  117 :  17 - 0x11
      11'h76: dout <= 8'b10110100; //  118 : 180 - 0xb4
      11'h77: dout <= 8'b10110101; //  119 : 181 - 0xb5
      11'h78: dout <= 8'b10110110; //  120 : 182 - 0xb6
      11'h79: dout <= 8'b10110111; //  121 : 183 - 0xb7
      11'h7A: dout <= 8'b10111000; //  122 : 184 - 0xb8
      11'h7B: dout <= 8'b10111001; //  123 : 185 - 0xb9
      11'h7C: dout <= 8'b10111010; //  124 : 186 - 0xba
      11'h7D: dout <= 8'b10111011; //  125 : 187 - 0xbb
      11'h7E: dout <= 8'b00100000; //  126 :  32 - 0x20
      11'h7F: dout <= 8'b00100000; //  127 :  32 - 0x20
      11'h80: dout <= 8'b00101101; //  128 :  45 - 0x2d -- line 0x4
      11'h81: dout <= 8'b00010001; //  129 :  17 - 0x11
      11'h82: dout <= 8'b00000011; //  130 :   3 - 0x3
      11'h83: dout <= 8'b00011111; //  131 :  31 - 0x1f
      11'h84: dout <= 8'b00010000; //  132 :  16 - 0x10
      11'h85: dout <= 8'b00011101; //  133 :  29 - 0x1d
      11'h86: dout <= 8'b00000011; //  134 :   3 - 0x3
      11'h87: dout <= 8'b00011111; //  135 :  31 - 0x1f
      11'h88: dout <= 8'b00010000; //  136 :  16 - 0x10
      11'h89: dout <= 8'b00011101; //  137 :  29 - 0x1d
      11'h8A: dout <= 8'b00000011; //  138 :   3 - 0x3
      11'h8B: dout <= 8'b00010001; //  139 :  17 - 0x11
      11'h8C: dout <= 8'b00000011; //  140 :   3 - 0x3
      11'h8D: dout <= 8'b00011111; //  141 :  31 - 0x1f
      11'h8E: dout <= 8'b00010000; //  142 :  16 - 0x10
      11'h8F: dout <= 8'b00011101; //  143 :  29 - 0x1d
      11'h90: dout <= 8'b00000011; //  144 :   3 - 0x3
      11'h91: dout <= 8'b00011111; //  145 :  31 - 0x1f
      11'h92: dout <= 8'b00010000; //  146 :  16 - 0x10
      11'h93: dout <= 8'b00011101; //  147 :  29 - 0x1d
      11'h94: dout <= 8'b00000011; //  148 :   3 - 0x3
      11'h95: dout <= 8'b00010001; //  149 :  17 - 0x11
      11'h96: dout <= 8'b00100000; //  150 :  32 - 0x20
      11'h97: dout <= 8'b00100000; //  151 :  32 - 0x20
      11'h98: dout <= 8'b00100000; //  152 :  32 - 0x20
      11'h99: dout <= 8'b00100000; //  153 :  32 - 0x20
      11'h9A: dout <= 8'b00100000; //  154 :  32 - 0x20
      11'h9B: dout <= 8'b00100000; //  155 :  32 - 0x20
      11'h9C: dout <= 8'b00100000; //  156 :  32 - 0x20
      11'h9D: dout <= 8'b00100000; //  157 :  32 - 0x20
      11'h9E: dout <= 8'b00100000; //  158 :  32 - 0x20
      11'h9F: dout <= 8'b00100000; //  159 :  32 - 0x20
      11'hA0: dout <= 8'b00101101; //  160 :  45 - 0x2d -- line 0x5
      11'hA1: dout <= 8'b00010001; //  161 :  17 - 0x11
      11'hA2: dout <= 8'b00000001; //  162 :   1 - 0x1
      11'hA3: dout <= 8'b00010001; //  163 :  17 - 0x11
      11'hA4: dout <= 8'b00100000; //  164 :  32 - 0x20
      11'hA5: dout <= 8'b00010001; //  165 :  17 - 0x11
      11'hA6: dout <= 8'b00000011; //  166 :   3 - 0x3
      11'hA7: dout <= 8'b00010001; //  167 :  17 - 0x11
      11'hA8: dout <= 8'b00100000; //  168 :  32 - 0x20
      11'hA9: dout <= 8'b00010001; //  169 :  17 - 0x11
      11'hAA: dout <= 8'b00000011; //  170 :   3 - 0x3
      11'hAB: dout <= 8'b00010001; //  171 :  17 - 0x11
      11'hAC: dout <= 8'b00000011; //  172 :   3 - 0x3
      11'hAD: dout <= 8'b00010001; //  173 :  17 - 0x11
      11'hAE: dout <= 8'b00100000; //  174 :  32 - 0x20
      11'hAF: dout <= 8'b00010001; //  175 :  17 - 0x11
      11'hB0: dout <= 8'b00000011; //  176 :   3 - 0x3
      11'hB1: dout <= 8'b00010001; //  177 :  17 - 0x11
      11'hB2: dout <= 8'b00100000; //  178 :  32 - 0x20
      11'hB3: dout <= 8'b00010001; //  179 :  17 - 0x11
      11'hB4: dout <= 8'b00000001; //  180 :   1 - 0x1
      11'hB5: dout <= 8'b00010001; //  181 :  17 - 0x11
      11'hB6: dout <= 8'b00100000; //  182 :  32 - 0x20
      11'hB7: dout <= 8'b00100000; //  183 :  32 - 0x20
      11'hB8: dout <= 8'b00110001; //  184 :  49 - 0x31
      11'hB9: dout <= 8'b00110000; //  185 :  48 - 0x30
      11'hBA: dout <= 8'b00110000; //  186 :  48 - 0x30
      11'hBB: dout <= 8'b00110000; //  187 :  48 - 0x30
      11'hBC: dout <= 8'b00110000; //  188 :  48 - 0x30
      11'hBD: dout <= 8'b00100000; //  189 :  32 - 0x20
      11'hBE: dout <= 8'b00100000; //  190 :  32 - 0x20
      11'hBF: dout <= 8'b00100000; //  191 :  32 - 0x20
      11'hC0: dout <= 8'b00101101; //  192 :  45 - 0x2d -- line 0x6
      11'hC1: dout <= 8'b00010001; //  193 :  17 - 0x11
      11'hC2: dout <= 8'b00000011; //  194 :   3 - 0x3
      11'hC3: dout <= 8'b00011110; //  195 :  30 - 0x1e
      11'hC4: dout <= 8'b00010000; //  196 :  16 - 0x10
      11'hC5: dout <= 8'b00011100; //  197 :  28 - 0x1c
      11'hC6: dout <= 8'b00000011; //  198 :   3 - 0x3
      11'hC7: dout <= 8'b00011110; //  199 :  30 - 0x1e
      11'hC8: dout <= 8'b00010000; //  200 :  16 - 0x10
      11'hC9: dout <= 8'b00011100; //  201 :  28 - 0x1c
      11'hCA: dout <= 8'b00000011; //  202 :   3 - 0x3
      11'hCB: dout <= 8'b00011010; //  203 :  26 - 0x1a
      11'hCC: dout <= 8'b00000011; //  204 :   3 - 0x3
      11'hCD: dout <= 8'b00011110; //  205 :  30 - 0x1e
      11'hCE: dout <= 8'b00010000; //  206 :  16 - 0x10
      11'hCF: dout <= 8'b00011100; //  207 :  28 - 0x1c
      11'hD0: dout <= 8'b00000011; //  208 :   3 - 0x3
      11'hD1: dout <= 8'b00011110; //  209 :  30 - 0x1e
      11'hD2: dout <= 8'b00010000; //  210 :  16 - 0x10
      11'hD3: dout <= 8'b00011100; //  211 :  28 - 0x1c
      11'hD4: dout <= 8'b00000011; //  212 :   3 - 0x3
      11'hD5: dout <= 8'b00010001; //  213 :  17 - 0x11
      11'hD6: dout <= 8'b00100000; //  214 :  32 - 0x20
      11'hD7: dout <= 8'b00100000; //  215 :  32 - 0x20
      11'hD8: dout <= 8'b00100000; //  216 :  32 - 0x20
      11'hD9: dout <= 8'b00100000; //  217 :  32 - 0x20
      11'hDA: dout <= 8'b00100000; //  218 :  32 - 0x20
      11'hDB: dout <= 8'b00100000; //  219 :  32 - 0x20
      11'hDC: dout <= 8'b00100000; //  220 :  32 - 0x20
      11'hDD: dout <= 8'b00100000; //  221 :  32 - 0x20
      11'hDE: dout <= 8'b00100000; //  222 :  32 - 0x20
      11'hDF: dout <= 8'b00100000; //  223 :  32 - 0x20
      11'hE0: dout <= 8'b00101101; //  224 :  45 - 0x2d -- line 0x7
      11'hE1: dout <= 8'b00010001; //  225 :  17 - 0x11
      11'hE2: dout <= 8'b00000011; //  226 :   3 - 0x3
      11'hE3: dout <= 8'b00000011; //  227 :   3 - 0x3
      11'hE4: dout <= 8'b00000011; //  228 :   3 - 0x3
      11'hE5: dout <= 8'b00000011; //  229 :   3 - 0x3
      11'hE6: dout <= 8'b00000011; //  230 :   3 - 0x3
      11'hE7: dout <= 8'b00000011; //  231 :   3 - 0x3
      11'hE8: dout <= 8'b00000011; //  232 :   3 - 0x3
      11'hE9: dout <= 8'b00000011; //  233 :   3 - 0x3
      11'hEA: dout <= 8'b00000011; //  234 :   3 - 0x3
      11'hEB: dout <= 8'b00000011; //  235 :   3 - 0x3
      11'hEC: dout <= 8'b00000011; //  236 :   3 - 0x3
      11'hED: dout <= 8'b00000011; //  237 :   3 - 0x3
      11'hEE: dout <= 8'b00000011; //  238 :   3 - 0x3
      11'hEF: dout <= 8'b00000011; //  239 :   3 - 0x3
      11'hF0: dout <= 8'b00000011; //  240 :   3 - 0x3
      11'hF1: dout <= 8'b00000011; //  241 :   3 - 0x3
      11'hF2: dout <= 8'b00000011; //  242 :   3 - 0x3
      11'hF3: dout <= 8'b00000011; //  243 :   3 - 0x3
      11'hF4: dout <= 8'b00000011; //  244 :   3 - 0x3
      11'hF5: dout <= 8'b00010001; //  245 :  17 - 0x11
      11'hF6: dout <= 8'b00100000; //  246 :  32 - 0x20
      11'hF7: dout <= 8'b00100000; //  247 :  32 - 0x20
      11'hF8: dout <= 8'b00100000; //  248 :  32 - 0x20
      11'hF9: dout <= 8'b00100000; //  249 :  32 - 0x20
      11'hFA: dout <= 8'b00100000; //  250 :  32 - 0x20
      11'hFB: dout <= 8'b00100000; //  251 :  32 - 0x20
      11'hFC: dout <= 8'b00100000; //  252 :  32 - 0x20
      11'hFD: dout <= 8'b00100000; //  253 :  32 - 0x20
      11'hFE: dout <= 8'b00100000; //  254 :  32 - 0x20
      11'hFF: dout <= 8'b00100000; //  255 :  32 - 0x20
      11'h100: dout <= 8'b00101101; //  256 :  45 - 0x2d -- line 0x8
      11'h101: dout <= 8'b00010001; //  257 :  17 - 0x11
      11'h102: dout <= 8'b00000011; //  258 :   3 - 0x3
      11'h103: dout <= 8'b00011111; //  259 :  31 - 0x1f
      11'h104: dout <= 8'b00010000; //  260 :  16 - 0x10
      11'h105: dout <= 8'b00011101; //  261 :  29 - 0x1d
      11'h106: dout <= 8'b00000011; //  262 :   3 - 0x3
      11'h107: dout <= 8'b00011011; //  263 :  27 - 0x1b
      11'h108: dout <= 8'b00000011; //  264 :   3 - 0x3
      11'h109: dout <= 8'b00011111; //  265 :  31 - 0x1f
      11'h10A: dout <= 8'b00010000; //  266 :  16 - 0x10
      11'h10B: dout <= 8'b00010000; //  267 :  16 - 0x10
      11'h10C: dout <= 8'b00010000; //  268 :  16 - 0x10
      11'h10D: dout <= 8'b00011101; //  269 :  29 - 0x1d
      11'h10E: dout <= 8'b00000011; //  270 :   3 - 0x3
      11'h10F: dout <= 8'b00011011; //  271 :  27 - 0x1b
      11'h110: dout <= 8'b00000011; //  272 :   3 - 0x3
      11'h111: dout <= 8'b00011111; //  273 :  31 - 0x1f
      11'h112: dout <= 8'b00010000; //  274 :  16 - 0x10
      11'h113: dout <= 8'b00011101; //  275 :  29 - 0x1d
      11'h114: dout <= 8'b00000011; //  276 :   3 - 0x3
      11'h115: dout <= 8'b00010001; //  277 :  17 - 0x11
      11'h116: dout <= 8'b00100000; //  278 :  32 - 0x20
      11'h117: dout <= 8'b00100000; //  279 :  32 - 0x20
      11'h118: dout <= 8'b00100000; //  280 :  32 - 0x20
      11'h119: dout <= 8'b00100000; //  281 :  32 - 0x20
      11'h11A: dout <= 8'b00100000; //  282 :  32 - 0x20
      11'h11B: dout <= 8'b00100000; //  283 :  32 - 0x20
      11'h11C: dout <= 8'b00100000; //  284 :  32 - 0x20
      11'h11D: dout <= 8'b00100000; //  285 :  32 - 0x20
      11'h11E: dout <= 8'b00100000; //  286 :  32 - 0x20
      11'h11F: dout <= 8'b00100000; //  287 :  32 - 0x20
      11'h120: dout <= 8'b00101101; //  288 :  45 - 0x2d -- line 0x9
      11'h121: dout <= 8'b00010001; //  289 :  17 - 0x11
      11'h122: dout <= 8'b00000011; //  290 :   3 - 0x3
      11'h123: dout <= 8'b00011110; //  291 :  30 - 0x1e
      11'h124: dout <= 8'b00010000; //  292 :  16 - 0x10
      11'h125: dout <= 8'b00011100; //  293 :  28 - 0x1c
      11'h126: dout <= 8'b00000011; //  294 :   3 - 0x3
      11'h127: dout <= 8'b00010001; //  295 :  17 - 0x11
      11'h128: dout <= 8'b00000011; //  296 :   3 - 0x3
      11'h129: dout <= 8'b00011110; //  297 :  30 - 0x1e
      11'h12A: dout <= 8'b00010000; //  298 :  16 - 0x10
      11'h12B: dout <= 8'b00010011; //  299 :  19 - 0x13
      11'h12C: dout <= 8'b00010000; //  300 :  16 - 0x10
      11'h12D: dout <= 8'b00011100; //  301 :  28 - 0x1c
      11'h12E: dout <= 8'b00000011; //  302 :   3 - 0x3
      11'h12F: dout <= 8'b00010001; //  303 :  17 - 0x11
      11'h130: dout <= 8'b00000011; //  304 :   3 - 0x3
      11'h131: dout <= 8'b00011110; //  305 :  30 - 0x1e
      11'h132: dout <= 8'b00010000; //  306 :  16 - 0x10
      11'h133: dout <= 8'b00011100; //  307 :  28 - 0x1c
      11'h134: dout <= 8'b00000011; //  308 :   3 - 0x3
      11'h135: dout <= 8'b00010001; //  309 :  17 - 0x11
      11'h136: dout <= 8'b00100000; //  310 :  32 - 0x20
      11'h137: dout <= 8'b00100000; //  311 :  32 - 0x20
      11'h138: dout <= 8'b00100000; //  312 :  32 - 0x20
      11'h139: dout <= 8'b00100000; //  313 :  32 - 0x20
      11'h13A: dout <= 8'b00100000; //  314 :  32 - 0x20
      11'h13B: dout <= 8'b00110000; //  315 :  48 - 0x30
      11'h13C: dout <= 8'b00110000; //  316 :  48 - 0x30
      11'h13D: dout <= 8'b00100000; //  317 :  32 - 0x20
      11'h13E: dout <= 8'b00100000; //  318 :  32 - 0x20
      11'h13F: dout <= 8'b00100000; //  319 :  32 - 0x20
      11'h140: dout <= 8'b00101101; //  320 :  45 - 0x2d -- line 0xa
      11'h141: dout <= 8'b00010001; //  321 :  17 - 0x11
      11'h142: dout <= 8'b00000011; //  322 :   3 - 0x3
      11'h143: dout <= 8'b00000011; //  323 :   3 - 0x3
      11'h144: dout <= 8'b00000011; //  324 :   3 - 0x3
      11'h145: dout <= 8'b00000011; //  325 :   3 - 0x3
      11'h146: dout <= 8'b00000011; //  326 :   3 - 0x3
      11'h147: dout <= 8'b00010001; //  327 :  17 - 0x11
      11'h148: dout <= 8'b00000011; //  328 :   3 - 0x3
      11'h149: dout <= 8'b00000011; //  329 :   3 - 0x3
      11'h14A: dout <= 8'b00000011; //  330 :   3 - 0x3
      11'h14B: dout <= 8'b00010001; //  331 :  17 - 0x11
      11'h14C: dout <= 8'b00000011; //  332 :   3 - 0x3
      11'h14D: dout <= 8'b00000011; //  333 :   3 - 0x3
      11'h14E: dout <= 8'b00000011; //  334 :   3 - 0x3
      11'h14F: dout <= 8'b00010001; //  335 :  17 - 0x11
      11'h150: dout <= 8'b00000011; //  336 :   3 - 0x3
      11'h151: dout <= 8'b00000011; //  337 :   3 - 0x3
      11'h152: dout <= 8'b00000011; //  338 :   3 - 0x3
      11'h153: dout <= 8'b00000011; //  339 :   3 - 0x3
      11'h154: dout <= 8'b00000011; //  340 :   3 - 0x3
      11'h155: dout <= 8'b00010001; //  341 :  17 - 0x11
      11'h156: dout <= 8'b00100000; //  342 :  32 - 0x20
      11'h157: dout <= 8'b00100000; //  343 :  32 - 0x20
      11'h158: dout <= 8'b00100000; //  344 :  32 - 0x20
      11'h159: dout <= 8'b00100000; //  345 :  32 - 0x20
      11'h15A: dout <= 8'b00100000; //  346 :  32 - 0x20
      11'h15B: dout <= 8'b00100000; //  347 :  32 - 0x20
      11'h15C: dout <= 8'b00100000; //  348 :  32 - 0x20
      11'h15D: dout <= 8'b00100000; //  349 :  32 - 0x20
      11'h15E: dout <= 8'b00100000; //  350 :  32 - 0x20
      11'h15F: dout <= 8'b00100000; //  351 :  32 - 0x20
      11'h160: dout <= 8'b00101101; //  352 :  45 - 0x2d -- line 0xb
      11'h161: dout <= 8'b00011110; //  353 :  30 - 0x1e
      11'h162: dout <= 8'b00010000; //  354 :  16 - 0x10
      11'h163: dout <= 8'b00010000; //  355 :  16 - 0x10
      11'h164: dout <= 8'b00010000; //  356 :  16 - 0x10
      11'h165: dout <= 8'b00011101; //  357 :  29 - 0x1d
      11'h166: dout <= 8'b00000011; //  358 :   3 - 0x3
      11'h167: dout <= 8'b00010101; //  359 :  21 - 0x15
      11'h168: dout <= 8'b00010000; //  360 :  16 - 0x10
      11'h169: dout <= 8'b00011000; //  361 :  24 - 0x18
      11'h16A: dout <= 8'b00001000; //  362 :   8 - 0x8
      11'h16B: dout <= 8'b00011010; //  363 :  26 - 0x1a
      11'h16C: dout <= 8'b00001000; //  364 :   8 - 0x8
      11'h16D: dout <= 8'b00011001; //  365 :  25 - 0x19
      11'h16E: dout <= 8'b00010000; //  366 :  16 - 0x10
      11'h16F: dout <= 8'b00010100; //  367 :  20 - 0x14
      11'h170: dout <= 8'b00000011; //  368 :   3 - 0x3
      11'h171: dout <= 8'b00011111; //  369 :  31 - 0x1f
      11'h172: dout <= 8'b00010000; //  370 :  16 - 0x10
      11'h173: dout <= 8'b00010000; //  371 :  16 - 0x10
      11'h174: dout <= 8'b00010000; //  372 :  16 - 0x10
      11'h175: dout <= 8'b00011100; //  373 :  28 - 0x1c
      11'h176: dout <= 8'b00100000; //  374 :  32 - 0x20
      11'h177: dout <= 8'b00100000; //  375 :  32 - 0x20
      11'h178: dout <= 8'b00100000; //  376 :  32 - 0x20
      11'h179: dout <= 8'b00100000; //  377 :  32 - 0x20
      11'h17A: dout <= 8'b00100000; //  378 :  32 - 0x20
      11'h17B: dout <= 8'b00100000; //  379 :  32 - 0x20
      11'h17C: dout <= 8'b00100000; //  380 :  32 - 0x20
      11'h17D: dout <= 8'b00100000; //  381 :  32 - 0x20
      11'h17E: dout <= 8'b00100000; //  382 :  32 - 0x20
      11'h17F: dout <= 8'b00100000; //  383 :  32 - 0x20
      11'h180: dout <= 8'b00101101; //  384 :  45 - 0x2d -- line 0xc
      11'h181: dout <= 8'b00100000; //  385 :  32 - 0x20
      11'h182: dout <= 8'b00100000; //  386 :  32 - 0x20
      11'h183: dout <= 8'b00100000; //  387 :  32 - 0x20
      11'h184: dout <= 8'b00100000; //  388 :  32 - 0x20
      11'h185: dout <= 8'b00010001; //  389 :  17 - 0x11
      11'h186: dout <= 8'b00000011; //  390 :   3 - 0x3
      11'h187: dout <= 8'b00010001; //  391 :  17 - 0x11
      11'h188: dout <= 8'b00000000; //  392 :   0 - 0x0
      11'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      11'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      11'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      11'h18F: dout <= 8'b00010001; //  399 :  17 - 0x11
      11'h190: dout <= 8'b00000011; //  400 :   3 - 0x3
      11'h191: dout <= 8'b00010001; //  401 :  17 - 0x11
      11'h192: dout <= 8'b00100000; //  402 :  32 - 0x20
      11'h193: dout <= 8'b00100000; //  403 :  32 - 0x20
      11'h194: dout <= 8'b00100000; //  404 :  32 - 0x20
      11'h195: dout <= 8'b00100000; //  405 :  32 - 0x20
      11'h196: dout <= 8'b00100000; //  406 :  32 - 0x20
      11'h197: dout <= 8'b00100000; //  407 :  32 - 0x20
      11'h198: dout <= 8'b00100000; //  408 :  32 - 0x20
      11'h199: dout <= 8'b00100000; //  409 :  32 - 0x20
      11'h19A: dout <= 8'b00100000; //  410 :  32 - 0x20
      11'h19B: dout <= 8'b00100000; //  411 :  32 - 0x20
      11'h19C: dout <= 8'b00100000; //  412 :  32 - 0x20
      11'h19D: dout <= 8'b00100000; //  413 :  32 - 0x20
      11'h19E: dout <= 8'b00100000; //  414 :  32 - 0x20
      11'h19F: dout <= 8'b00100000; //  415 :  32 - 0x20
      11'h1A0: dout <= 8'b00101101; //  416 :  45 - 0x2d -- line 0xd
      11'h1A1: dout <= 8'b00100000; //  417 :  32 - 0x20
      11'h1A2: dout <= 8'b00100000; //  418 :  32 - 0x20
      11'h1A3: dout <= 8'b00100000; //  419 :  32 - 0x20
      11'h1A4: dout <= 8'b00100000; //  420 :  32 - 0x20
      11'h1A5: dout <= 8'b00010001; //  421 :  17 - 0x11
      11'h1A6: dout <= 8'b00000011; //  422 :   3 - 0x3
      11'h1A7: dout <= 8'b00010001; //  423 :  17 - 0x11
      11'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0
      11'h1A9: dout <= 8'b00011111; //  425 :  31 - 0x1f
      11'h1AA: dout <= 8'b00010111; //  426 :  23 - 0x17
      11'h1AB: dout <= 8'b00101100; //  427 :  44 - 0x2c
      11'h1AC: dout <= 8'b00010110; //  428 :  22 - 0x16
      11'h1AD: dout <= 8'b00011101; //  429 :  29 - 0x1d
      11'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout <= 8'b00010001; //  431 :  17 - 0x11
      11'h1B0: dout <= 8'b00000011; //  432 :   3 - 0x3
      11'h1B1: dout <= 8'b00010001; //  433 :  17 - 0x11
      11'h1B2: dout <= 8'b00100000; //  434 :  32 - 0x20
      11'h1B3: dout <= 8'b00100000; //  435 :  32 - 0x20
      11'h1B4: dout <= 8'b00100000; //  436 :  32 - 0x20
      11'h1B5: dout <= 8'b00100000; //  437 :  32 - 0x20
      11'h1B6: dout <= 8'b00100000; //  438 :  32 - 0x20
      11'h1B7: dout <= 8'b00100000; //  439 :  32 - 0x20
      11'h1B8: dout <= 8'b00100000; //  440 :  32 - 0x20
      11'h1B9: dout <= 8'b00100000; //  441 :  32 - 0x20
      11'h1BA: dout <= 8'b00100000; //  442 :  32 - 0x20
      11'h1BB: dout <= 8'b00100000; //  443 :  32 - 0x20
      11'h1BC: dout <= 8'b00100000; //  444 :  32 - 0x20
      11'h1BD: dout <= 8'b00100000; //  445 :  32 - 0x20
      11'h1BE: dout <= 8'b00100000; //  446 :  32 - 0x20
      11'h1BF: dout <= 8'b00100000; //  447 :  32 - 0x20
      11'h1C0: dout <= 8'b00101101; //  448 :  45 - 0x2d -- line 0xe
      11'h1C1: dout <= 8'b00100010; //  449 :  34 - 0x22
      11'h1C2: dout <= 8'b00010000; //  450 :  16 - 0x10
      11'h1C3: dout <= 8'b00010000; //  451 :  16 - 0x10
      11'h1C4: dout <= 8'b00010000; //  452 :  16 - 0x10
      11'h1C5: dout <= 8'b00011100; //  453 :  28 - 0x1c
      11'h1C6: dout <= 8'b00000011; //  454 :   3 - 0x3
      11'h1C7: dout <= 8'b00011010; //  455 :  26 - 0x1a
      11'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0
      11'h1C9: dout <= 8'b00010001; //  457 :  17 - 0x11
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00010001; //  461 :  17 - 0x11
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00011010; //  463 :  26 - 0x1a
      11'h1D0: dout <= 8'b00000011; //  464 :   3 - 0x3
      11'h1D1: dout <= 8'b00011110; //  465 :  30 - 0x1e
      11'h1D2: dout <= 8'b00010000; //  466 :  16 - 0x10
      11'h1D3: dout <= 8'b00010000; //  467 :  16 - 0x10
      11'h1D4: dout <= 8'b00010000; //  468 :  16 - 0x10
      11'h1D5: dout <= 8'b00100001; //  469 :  33 - 0x21
      11'h1D6: dout <= 8'b00101101; //  470 :  45 - 0x2d
      11'h1D7: dout <= 8'b00101101; //  471 :  45 - 0x2d
      11'h1D8: dout <= 8'b00101101; //  472 :  45 - 0x2d
      11'h1D9: dout <= 8'b00101101; //  473 :  45 - 0x2d
      11'h1DA: dout <= 8'b00101101; //  474 :  45 - 0x2d
      11'h1DB: dout <= 8'b00101101; //  475 :  45 - 0x2d
      11'h1DC: dout <= 8'b00101101; //  476 :  45 - 0x2d
      11'h1DD: dout <= 8'b00101101; //  477 :  45 - 0x2d
      11'h1DE: dout <= 8'b00100000; //  478 :  32 - 0x20
      11'h1DF: dout <= 8'b00100000; //  479 :  32 - 0x20
      11'h1E0: dout <= 8'b00000100; //  480 :   4 - 0x4 -- line 0xf
      11'h1E1: dout <= 8'b00000110; //  481 :   6 - 0x6
      11'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout <= 8'b00000011; //  486 :   3 - 0x3
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0
      11'h1E9: dout <= 8'b00010001; //  489 :  17 - 0x11
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b00010001; //  493 :  17 - 0x11
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b00000011; //  496 :   3 - 0x3
      11'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout <= 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout <= 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout <= 8'b00000101; //  501 :   5 - 0x5
      11'h1F6: dout <= 8'b00000100; //  502 :   4 - 0x4
      11'h1F7: dout <= 8'b00000100; //  503 :   4 - 0x4
      11'h1F8: dout <= 8'b00000100; //  504 :   4 - 0x4
      11'h1F9: dout <= 8'b00000100; //  505 :   4 - 0x4
      11'h1FA: dout <= 8'b00000100; //  506 :   4 - 0x4
      11'h1FB: dout <= 8'b00000100; //  507 :   4 - 0x4
      11'h1FC: dout <= 8'b00000100; //  508 :   4 - 0x4
      11'h1FD: dout <= 8'b00000100; //  509 :   4 - 0x4
      11'h1FE: dout <= 8'b00100000; //  510 :  32 - 0x20
      11'h1FF: dout <= 8'b00100000; //  511 :  32 - 0x20
      11'h200: dout <= 8'b00101101; //  512 :  45 - 0x2d -- line 0x10
      11'h201: dout <= 8'b00100010; //  513 :  34 - 0x22
      11'h202: dout <= 8'b00010000; //  514 :  16 - 0x10
      11'h203: dout <= 8'b00010000; //  515 :  16 - 0x10
      11'h204: dout <= 8'b00010000; //  516 :  16 - 0x10
      11'h205: dout <= 8'b00011101; //  517 :  29 - 0x1d
      11'h206: dout <= 8'b00000011; //  518 :   3 - 0x3
      11'h207: dout <= 8'b00011011; //  519 :  27 - 0x1b
      11'h208: dout <= 8'b00000000; //  520 :   0 - 0x0
      11'h209: dout <= 8'b00011110; //  521 :  30 - 0x1e
      11'h20A: dout <= 8'b00010000; //  522 :  16 - 0x10
      11'h20B: dout <= 8'b00010000; //  523 :  16 - 0x10
      11'h20C: dout <= 8'b00010000; //  524 :  16 - 0x10
      11'h20D: dout <= 8'b00011100; //  525 :  28 - 0x1c
      11'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      11'h20F: dout <= 8'b00011011; //  527 :  27 - 0x1b
      11'h210: dout <= 8'b00000011; //  528 :   3 - 0x3
      11'h211: dout <= 8'b00011111; //  529 :  31 - 0x1f
      11'h212: dout <= 8'b00010000; //  530 :  16 - 0x10
      11'h213: dout <= 8'b00010000; //  531 :  16 - 0x10
      11'h214: dout <= 8'b00010000; //  532 :  16 - 0x10
      11'h215: dout <= 8'b00100001; //  533 :  33 - 0x21
      11'h216: dout <= 8'b00101101; //  534 :  45 - 0x2d
      11'h217: dout <= 8'b00101101; //  535 :  45 - 0x2d
      11'h218: dout <= 8'b00101101; //  536 :  45 - 0x2d
      11'h219: dout <= 8'b00101101; //  537 :  45 - 0x2d
      11'h21A: dout <= 8'b00101101; //  538 :  45 - 0x2d
      11'h21B: dout <= 8'b00101101; //  539 :  45 - 0x2d
      11'h21C: dout <= 8'b00101101; //  540 :  45 - 0x2d
      11'h21D: dout <= 8'b00101101; //  541 :  45 - 0x2d
      11'h21E: dout <= 8'b00100000; //  542 :  32 - 0x20
      11'h21F: dout <= 8'b00100000; //  543 :  32 - 0x20
      11'h220: dout <= 8'b00101101; //  544 :  45 - 0x2d -- line 0x11
      11'h221: dout <= 8'b00100000; //  545 :  32 - 0x20
      11'h222: dout <= 8'b00100000; //  546 :  32 - 0x20
      11'h223: dout <= 8'b00100000; //  547 :  32 - 0x20
      11'h224: dout <= 8'b00100000; //  548 :  32 - 0x20
      11'h225: dout <= 8'b00010001; //  549 :  17 - 0x11
      11'h226: dout <= 8'b00000011; //  550 :   3 - 0x3
      11'h227: dout <= 8'b00010001; //  551 :  17 - 0x11
      11'h228: dout <= 8'b00000000; //  552 :   0 - 0x0
      11'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      11'h22A: dout <= 8'b00000000; //  554 :   0 - 0x0
      11'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      11'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      11'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout <= 8'b00010001; //  559 :  17 - 0x11
      11'h230: dout <= 8'b00000011; //  560 :   3 - 0x3
      11'h231: dout <= 8'b00010001; //  561 :  17 - 0x11
      11'h232: dout <= 8'b00100000; //  562 :  32 - 0x20
      11'h233: dout <= 8'b00100000; //  563 :  32 - 0x20
      11'h234: dout <= 8'b00100000; //  564 :  32 - 0x20
      11'h235: dout <= 8'b00100000; //  565 :  32 - 0x20
      11'h236: dout <= 8'b00100000; //  566 :  32 - 0x20
      11'h237: dout <= 8'b00100000; //  567 :  32 - 0x20
      11'h238: dout <= 8'b00100000; //  568 :  32 - 0x20
      11'h239: dout <= 8'b00100000; //  569 :  32 - 0x20
      11'h23A: dout <= 8'b00100000; //  570 :  32 - 0x20
      11'h23B: dout <= 8'b00100000; //  571 :  32 - 0x20
      11'h23C: dout <= 8'b00100000; //  572 :  32 - 0x20
      11'h23D: dout <= 8'b00100000; //  573 :  32 - 0x20
      11'h23E: dout <= 8'b00100000; //  574 :  32 - 0x20
      11'h23F: dout <= 8'b00100000; //  575 :  32 - 0x20
      11'h240: dout <= 8'b00101101; //  576 :  45 - 0x2d -- line 0x12
      11'h241: dout <= 8'b00100000; //  577 :  32 - 0x20
      11'h242: dout <= 8'b00100000; //  578 :  32 - 0x20
      11'h243: dout <= 8'b00100000; //  579 :  32 - 0x20
      11'h244: dout <= 8'b00100000; //  580 :  32 - 0x20
      11'h245: dout <= 8'b00010001; //  581 :  17 - 0x11
      11'h246: dout <= 8'b00000011; //  582 :   3 - 0x3
      11'h247: dout <= 8'b00010001; //  583 :  17 - 0x11
      11'h248: dout <= 8'b00000000; //  584 :   0 - 0x0
      11'h249: dout <= 8'b00011111; //  585 :  31 - 0x1f
      11'h24A: dout <= 8'b00010000; //  586 :  16 - 0x10
      11'h24B: dout <= 8'b00010000; //  587 :  16 - 0x10
      11'h24C: dout <= 8'b00010000; //  588 :  16 - 0x10
      11'h24D: dout <= 8'b00011101; //  589 :  29 - 0x1d
      11'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout <= 8'b00010001; //  591 :  17 - 0x11
      11'h250: dout <= 8'b00000011; //  592 :   3 - 0x3
      11'h251: dout <= 8'b00010001; //  593 :  17 - 0x11
      11'h252: dout <= 8'b00100000; //  594 :  32 - 0x20
      11'h253: dout <= 8'b00100000; //  595 :  32 - 0x20
      11'h254: dout <= 8'b00100000; //  596 :  32 - 0x20
      11'h255: dout <= 8'b00100000; //  597 :  32 - 0x20
      11'h256: dout <= 8'b01100000; //  598 :  96 - 0x60
      11'h257: dout <= 8'b01100001; //  599 :  97 - 0x61
      11'h258: dout <= 8'b00100000; //  600 :  32 - 0x20
      11'h259: dout <= 8'b00100000; //  601 :  32 - 0x20
      11'h25A: dout <= 8'b00100000; //  602 :  32 - 0x20
      11'h25B: dout <= 8'b00100000; //  603 :  32 - 0x20
      11'h25C: dout <= 8'b00101101; //  604 :  45 - 0x2d
      11'h25D: dout <= 8'b00101101; //  605 :  45 - 0x2d
      11'h25E: dout <= 8'b00100000; //  606 :  32 - 0x20
      11'h25F: dout <= 8'b00100000; //  607 :  32 - 0x20
      11'h260: dout <= 8'b00101101; //  608 :  45 - 0x2d -- line 0x13
      11'h261: dout <= 8'b00011111; //  609 :  31 - 0x1f
      11'h262: dout <= 8'b00010000; //  610 :  16 - 0x10
      11'h263: dout <= 8'b00010000; //  611 :  16 - 0x10
      11'h264: dout <= 8'b00010000; //  612 :  16 - 0x10
      11'h265: dout <= 8'b00011100; //  613 :  28 - 0x1c
      11'h266: dout <= 8'b00000011; //  614 :   3 - 0x3
      11'h267: dout <= 8'b00011010; //  615 :  26 - 0x1a
      11'h268: dout <= 8'b00000000; //  616 :   0 - 0x0
      11'h269: dout <= 8'b00011110; //  617 :  30 - 0x1e
      11'h26A: dout <= 8'b00010000; //  618 :  16 - 0x10
      11'h26B: dout <= 8'b00010011; //  619 :  19 - 0x13
      11'h26C: dout <= 8'b00010000; //  620 :  16 - 0x10
      11'h26D: dout <= 8'b00011100; //  621 :  28 - 0x1c
      11'h26E: dout <= 8'b00000000; //  622 :   0 - 0x0
      11'h26F: dout <= 8'b00011010; //  623 :  26 - 0x1a
      11'h270: dout <= 8'b00000011; //  624 :   3 - 0x3
      11'h271: dout <= 8'b00011110; //  625 :  30 - 0x1e
      11'h272: dout <= 8'b00010000; //  626 :  16 - 0x10
      11'h273: dout <= 8'b00010000; //  627 :  16 - 0x10
      11'h274: dout <= 8'b00010000; //  628 :  16 - 0x10
      11'h275: dout <= 8'b00011101; //  629 :  29 - 0x1d
      11'h276: dout <= 8'b01100010; //  630 :  98 - 0x62
      11'h277: dout <= 8'b01100011; //  631 :  99 - 0x63
      11'h278: dout <= 8'b00100000; //  632 :  32 - 0x20
      11'h279: dout <= 8'b00100000; //  633 :  32 - 0x20
      11'h27A: dout <= 8'b00100000; //  634 :  32 - 0x20
      11'h27B: dout <= 8'b00100000; //  635 :  32 - 0x20
      11'h27C: dout <= 8'b00101101; //  636 :  45 - 0x2d
      11'h27D: dout <= 8'b00101101; //  637 :  45 - 0x2d
      11'h27E: dout <= 8'b00100000; //  638 :  32 - 0x20
      11'h27F: dout <= 8'b00100000; //  639 :  32 - 0x20
      11'h280: dout <= 8'b00101101; //  640 :  45 - 0x2d -- line 0x14
      11'h281: dout <= 8'b00010001; //  641 :  17 - 0x11
      11'h282: dout <= 8'b00000011; //  642 :   3 - 0x3
      11'h283: dout <= 8'b00000011; //  643 :   3 - 0x3
      11'h284: dout <= 8'b00000011; //  644 :   3 - 0x3
      11'h285: dout <= 8'b00000011; //  645 :   3 - 0x3
      11'h286: dout <= 8'b00000011; //  646 :   3 - 0x3
      11'h287: dout <= 8'b00000011; //  647 :   3 - 0x3
      11'h288: dout <= 8'b00000011; //  648 :   3 - 0x3
      11'h289: dout <= 8'b00000011; //  649 :   3 - 0x3
      11'h28A: dout <= 8'b00000011; //  650 :   3 - 0x3
      11'h28B: dout <= 8'b00010001; //  651 :  17 - 0x11
      11'h28C: dout <= 8'b00000011; //  652 :   3 - 0x3
      11'h28D: dout <= 8'b00000011; //  653 :   3 - 0x3
      11'h28E: dout <= 8'b00000011; //  654 :   3 - 0x3
      11'h28F: dout <= 8'b00000011; //  655 :   3 - 0x3
      11'h290: dout <= 8'b00000011; //  656 :   3 - 0x3
      11'h291: dout <= 8'b00000011; //  657 :   3 - 0x3
      11'h292: dout <= 8'b00000011; //  658 :   3 - 0x3
      11'h293: dout <= 8'b00000011; //  659 :   3 - 0x3
      11'h294: dout <= 8'b00000011; //  660 :   3 - 0x3
      11'h295: dout <= 8'b00010001; //  661 :  17 - 0x11
      11'h296: dout <= 8'b00100000; //  662 :  32 - 0x20
      11'h297: dout <= 8'b00100000; //  663 :  32 - 0x20
      11'h298: dout <= 8'b00100000; //  664 :  32 - 0x20
      11'h299: dout <= 8'b00100000; //  665 :  32 - 0x20
      11'h29A: dout <= 8'b00100000; //  666 :  32 - 0x20
      11'h29B: dout <= 8'b00100000; //  667 :  32 - 0x20
      11'h29C: dout <= 8'b00101101; //  668 :  45 - 0x2d
      11'h29D: dout <= 8'b00101101; //  669 :  45 - 0x2d
      11'h29E: dout <= 8'b00100000; //  670 :  32 - 0x20
      11'h29F: dout <= 8'b00100000; //  671 :  32 - 0x20
      11'h2A0: dout <= 8'b00101101; //  672 :  45 - 0x2d -- line 0x15
      11'h2A1: dout <= 8'b00010001; //  673 :  17 - 0x11
      11'h2A2: dout <= 8'b00000011; //  674 :   3 - 0x3
      11'h2A3: dout <= 8'b00011001; //  675 :  25 - 0x19
      11'h2A4: dout <= 8'b00010000; //  676 :  16 - 0x10
      11'h2A5: dout <= 8'b00011101; //  677 :  29 - 0x1d
      11'h2A6: dout <= 8'b00000011; //  678 :   3 - 0x3
      11'h2A7: dout <= 8'b00011001; //  679 :  25 - 0x19
      11'h2A8: dout <= 8'b00010000; //  680 :  16 - 0x10
      11'h2A9: dout <= 8'b00011000; //  681 :  24 - 0x18
      11'h2AA: dout <= 8'b00001001; //  682 :   9 - 0x9
      11'h2AB: dout <= 8'b00011010; //  683 :  26 - 0x1a
      11'h2AC: dout <= 8'b00001001; //  684 :   9 - 0x9
      11'h2AD: dout <= 8'b00011001; //  685 :  25 - 0x19
      11'h2AE: dout <= 8'b00010000; //  686 :  16 - 0x10
      11'h2AF: dout <= 8'b00011000; //  687 :  24 - 0x18
      11'h2B0: dout <= 8'b00000011; //  688 :   3 - 0x3
      11'h2B1: dout <= 8'b00011111; //  689 :  31 - 0x1f
      11'h2B2: dout <= 8'b00010000; //  690 :  16 - 0x10
      11'h2B3: dout <= 8'b00011000; //  691 :  24 - 0x18
      11'h2B4: dout <= 8'b00000011; //  692 :   3 - 0x3
      11'h2B5: dout <= 8'b00010001; //  693 :  17 - 0x11
      11'h2B6: dout <= 8'b00100000; //  694 :  32 - 0x20
      11'h2B7: dout <= 8'b00100000; //  695 :  32 - 0x20
      11'h2B8: dout <= 8'b00100000; //  696 :  32 - 0x20
      11'h2B9: dout <= 8'b00100000; //  697 :  32 - 0x20
      11'h2BA: dout <= 8'b00100000; //  698 :  32 - 0x20
      11'h2BB: dout <= 8'b00100000; //  699 :  32 - 0x20
      11'h2BC: dout <= 8'b00101101; //  700 :  45 - 0x2d
      11'h2BD: dout <= 8'b00101101; //  701 :  45 - 0x2d
      11'h2BE: dout <= 8'b00100000; //  702 :  32 - 0x20
      11'h2BF: dout <= 8'b00100000; //  703 :  32 - 0x20
      11'h2C0: dout <= 8'b00101101; //  704 :  45 - 0x2d -- line 0x16
      11'h2C1: dout <= 8'b00010001; //  705 :  17 - 0x11
      11'h2C2: dout <= 8'b00000001; //  706 :   1 - 0x1
      11'h2C3: dout <= 8'b00000011; //  707 :   3 - 0x3
      11'h2C4: dout <= 8'b00000011; //  708 :   3 - 0x3
      11'h2C5: dout <= 8'b00010001; //  709 :  17 - 0x11
      11'h2C6: dout <= 8'b00000011; //  710 :   3 - 0x3
      11'h2C7: dout <= 8'b00000011; //  711 :   3 - 0x3
      11'h2C8: dout <= 8'b00000011; //  712 :   3 - 0x3
      11'h2C9: dout <= 8'b00000011; //  713 :   3 - 0x3
      11'h2CA: dout <= 8'b00000011; //  714 :   3 - 0x3
      11'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      11'h2CC: dout <= 8'b00000011; //  716 :   3 - 0x3
      11'h2CD: dout <= 8'b00000011; //  717 :   3 - 0x3
      11'h2CE: dout <= 8'b00000011; //  718 :   3 - 0x3
      11'h2CF: dout <= 8'b00000011; //  719 :   3 - 0x3
      11'h2D0: dout <= 8'b00000011; //  720 :   3 - 0x3
      11'h2D1: dout <= 8'b00010001; //  721 :  17 - 0x11
      11'h2D2: dout <= 8'b00000011; //  722 :   3 - 0x3
      11'h2D3: dout <= 8'b00000011; //  723 :   3 - 0x3
      11'h2D4: dout <= 8'b00000001; //  724 :   1 - 0x1
      11'h2D5: dout <= 8'b00010001; //  725 :  17 - 0x11
      11'h2D6: dout <= 8'b00100000; //  726 :  32 - 0x20
      11'h2D7: dout <= 8'b00100000; //  727 :  32 - 0x20
      11'h2D8: dout <= 8'b00100000; //  728 :  32 - 0x20
      11'h2D9: dout <= 8'b00100000; //  729 :  32 - 0x20
      11'h2DA: dout <= 8'b00100000; //  730 :  32 - 0x20
      11'h2DB: dout <= 8'b00100000; //  731 :  32 - 0x20
      11'h2DC: dout <= 8'b00101101; //  732 :  45 - 0x2d
      11'h2DD: dout <= 8'b00101101; //  733 :  45 - 0x2d
      11'h2DE: dout <= 8'b00100000; //  734 :  32 - 0x20
      11'h2DF: dout <= 8'b00100000; //  735 :  32 - 0x20
      11'h2E0: dout <= 8'b00101101; //  736 :  45 - 0x2d -- line 0x17
      11'h2E1: dout <= 8'b00010101; //  737 :  21 - 0x15
      11'h2E2: dout <= 8'b00010000; //  738 :  16 - 0x10
      11'h2E3: dout <= 8'b00011101; //  739 :  29 - 0x1d
      11'h2E4: dout <= 8'b00000011; //  740 :   3 - 0x3
      11'h2E5: dout <= 8'b00010001; //  741 :  17 - 0x11
      11'h2E6: dout <= 8'b00000011; //  742 :   3 - 0x3
      11'h2E7: dout <= 8'b00011011; //  743 :  27 - 0x1b
      11'h2E8: dout <= 8'b00000011; //  744 :   3 - 0x3
      11'h2E9: dout <= 8'b00011111; //  745 :  31 - 0x1f
      11'h2EA: dout <= 8'b00010000; //  746 :  16 - 0x10
      11'h2EB: dout <= 8'b00010000; //  747 :  16 - 0x10
      11'h2EC: dout <= 8'b00010000; //  748 :  16 - 0x10
      11'h2ED: dout <= 8'b00011101; //  749 :  29 - 0x1d
      11'h2EE: dout <= 8'b00000011; //  750 :   3 - 0x3
      11'h2EF: dout <= 8'b00011011; //  751 :  27 - 0x1b
      11'h2F0: dout <= 8'b00000011; //  752 :   3 - 0x3
      11'h2F1: dout <= 8'b00010001; //  753 :  17 - 0x11
      11'h2F2: dout <= 8'b00000011; //  754 :   3 - 0x3
      11'h2F3: dout <= 8'b00011111; //  755 :  31 - 0x1f
      11'h2F4: dout <= 8'b00010000; //  756 :  16 - 0x10
      11'h2F5: dout <= 8'b00010100; //  757 :  20 - 0x14
      11'h2F6: dout <= 8'b00100000; //  758 :  32 - 0x20
      11'h2F7: dout <= 8'b00100000; //  759 :  32 - 0x20
      11'h2F8: dout <= 8'b00100000; //  760 :  32 - 0x20
      11'h2F9: dout <= 8'b00100000; //  761 :  32 - 0x20
      11'h2FA: dout <= 8'b00100000; //  762 :  32 - 0x20
      11'h2FB: dout <= 8'b00100000; //  763 :  32 - 0x20
      11'h2FC: dout <= 8'b00101101; //  764 :  45 - 0x2d
      11'h2FD: dout <= 8'b00101101; //  765 :  45 - 0x2d
      11'h2FE: dout <= 8'b00100000; //  766 :  32 - 0x20
      11'h2FF: dout <= 8'b00100000; //  767 :  32 - 0x20
      11'h300: dout <= 8'b00101101; //  768 :  45 - 0x2d -- line 0x18
      11'h301: dout <= 8'b00010101; //  769 :  21 - 0x15
      11'h302: dout <= 8'b00010000; //  770 :  16 - 0x10
      11'h303: dout <= 8'b00011100; //  771 :  28 - 0x1c
      11'h304: dout <= 8'b00000011; //  772 :   3 - 0x3
      11'h305: dout <= 8'b00011010; //  773 :  26 - 0x1a
      11'h306: dout <= 8'b00000011; //  774 :   3 - 0x3
      11'h307: dout <= 8'b00010001; //  775 :  17 - 0x11
      11'h308: dout <= 8'b00000011; //  776 :   3 - 0x3
      11'h309: dout <= 8'b00011110; //  777 :  30 - 0x1e
      11'h30A: dout <= 8'b00010000; //  778 :  16 - 0x10
      11'h30B: dout <= 8'b00010011; //  779 :  19 - 0x13
      11'h30C: dout <= 8'b00010000; //  780 :  16 - 0x10
      11'h30D: dout <= 8'b00011100; //  781 :  28 - 0x1c
      11'h30E: dout <= 8'b00000011; //  782 :   3 - 0x3
      11'h30F: dout <= 8'b00010001; //  783 :  17 - 0x11
      11'h310: dout <= 8'b00000011; //  784 :   3 - 0x3
      11'h311: dout <= 8'b00011010; //  785 :  26 - 0x1a
      11'h312: dout <= 8'b00000011; //  786 :   3 - 0x3
      11'h313: dout <= 8'b00011110; //  787 :  30 - 0x1e
      11'h314: dout <= 8'b00010000; //  788 :  16 - 0x10
      11'h315: dout <= 8'b00010100; //  789 :  20 - 0x14
      11'h316: dout <= 8'b00100000; //  790 :  32 - 0x20
      11'h317: dout <= 8'b00111100; //  791 :  60 - 0x3c
      11'h318: dout <= 8'b00111101; //  792 :  61 - 0x3d
      11'h319: dout <= 8'b00111100; //  793 :  60 - 0x3c
      11'h31A: dout <= 8'b00111101; //  794 :  61 - 0x3d
      11'h31B: dout <= 8'b00101101; //  795 :  45 - 0x2d
      11'h31C: dout <= 8'b00101101; //  796 :  45 - 0x2d
      11'h31D: dout <= 8'b00101101; //  797 :  45 - 0x2d
      11'h31E: dout <= 8'b00100000; //  798 :  32 - 0x20
      11'h31F: dout <= 8'b00100000; //  799 :  32 - 0x20
      11'h320: dout <= 8'b00101101; //  800 :  45 - 0x2d -- line 0x19
      11'h321: dout <= 8'b00010001; //  801 :  17 - 0x11
      11'h322: dout <= 8'b00000011; //  802 :   3 - 0x3
      11'h323: dout <= 8'b00000011; //  803 :   3 - 0x3
      11'h324: dout <= 8'b00000011; //  804 :   3 - 0x3
      11'h325: dout <= 8'b00000011; //  805 :   3 - 0x3
      11'h326: dout <= 8'b00000011; //  806 :   3 - 0x3
      11'h327: dout <= 8'b00010001; //  807 :  17 - 0x11
      11'h328: dout <= 8'b00000011; //  808 :   3 - 0x3
      11'h329: dout <= 8'b00000011; //  809 :   3 - 0x3
      11'h32A: dout <= 8'b00000011; //  810 :   3 - 0x3
      11'h32B: dout <= 8'b00010001; //  811 :  17 - 0x11
      11'h32C: dout <= 8'b00000011; //  812 :   3 - 0x3
      11'h32D: dout <= 8'b00000011; //  813 :   3 - 0x3
      11'h32E: dout <= 8'b00000011; //  814 :   3 - 0x3
      11'h32F: dout <= 8'b00010001; //  815 :  17 - 0x11
      11'h330: dout <= 8'b00000011; //  816 :   3 - 0x3
      11'h331: dout <= 8'b00000011; //  817 :   3 - 0x3
      11'h332: dout <= 8'b00000011; //  818 :   3 - 0x3
      11'h333: dout <= 8'b00000011; //  819 :   3 - 0x3
      11'h334: dout <= 8'b00000011; //  820 :   3 - 0x3
      11'h335: dout <= 8'b00010001; //  821 :  17 - 0x11
      11'h336: dout <= 8'b00100000; //  822 :  32 - 0x20
      11'h337: dout <= 8'b00111110; //  823 :  62 - 0x3e
      11'h338: dout <= 8'b00111111; //  824 :  63 - 0x3f
      11'h339: dout <= 8'b00111110; //  825 :  62 - 0x3e
      11'h33A: dout <= 8'b00111111; //  826 :  63 - 0x3f
      11'h33B: dout <= 8'b00101101; //  827 :  45 - 0x2d
      11'h33C: dout <= 8'b00101101; //  828 :  45 - 0x2d
      11'h33D: dout <= 8'b00101101; //  829 :  45 - 0x2d
      11'h33E: dout <= 8'b00100000; //  830 :  32 - 0x20
      11'h33F: dout <= 8'b00100000; //  831 :  32 - 0x20
      11'h340: dout <= 8'b00101101; //  832 :  45 - 0x2d -- line 0x1a
      11'h341: dout <= 8'b00010001; //  833 :  17 - 0x11
      11'h342: dout <= 8'b00000011; //  834 :   3 - 0x3
      11'h343: dout <= 8'b00011001; //  835 :  25 - 0x19
      11'h344: dout <= 8'b00010000; //  836 :  16 - 0x10
      11'h345: dout <= 8'b00010000; //  837 :  16 - 0x10
      11'h346: dout <= 8'b00010000; //  838 :  16 - 0x10
      11'h347: dout <= 8'b00010010; //  839 :  18 - 0x12
      11'h348: dout <= 8'b00010000; //  840 :  16 - 0x10
      11'h349: dout <= 8'b00011000; //  841 :  24 - 0x18
      11'h34A: dout <= 8'b00000011; //  842 :   3 - 0x3
      11'h34B: dout <= 8'b00011010; //  843 :  26 - 0x1a
      11'h34C: dout <= 8'b00000011; //  844 :   3 - 0x3
      11'h34D: dout <= 8'b00011001; //  845 :  25 - 0x19
      11'h34E: dout <= 8'b00010000; //  846 :  16 - 0x10
      11'h34F: dout <= 8'b00010010; //  847 :  18 - 0x12
      11'h350: dout <= 8'b00010000; //  848 :  16 - 0x10
      11'h351: dout <= 8'b00010000; //  849 :  16 - 0x10
      11'h352: dout <= 8'b00010000; //  850 :  16 - 0x10
      11'h353: dout <= 8'b00011000; //  851 :  24 - 0x18
      11'h354: dout <= 8'b00000011; //  852 :   3 - 0x3
      11'h355: dout <= 8'b00010001; //  853 :  17 - 0x11
      11'h356: dout <= 8'b00100000; //  854 :  32 - 0x20
      11'h357: dout <= 8'b00100000; //  855 :  32 - 0x20
      11'h358: dout <= 8'b00100000; //  856 :  32 - 0x20
      11'h359: dout <= 8'b00100000; //  857 :  32 - 0x20
      11'h35A: dout <= 8'b00100000; //  858 :  32 - 0x20
      11'h35B: dout <= 8'b00100000; //  859 :  32 - 0x20
      11'h35C: dout <= 8'b00101101; //  860 :  45 - 0x2d
      11'h35D: dout <= 8'b00101101; //  861 :  45 - 0x2d
      11'h35E: dout <= 8'b00100000; //  862 :  32 - 0x20
      11'h35F: dout <= 8'b00100000; //  863 :  32 - 0x20
      11'h360: dout <= 8'b00101101; //  864 :  45 - 0x2d -- line 0x1b
      11'h361: dout <= 8'b00010001; //  865 :  17 - 0x11
      11'h362: dout <= 8'b00000011; //  866 :   3 - 0x3
      11'h363: dout <= 8'b00000011; //  867 :   3 - 0x3
      11'h364: dout <= 8'b00000011; //  868 :   3 - 0x3
      11'h365: dout <= 8'b00000011; //  869 :   3 - 0x3
      11'h366: dout <= 8'b00000011; //  870 :   3 - 0x3
      11'h367: dout <= 8'b00000011; //  871 :   3 - 0x3
      11'h368: dout <= 8'b00000011; //  872 :   3 - 0x3
      11'h369: dout <= 8'b00000011; //  873 :   3 - 0x3
      11'h36A: dout <= 8'b00000011; //  874 :   3 - 0x3
      11'h36B: dout <= 8'b00000011; //  875 :   3 - 0x3
      11'h36C: dout <= 8'b00000011; //  876 :   3 - 0x3
      11'h36D: dout <= 8'b00000011; //  877 :   3 - 0x3
      11'h36E: dout <= 8'b00000011; //  878 :   3 - 0x3
      11'h36F: dout <= 8'b00000011; //  879 :   3 - 0x3
      11'h370: dout <= 8'b00000011; //  880 :   3 - 0x3
      11'h371: dout <= 8'b00000011; //  881 :   3 - 0x3
      11'h372: dout <= 8'b00000011; //  882 :   3 - 0x3
      11'h373: dout <= 8'b00000011; //  883 :   3 - 0x3
      11'h374: dout <= 8'b00000011; //  884 :   3 - 0x3
      11'h375: dout <= 8'b00010001; //  885 :  17 - 0x11
      11'h376: dout <= 8'b00100000; //  886 :  32 - 0x20
      11'h377: dout <= 8'b00100000; //  887 :  32 - 0x20
      11'h378: dout <= 8'b00100000; //  888 :  32 - 0x20
      11'h379: dout <= 8'b00100000; //  889 :  32 - 0x20
      11'h37A: dout <= 8'b00100000; //  890 :  32 - 0x20
      11'h37B: dout <= 8'b00100000; //  891 :  32 - 0x20
      11'h37C: dout <= 8'b00101101; //  892 :  45 - 0x2d
      11'h37D: dout <= 8'b00101101; //  893 :  45 - 0x2d
      11'h37E: dout <= 8'b00100000; //  894 :  32 - 0x20
      11'h37F: dout <= 8'b00100000; //  895 :  32 - 0x20
      11'h380: dout <= 8'b00101101; //  896 :  45 - 0x2d -- line 0x1c
      11'h381: dout <= 8'b00011110; //  897 :  30 - 0x1e
      11'h382: dout <= 8'b00010000; //  898 :  16 - 0x10
      11'h383: dout <= 8'b00010000; //  899 :  16 - 0x10
      11'h384: dout <= 8'b00010000; //  900 :  16 - 0x10
      11'h385: dout <= 8'b00010000; //  901 :  16 - 0x10
      11'h386: dout <= 8'b00010000; //  902 :  16 - 0x10
      11'h387: dout <= 8'b00010000; //  903 :  16 - 0x10
      11'h388: dout <= 8'b00010000; //  904 :  16 - 0x10
      11'h389: dout <= 8'b00010000; //  905 :  16 - 0x10
      11'h38A: dout <= 8'b00010000; //  906 :  16 - 0x10
      11'h38B: dout <= 8'b00010000; //  907 :  16 - 0x10
      11'h38C: dout <= 8'b00010000; //  908 :  16 - 0x10
      11'h38D: dout <= 8'b00010000; //  909 :  16 - 0x10
      11'h38E: dout <= 8'b00010000; //  910 :  16 - 0x10
      11'h38F: dout <= 8'b00010000; //  911 :  16 - 0x10
      11'h390: dout <= 8'b00010000; //  912 :  16 - 0x10
      11'h391: dout <= 8'b00010000; //  913 :  16 - 0x10
      11'h392: dout <= 8'b00010000; //  914 :  16 - 0x10
      11'h393: dout <= 8'b00010000; //  915 :  16 - 0x10
      11'h394: dout <= 8'b00010000; //  916 :  16 - 0x10
      11'h395: dout <= 8'b00011100; //  917 :  28 - 0x1c
      11'h396: dout <= 8'b00100000; //  918 :  32 - 0x20
      11'h397: dout <= 8'b00100000; //  919 :  32 - 0x20
      11'h398: dout <= 8'b00100000; //  920 :  32 - 0x20
      11'h399: dout <= 8'b00100000; //  921 :  32 - 0x20
      11'h39A: dout <= 8'b00100000; //  922 :  32 - 0x20
      11'h39B: dout <= 8'b00100000; //  923 :  32 - 0x20
      11'h39C: dout <= 8'b00100000; //  924 :  32 - 0x20
      11'h39D: dout <= 8'b00100000; //  925 :  32 - 0x20
      11'h39E: dout <= 8'b00100000; //  926 :  32 - 0x20
      11'h39F: dout <= 8'b00100000; //  927 :  32 - 0x20
      11'h3A0: dout <= 8'b00100000; //  928 :  32 - 0x20 -- line 0x1d
      11'h3A1: dout <= 8'b00100000; //  929 :  32 - 0x20
      11'h3A2: dout <= 8'b00100000; //  930 :  32 - 0x20
      11'h3A3: dout <= 8'b00100000; //  931 :  32 - 0x20
      11'h3A4: dout <= 8'b00100000; //  932 :  32 - 0x20
      11'h3A5: dout <= 8'b00100000; //  933 :  32 - 0x20
      11'h3A6: dout <= 8'b00100000; //  934 :  32 - 0x20
      11'h3A7: dout <= 8'b00100000; //  935 :  32 - 0x20
      11'h3A8: dout <= 8'b00100000; //  936 :  32 - 0x20
      11'h3A9: dout <= 8'b00100000; //  937 :  32 - 0x20
      11'h3AA: dout <= 8'b00100000; //  938 :  32 - 0x20
      11'h3AB: dout <= 8'b00100000; //  939 :  32 - 0x20
      11'h3AC: dout <= 8'b00100000; //  940 :  32 - 0x20
      11'h3AD: dout <= 8'b00100000; //  941 :  32 - 0x20
      11'h3AE: dout <= 8'b00100000; //  942 :  32 - 0x20
      11'h3AF: dout <= 8'b00100000; //  943 :  32 - 0x20
      11'h3B0: dout <= 8'b00100000; //  944 :  32 - 0x20
      11'h3B1: dout <= 8'b00100000; //  945 :  32 - 0x20
      11'h3B2: dout <= 8'b00100000; //  946 :  32 - 0x20
      11'h3B3: dout <= 8'b00100000; //  947 :  32 - 0x20
      11'h3B4: dout <= 8'b00100000; //  948 :  32 - 0x20
      11'h3B5: dout <= 8'b00100000; //  949 :  32 - 0x20
      11'h3B6: dout <= 8'b00100000; //  950 :  32 - 0x20
      11'h3B7: dout <= 8'b00100000; //  951 :  32 - 0x20
      11'h3B8: dout <= 8'b00100000; //  952 :  32 - 0x20
      11'h3B9: dout <= 8'b00100000; //  953 :  32 - 0x20
      11'h3BA: dout <= 8'b00100000; //  954 :  32 - 0x20
      11'h3BB: dout <= 8'b00100000; //  955 :  32 - 0x20
      11'h3BC: dout <= 8'b00100000; //  956 :  32 - 0x20
      11'h3BD: dout <= 8'b00100000; //  957 :  32 - 0x20
      11'h3BE: dout <= 8'b00100000; //  958 :  32 - 0x20
      11'h3BF: dout <= 8'b00100000; //  959 :  32 - 0x20
        //-- Attribute Table 0----
      11'h3C0: dout <= 8'b01010101; //  960 :  85 - 0x55
      11'h3C1: dout <= 8'b01010101; //  961 :  85 - 0x55
      11'h3C2: dout <= 8'b01010101; //  962 :  85 - 0x55
      11'h3C3: dout <= 8'b01010101; //  963 :  85 - 0x55
      11'h3C4: dout <= 8'b01010101; //  964 :  85 - 0x55
      11'h3C5: dout <= 8'b00010001; //  965 :  17 - 0x11
      11'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout <= 8'b01010101; //  968 :  85 - 0x55
      11'h3C9: dout <= 8'b01010101; //  969 :  85 - 0x55
      11'h3CA: dout <= 8'b01010101; //  970 :  85 - 0x55
      11'h3CB: dout <= 8'b01010101; //  971 :  85 - 0x55
      11'h3CC: dout <= 8'b01010101; //  972 :  85 - 0x55
      11'h3CD: dout <= 8'b00010001; //  973 :  17 - 0x11
      11'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout <= 8'b01010101; //  976 :  85 - 0x55
      11'h3D1: dout <= 8'b01010101; //  977 :  85 - 0x55
      11'h3D2: dout <= 8'b01010101; //  978 :  85 - 0x55
      11'h3D3: dout <= 8'b01010101; //  979 :  85 - 0x55
      11'h3D4: dout <= 8'b01010101; //  980 :  85 - 0x55
      11'h3D5: dout <= 8'b00010001; //  981 :  17 - 0x11
      11'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout <= 8'b01010101; //  984 :  85 - 0x55
      11'h3D9: dout <= 8'b01010101; //  985 :  85 - 0x55
      11'h3DA: dout <= 8'b01010101; //  986 :  85 - 0x55
      11'h3DB: dout <= 8'b01010101; //  987 :  85 - 0x55
      11'h3DC: dout <= 8'b01010101; //  988 :  85 - 0x55
      11'h3DD: dout <= 8'b01010001; //  989 :  81 - 0x51
      11'h3DE: dout <= 8'b01010000; //  990 :  80 - 0x50
      11'h3DF: dout <= 8'b01010000; //  991 :  80 - 0x50
      11'h3E0: dout <= 8'b01010101; //  992 :  85 - 0x55
      11'h3E1: dout <= 8'b01010101; //  993 :  85 - 0x55
      11'h3E2: dout <= 8'b01010101; //  994 :  85 - 0x55
      11'h3E3: dout <= 8'b01010101; //  995 :  85 - 0x55
      11'h3E4: dout <= 8'b01010101; //  996 :  85 - 0x55
      11'h3E5: dout <= 8'b10010101; //  997 : 149 - 0x95
      11'h3E6: dout <= 8'b00000101; //  998 :   5 - 0x5
      11'h3E7: dout <= 8'b00000101; //  999 :   5 - 0x5
      11'h3E8: dout <= 8'b01010101; // 1000 :  85 - 0x55
      11'h3E9: dout <= 8'b01010101; // 1001 :  85 - 0x55
      11'h3EA: dout <= 8'b01010101; // 1002 :  85 - 0x55
      11'h3EB: dout <= 8'b01010101; // 1003 :  85 - 0x55
      11'h3EC: dout <= 8'b01010101; // 1004 :  85 - 0x55
      11'h3ED: dout <= 8'b00010001; // 1005 :  17 - 0x11
      11'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      11'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout <= 8'b01010101; // 1008 :  85 - 0x55
      11'h3F1: dout <= 8'b01010101; // 1009 :  85 - 0x55
      11'h3F2: dout <= 8'b01010101; // 1010 :  85 - 0x55
      11'h3F3: dout <= 8'b01010101; // 1011 :  85 - 0x55
      11'h3F4: dout <= 8'b01010101; // 1012 :  85 - 0x55
      11'h3F5: dout <= 8'b01010101; // 1013 :  85 - 0x55
      11'h3F6: dout <= 8'b01010101; // 1014 :  85 - 0x55
      11'h3F7: dout <= 8'b01010101; // 1015 :  85 - 0x55
      11'h3F8: dout <= 8'b01010101; // 1016 :  85 - 0x55
      11'h3F9: dout <= 8'b01010101; // 1017 :  85 - 0x55
      11'h3FA: dout <= 8'b01010101; // 1018 :  85 - 0x55
      11'h3FB: dout <= 8'b01010101; // 1019 :  85 - 0x55
      11'h3FC: dout <= 8'b01010101; // 1020 :  85 - 0x55
      11'h3FD: dout <= 8'b01010101; // 1021 :  85 - 0x55
      11'h3FE: dout <= 8'b01010101; // 1022 :  85 - 0x55
      11'h3FF: dout <= 8'b01010101; // 1023 :  85 - 0x55
     //----- Name Table 1---------
      11'h400: dout <= 8'b00100000; // 1024 :  32 - 0x20 -- line 0x0
      11'h401: dout <= 8'b00100000; // 1025 :  32 - 0x20
      11'h402: dout <= 8'b00100000; // 1026 :  32 - 0x20
      11'h403: dout <= 8'b00100000; // 1027 :  32 - 0x20
      11'h404: dout <= 8'b00100000; // 1028 :  32 - 0x20
      11'h405: dout <= 8'b00100000; // 1029 :  32 - 0x20
      11'h406: dout <= 8'b00100000; // 1030 :  32 - 0x20
      11'h407: dout <= 8'b00100000; // 1031 :  32 - 0x20
      11'h408: dout <= 8'b00100000; // 1032 :  32 - 0x20
      11'h409: dout <= 8'b00100000; // 1033 :  32 - 0x20
      11'h40A: dout <= 8'b00100000; // 1034 :  32 - 0x20
      11'h40B: dout <= 8'b00100000; // 1035 :  32 - 0x20
      11'h40C: dout <= 8'b00100000; // 1036 :  32 - 0x20
      11'h40D: dout <= 8'b00100000; // 1037 :  32 - 0x20
      11'h40E: dout <= 8'b00100000; // 1038 :  32 - 0x20
      11'h40F: dout <= 8'b00100000; // 1039 :  32 - 0x20
      11'h410: dout <= 8'b00100000; // 1040 :  32 - 0x20
      11'h411: dout <= 8'b00100000; // 1041 :  32 - 0x20
      11'h412: dout <= 8'b00100000; // 1042 :  32 - 0x20
      11'h413: dout <= 8'b00100000; // 1043 :  32 - 0x20
      11'h414: dout <= 8'b00100000; // 1044 :  32 - 0x20
      11'h415: dout <= 8'b00100000; // 1045 :  32 - 0x20
      11'h416: dout <= 8'b00100000; // 1046 :  32 - 0x20
      11'h417: dout <= 8'b00100000; // 1047 :  32 - 0x20
      11'h418: dout <= 8'b00100000; // 1048 :  32 - 0x20
      11'h419: dout <= 8'b00100000; // 1049 :  32 - 0x20
      11'h41A: dout <= 8'b00100000; // 1050 :  32 - 0x20
      11'h41B: dout <= 8'b00100000; // 1051 :  32 - 0x20
      11'h41C: dout <= 8'b00100000; // 1052 :  32 - 0x20
      11'h41D: dout <= 8'b00100000; // 1053 :  32 - 0x20
      11'h41E: dout <= 8'b00100000; // 1054 :  32 - 0x20
      11'h41F: dout <= 8'b00100000; // 1055 :  32 - 0x20
      11'h420: dout <= 8'b00100000; // 1056 :  32 - 0x20 -- line 0x1
      11'h421: dout <= 8'b00100000; // 1057 :  32 - 0x20
      11'h422: dout <= 8'b00100000; // 1058 :  32 - 0x20
      11'h423: dout <= 8'b00100000; // 1059 :  32 - 0x20
      11'h424: dout <= 8'b00100000; // 1060 :  32 - 0x20
      11'h425: dout <= 8'b00100000; // 1061 :  32 - 0x20
      11'h426: dout <= 8'b00100000; // 1062 :  32 - 0x20
      11'h427: dout <= 8'b00100000; // 1063 :  32 - 0x20
      11'h428: dout <= 8'b00100000; // 1064 :  32 - 0x20
      11'h429: dout <= 8'b00100000; // 1065 :  32 - 0x20
      11'h42A: dout <= 8'b00100000; // 1066 :  32 - 0x20
      11'h42B: dout <= 8'b00100000; // 1067 :  32 - 0x20
      11'h42C: dout <= 8'b00100000; // 1068 :  32 - 0x20
      11'h42D: dout <= 8'b00100000; // 1069 :  32 - 0x20
      11'h42E: dout <= 8'b00100000; // 1070 :  32 - 0x20
      11'h42F: dout <= 8'b00100000; // 1071 :  32 - 0x20
      11'h430: dout <= 8'b00100000; // 1072 :  32 - 0x20
      11'h431: dout <= 8'b00100000; // 1073 :  32 - 0x20
      11'h432: dout <= 8'b00100000; // 1074 :  32 - 0x20
      11'h433: dout <= 8'b00100000; // 1075 :  32 - 0x20
      11'h434: dout <= 8'b00100000; // 1076 :  32 - 0x20
      11'h435: dout <= 8'b00100000; // 1077 :  32 - 0x20
      11'h436: dout <= 8'b00100000; // 1078 :  32 - 0x20
      11'h437: dout <= 8'b00100000; // 1079 :  32 - 0x20
      11'h438: dout <= 8'b00100000; // 1080 :  32 - 0x20
      11'h439: dout <= 8'b00100000; // 1081 :  32 - 0x20
      11'h43A: dout <= 8'b00100000; // 1082 :  32 - 0x20
      11'h43B: dout <= 8'b00100000; // 1083 :  32 - 0x20
      11'h43C: dout <= 8'b00100000; // 1084 :  32 - 0x20
      11'h43D: dout <= 8'b00100000; // 1085 :  32 - 0x20
      11'h43E: dout <= 8'b00100000; // 1086 :  32 - 0x20
      11'h43F: dout <= 8'b00100000; // 1087 :  32 - 0x20
      11'h440: dout <= 8'b00100000; // 1088 :  32 - 0x20 -- line 0x2
      11'h441: dout <= 8'b00100000; // 1089 :  32 - 0x20
      11'h442: dout <= 8'b00100000; // 1090 :  32 - 0x20
      11'h443: dout <= 8'b00100000; // 1091 :  32 - 0x20
      11'h444: dout <= 8'b00100000; // 1092 :  32 - 0x20
      11'h445: dout <= 8'b00100000; // 1093 :  32 - 0x20
      11'h446: dout <= 8'b00100000; // 1094 :  32 - 0x20
      11'h447: dout <= 8'b00100000; // 1095 :  32 - 0x20
      11'h448: dout <= 8'b00100000; // 1096 :  32 - 0x20
      11'h449: dout <= 8'b00100000; // 1097 :  32 - 0x20
      11'h44A: dout <= 8'b00100000; // 1098 :  32 - 0x20
      11'h44B: dout <= 8'b00100000; // 1099 :  32 - 0x20
      11'h44C: dout <= 8'b00100000; // 1100 :  32 - 0x20
      11'h44D: dout <= 8'b00100000; // 1101 :  32 - 0x20
      11'h44E: dout <= 8'b00100000; // 1102 :  32 - 0x20
      11'h44F: dout <= 8'b00100000; // 1103 :  32 - 0x20
      11'h450: dout <= 8'b00100000; // 1104 :  32 - 0x20
      11'h451: dout <= 8'b00100000; // 1105 :  32 - 0x20
      11'h452: dout <= 8'b00100000; // 1106 :  32 - 0x20
      11'h453: dout <= 8'b00100000; // 1107 :  32 - 0x20
      11'h454: dout <= 8'b00100000; // 1108 :  32 - 0x20
      11'h455: dout <= 8'b00100000; // 1109 :  32 - 0x20
      11'h456: dout <= 8'b00100000; // 1110 :  32 - 0x20
      11'h457: dout <= 8'b00100000; // 1111 :  32 - 0x20
      11'h458: dout <= 8'b00100000; // 1112 :  32 - 0x20
      11'h459: dout <= 8'b00100000; // 1113 :  32 - 0x20
      11'h45A: dout <= 8'b00100000; // 1114 :  32 - 0x20
      11'h45B: dout <= 8'b00100000; // 1115 :  32 - 0x20
      11'h45C: dout <= 8'b00100000; // 1116 :  32 - 0x20
      11'h45D: dout <= 8'b00100000; // 1117 :  32 - 0x20
      11'h45E: dout <= 8'b00100000; // 1118 :  32 - 0x20
      11'h45F: dout <= 8'b00100000; // 1119 :  32 - 0x20
      11'h460: dout <= 8'b00100000; // 1120 :  32 - 0x20 -- line 0x3
      11'h461: dout <= 8'b00100000; // 1121 :  32 - 0x20
      11'h462: dout <= 8'b00100000; // 1122 :  32 - 0x20
      11'h463: dout <= 8'b00100000; // 1123 :  32 - 0x20
      11'h464: dout <= 8'b00100000; // 1124 :  32 - 0x20
      11'h465: dout <= 8'b00100000; // 1125 :  32 - 0x20
      11'h466: dout <= 8'b00100000; // 1126 :  32 - 0x20
      11'h467: dout <= 8'b00100000; // 1127 :  32 - 0x20
      11'h468: dout <= 8'b00100000; // 1128 :  32 - 0x20
      11'h469: dout <= 8'b00100000; // 1129 :  32 - 0x20
      11'h46A: dout <= 8'b00100000; // 1130 :  32 - 0x20
      11'h46B: dout <= 8'b00100000; // 1131 :  32 - 0x20
      11'h46C: dout <= 8'b00100000; // 1132 :  32 - 0x20
      11'h46D: dout <= 8'b00100000; // 1133 :  32 - 0x20
      11'h46E: dout <= 8'b00100000; // 1134 :  32 - 0x20
      11'h46F: dout <= 8'b00100000; // 1135 :  32 - 0x20
      11'h470: dout <= 8'b00100000; // 1136 :  32 - 0x20
      11'h471: dout <= 8'b00100000; // 1137 :  32 - 0x20
      11'h472: dout <= 8'b00100000; // 1138 :  32 - 0x20
      11'h473: dout <= 8'b00100000; // 1139 :  32 - 0x20
      11'h474: dout <= 8'b00100000; // 1140 :  32 - 0x20
      11'h475: dout <= 8'b00100000; // 1141 :  32 - 0x20
      11'h476: dout <= 8'b00100000; // 1142 :  32 - 0x20
      11'h477: dout <= 8'b00100000; // 1143 :  32 - 0x20
      11'h478: dout <= 8'b00100000; // 1144 :  32 - 0x20
      11'h479: dout <= 8'b00100000; // 1145 :  32 - 0x20
      11'h47A: dout <= 8'b00100000; // 1146 :  32 - 0x20
      11'h47B: dout <= 8'b00100000; // 1147 :  32 - 0x20
      11'h47C: dout <= 8'b00100000; // 1148 :  32 - 0x20
      11'h47D: dout <= 8'b00100000; // 1149 :  32 - 0x20
      11'h47E: dout <= 8'b00100000; // 1150 :  32 - 0x20
      11'h47F: dout <= 8'b00100000; // 1151 :  32 - 0x20
      11'h480: dout <= 8'b00100000; // 1152 :  32 - 0x20 -- line 0x4
      11'h481: dout <= 8'b00100000; // 1153 :  32 - 0x20
      11'h482: dout <= 8'b00100000; // 1154 :  32 - 0x20
      11'h483: dout <= 8'b00100000; // 1155 :  32 - 0x20
      11'h484: dout <= 8'b00100000; // 1156 :  32 - 0x20
      11'h485: dout <= 8'b00100000; // 1157 :  32 - 0x20
      11'h486: dout <= 8'b00100000; // 1158 :  32 - 0x20
      11'h487: dout <= 8'b00100000; // 1159 :  32 - 0x20
      11'h488: dout <= 8'b00100000; // 1160 :  32 - 0x20
      11'h489: dout <= 8'b00100000; // 1161 :  32 - 0x20
      11'h48A: dout <= 8'b00100000; // 1162 :  32 - 0x20
      11'h48B: dout <= 8'b00100000; // 1163 :  32 - 0x20
      11'h48C: dout <= 8'b00100000; // 1164 :  32 - 0x20
      11'h48D: dout <= 8'b00100000; // 1165 :  32 - 0x20
      11'h48E: dout <= 8'b00100000; // 1166 :  32 - 0x20
      11'h48F: dout <= 8'b00100000; // 1167 :  32 - 0x20
      11'h490: dout <= 8'b00100000; // 1168 :  32 - 0x20
      11'h491: dout <= 8'b00100000; // 1169 :  32 - 0x20
      11'h492: dout <= 8'b00100000; // 1170 :  32 - 0x20
      11'h493: dout <= 8'b00100000; // 1171 :  32 - 0x20
      11'h494: dout <= 8'b00100000; // 1172 :  32 - 0x20
      11'h495: dout <= 8'b00100000; // 1173 :  32 - 0x20
      11'h496: dout <= 8'b00100000; // 1174 :  32 - 0x20
      11'h497: dout <= 8'b00100000; // 1175 :  32 - 0x20
      11'h498: dout <= 8'b00100000; // 1176 :  32 - 0x20
      11'h499: dout <= 8'b00100000; // 1177 :  32 - 0x20
      11'h49A: dout <= 8'b00100000; // 1178 :  32 - 0x20
      11'h49B: dout <= 8'b00100000; // 1179 :  32 - 0x20
      11'h49C: dout <= 8'b00100000; // 1180 :  32 - 0x20
      11'h49D: dout <= 8'b00100000; // 1181 :  32 - 0x20
      11'h49E: dout <= 8'b00100000; // 1182 :  32 - 0x20
      11'h49F: dout <= 8'b00100000; // 1183 :  32 - 0x20
      11'h4A0: dout <= 8'b00100000; // 1184 :  32 - 0x20 -- line 0x5
      11'h4A1: dout <= 8'b00100000; // 1185 :  32 - 0x20
      11'h4A2: dout <= 8'b00100000; // 1186 :  32 - 0x20
      11'h4A3: dout <= 8'b00100000; // 1187 :  32 - 0x20
      11'h4A4: dout <= 8'b00100000; // 1188 :  32 - 0x20
      11'h4A5: dout <= 8'b00100000; // 1189 :  32 - 0x20
      11'h4A6: dout <= 8'b00100000; // 1190 :  32 - 0x20
      11'h4A7: dout <= 8'b00100000; // 1191 :  32 - 0x20
      11'h4A8: dout <= 8'b00100000; // 1192 :  32 - 0x20
      11'h4A9: dout <= 8'b00100000; // 1193 :  32 - 0x20
      11'h4AA: dout <= 8'b00100000; // 1194 :  32 - 0x20
      11'h4AB: dout <= 8'b00100000; // 1195 :  32 - 0x20
      11'h4AC: dout <= 8'b00100000; // 1196 :  32 - 0x20
      11'h4AD: dout <= 8'b00100000; // 1197 :  32 - 0x20
      11'h4AE: dout <= 8'b00100000; // 1198 :  32 - 0x20
      11'h4AF: dout <= 8'b00100000; // 1199 :  32 - 0x20
      11'h4B0: dout <= 8'b00100000; // 1200 :  32 - 0x20
      11'h4B1: dout <= 8'b00100000; // 1201 :  32 - 0x20
      11'h4B2: dout <= 8'b00100000; // 1202 :  32 - 0x20
      11'h4B3: dout <= 8'b00100000; // 1203 :  32 - 0x20
      11'h4B4: dout <= 8'b00100000; // 1204 :  32 - 0x20
      11'h4B5: dout <= 8'b00100000; // 1205 :  32 - 0x20
      11'h4B6: dout <= 8'b00100000; // 1206 :  32 - 0x20
      11'h4B7: dout <= 8'b00100000; // 1207 :  32 - 0x20
      11'h4B8: dout <= 8'b00100000; // 1208 :  32 - 0x20
      11'h4B9: dout <= 8'b00100000; // 1209 :  32 - 0x20
      11'h4BA: dout <= 8'b00100000; // 1210 :  32 - 0x20
      11'h4BB: dout <= 8'b00100000; // 1211 :  32 - 0x20
      11'h4BC: dout <= 8'b00100000; // 1212 :  32 - 0x20
      11'h4BD: dout <= 8'b00100000; // 1213 :  32 - 0x20
      11'h4BE: dout <= 8'b00100000; // 1214 :  32 - 0x20
      11'h4BF: dout <= 8'b00100000; // 1215 :  32 - 0x20
      11'h4C0: dout <= 8'b00100000; // 1216 :  32 - 0x20 -- line 0x6
      11'h4C1: dout <= 8'b00100000; // 1217 :  32 - 0x20
      11'h4C2: dout <= 8'b00100000; // 1218 :  32 - 0x20
      11'h4C3: dout <= 8'b00100000; // 1219 :  32 - 0x20
      11'h4C4: dout <= 8'b00100000; // 1220 :  32 - 0x20
      11'h4C5: dout <= 8'b00100000; // 1221 :  32 - 0x20
      11'h4C6: dout <= 8'b00100000; // 1222 :  32 - 0x20
      11'h4C7: dout <= 8'b00100000; // 1223 :  32 - 0x20
      11'h4C8: dout <= 8'b00100000; // 1224 :  32 - 0x20
      11'h4C9: dout <= 8'b00100000; // 1225 :  32 - 0x20
      11'h4CA: dout <= 8'b00100000; // 1226 :  32 - 0x20
      11'h4CB: dout <= 8'b00100000; // 1227 :  32 - 0x20
      11'h4CC: dout <= 8'b00100000; // 1228 :  32 - 0x20
      11'h4CD: dout <= 8'b00100000; // 1229 :  32 - 0x20
      11'h4CE: dout <= 8'b00100000; // 1230 :  32 - 0x20
      11'h4CF: dout <= 8'b00100000; // 1231 :  32 - 0x20
      11'h4D0: dout <= 8'b00100000; // 1232 :  32 - 0x20
      11'h4D1: dout <= 8'b00100000; // 1233 :  32 - 0x20
      11'h4D2: dout <= 8'b00100000; // 1234 :  32 - 0x20
      11'h4D3: dout <= 8'b00100000; // 1235 :  32 - 0x20
      11'h4D4: dout <= 8'b00100000; // 1236 :  32 - 0x20
      11'h4D5: dout <= 8'b00100000; // 1237 :  32 - 0x20
      11'h4D6: dout <= 8'b00100000; // 1238 :  32 - 0x20
      11'h4D7: dout <= 8'b00100000; // 1239 :  32 - 0x20
      11'h4D8: dout <= 8'b00100000; // 1240 :  32 - 0x20
      11'h4D9: dout <= 8'b00100000; // 1241 :  32 - 0x20
      11'h4DA: dout <= 8'b00100000; // 1242 :  32 - 0x20
      11'h4DB: dout <= 8'b00100000; // 1243 :  32 - 0x20
      11'h4DC: dout <= 8'b00100000; // 1244 :  32 - 0x20
      11'h4DD: dout <= 8'b00100000; // 1245 :  32 - 0x20
      11'h4DE: dout <= 8'b00100000; // 1246 :  32 - 0x20
      11'h4DF: dout <= 8'b00100000; // 1247 :  32 - 0x20
      11'h4E0: dout <= 8'b00100000; // 1248 :  32 - 0x20 -- line 0x7
      11'h4E1: dout <= 8'b00100000; // 1249 :  32 - 0x20
      11'h4E2: dout <= 8'b00100000; // 1250 :  32 - 0x20
      11'h4E3: dout <= 8'b00100000; // 1251 :  32 - 0x20
      11'h4E4: dout <= 8'b00100000; // 1252 :  32 - 0x20
      11'h4E5: dout <= 8'b00100000; // 1253 :  32 - 0x20
      11'h4E6: dout <= 8'b00100000; // 1254 :  32 - 0x20
      11'h4E7: dout <= 8'b00100000; // 1255 :  32 - 0x20
      11'h4E8: dout <= 8'b00100000; // 1256 :  32 - 0x20
      11'h4E9: dout <= 8'b00100000; // 1257 :  32 - 0x20
      11'h4EA: dout <= 8'b00100000; // 1258 :  32 - 0x20
      11'h4EB: dout <= 8'b00100000; // 1259 :  32 - 0x20
      11'h4EC: dout <= 8'b00100000; // 1260 :  32 - 0x20
      11'h4ED: dout <= 8'b00100000; // 1261 :  32 - 0x20
      11'h4EE: dout <= 8'b00100000; // 1262 :  32 - 0x20
      11'h4EF: dout <= 8'b00100000; // 1263 :  32 - 0x20
      11'h4F0: dout <= 8'b00100000; // 1264 :  32 - 0x20
      11'h4F1: dout <= 8'b00100000; // 1265 :  32 - 0x20
      11'h4F2: dout <= 8'b00100000; // 1266 :  32 - 0x20
      11'h4F3: dout <= 8'b00100000; // 1267 :  32 - 0x20
      11'h4F4: dout <= 8'b00100000; // 1268 :  32 - 0x20
      11'h4F5: dout <= 8'b00100000; // 1269 :  32 - 0x20
      11'h4F6: dout <= 8'b00100000; // 1270 :  32 - 0x20
      11'h4F7: dout <= 8'b00100000; // 1271 :  32 - 0x20
      11'h4F8: dout <= 8'b00100000; // 1272 :  32 - 0x20
      11'h4F9: dout <= 8'b00100000; // 1273 :  32 - 0x20
      11'h4FA: dout <= 8'b00100000; // 1274 :  32 - 0x20
      11'h4FB: dout <= 8'b00100000; // 1275 :  32 - 0x20
      11'h4FC: dout <= 8'b00100000; // 1276 :  32 - 0x20
      11'h4FD: dout <= 8'b00100000; // 1277 :  32 - 0x20
      11'h4FE: dout <= 8'b00100000; // 1278 :  32 - 0x20
      11'h4FF: dout <= 8'b00100000; // 1279 :  32 - 0x20
      11'h500: dout <= 8'b00100000; // 1280 :  32 - 0x20 -- line 0x8
      11'h501: dout <= 8'b00100000; // 1281 :  32 - 0x20
      11'h502: dout <= 8'b00100000; // 1282 :  32 - 0x20
      11'h503: dout <= 8'b00100000; // 1283 :  32 - 0x20
      11'h504: dout <= 8'b00100000; // 1284 :  32 - 0x20
      11'h505: dout <= 8'b00100000; // 1285 :  32 - 0x20
      11'h506: dout <= 8'b00100000; // 1286 :  32 - 0x20
      11'h507: dout <= 8'b00100000; // 1287 :  32 - 0x20
      11'h508: dout <= 8'b00100000; // 1288 :  32 - 0x20
      11'h509: dout <= 8'b00100000; // 1289 :  32 - 0x20
      11'h50A: dout <= 8'b00100000; // 1290 :  32 - 0x20
      11'h50B: dout <= 8'b00100000; // 1291 :  32 - 0x20
      11'h50C: dout <= 8'b00100000; // 1292 :  32 - 0x20
      11'h50D: dout <= 8'b00100000; // 1293 :  32 - 0x20
      11'h50E: dout <= 8'b00100000; // 1294 :  32 - 0x20
      11'h50F: dout <= 8'b00100000; // 1295 :  32 - 0x20
      11'h510: dout <= 8'b00100000; // 1296 :  32 - 0x20
      11'h511: dout <= 8'b00100000; // 1297 :  32 - 0x20
      11'h512: dout <= 8'b00100000; // 1298 :  32 - 0x20
      11'h513: dout <= 8'b00100000; // 1299 :  32 - 0x20
      11'h514: dout <= 8'b00100000; // 1300 :  32 - 0x20
      11'h515: dout <= 8'b00100000; // 1301 :  32 - 0x20
      11'h516: dout <= 8'b00100000; // 1302 :  32 - 0x20
      11'h517: dout <= 8'b00100000; // 1303 :  32 - 0x20
      11'h518: dout <= 8'b00100000; // 1304 :  32 - 0x20
      11'h519: dout <= 8'b00100000; // 1305 :  32 - 0x20
      11'h51A: dout <= 8'b00100000; // 1306 :  32 - 0x20
      11'h51B: dout <= 8'b00100000; // 1307 :  32 - 0x20
      11'h51C: dout <= 8'b00100000; // 1308 :  32 - 0x20
      11'h51D: dout <= 8'b00100000; // 1309 :  32 - 0x20
      11'h51E: dout <= 8'b00100000; // 1310 :  32 - 0x20
      11'h51F: dout <= 8'b00100000; // 1311 :  32 - 0x20
      11'h520: dout <= 8'b00100000; // 1312 :  32 - 0x20 -- line 0x9
      11'h521: dout <= 8'b00100000; // 1313 :  32 - 0x20
      11'h522: dout <= 8'b00100000; // 1314 :  32 - 0x20
      11'h523: dout <= 8'b00100000; // 1315 :  32 - 0x20
      11'h524: dout <= 8'b00100000; // 1316 :  32 - 0x20
      11'h525: dout <= 8'b00100000; // 1317 :  32 - 0x20
      11'h526: dout <= 8'b00100000; // 1318 :  32 - 0x20
      11'h527: dout <= 8'b00100000; // 1319 :  32 - 0x20
      11'h528: dout <= 8'b00100000; // 1320 :  32 - 0x20
      11'h529: dout <= 8'b00100000; // 1321 :  32 - 0x20
      11'h52A: dout <= 8'b00100000; // 1322 :  32 - 0x20
      11'h52B: dout <= 8'b00100000; // 1323 :  32 - 0x20
      11'h52C: dout <= 8'b00100000; // 1324 :  32 - 0x20
      11'h52D: dout <= 8'b00100000; // 1325 :  32 - 0x20
      11'h52E: dout <= 8'b00100000; // 1326 :  32 - 0x20
      11'h52F: dout <= 8'b00100000; // 1327 :  32 - 0x20
      11'h530: dout <= 8'b00100000; // 1328 :  32 - 0x20
      11'h531: dout <= 8'b00100000; // 1329 :  32 - 0x20
      11'h532: dout <= 8'b00100000; // 1330 :  32 - 0x20
      11'h533: dout <= 8'b00100000; // 1331 :  32 - 0x20
      11'h534: dout <= 8'b00100000; // 1332 :  32 - 0x20
      11'h535: dout <= 8'b00100000; // 1333 :  32 - 0x20
      11'h536: dout <= 8'b00100000; // 1334 :  32 - 0x20
      11'h537: dout <= 8'b00100000; // 1335 :  32 - 0x20
      11'h538: dout <= 8'b00100000; // 1336 :  32 - 0x20
      11'h539: dout <= 8'b00100000; // 1337 :  32 - 0x20
      11'h53A: dout <= 8'b00100000; // 1338 :  32 - 0x20
      11'h53B: dout <= 8'b00100000; // 1339 :  32 - 0x20
      11'h53C: dout <= 8'b00100000; // 1340 :  32 - 0x20
      11'h53D: dout <= 8'b00100000; // 1341 :  32 - 0x20
      11'h53E: dout <= 8'b00100000; // 1342 :  32 - 0x20
      11'h53F: dout <= 8'b00100000; // 1343 :  32 - 0x20
      11'h540: dout <= 8'b00100000; // 1344 :  32 - 0x20 -- line 0xa
      11'h541: dout <= 8'b00100000; // 1345 :  32 - 0x20
      11'h542: dout <= 8'b00100000; // 1346 :  32 - 0x20
      11'h543: dout <= 8'b00100000; // 1347 :  32 - 0x20
      11'h544: dout <= 8'b00100000; // 1348 :  32 - 0x20
      11'h545: dout <= 8'b00100000; // 1349 :  32 - 0x20
      11'h546: dout <= 8'b00100000; // 1350 :  32 - 0x20
      11'h547: dout <= 8'b00100000; // 1351 :  32 - 0x20
      11'h548: dout <= 8'b00100000; // 1352 :  32 - 0x20
      11'h549: dout <= 8'b00100000; // 1353 :  32 - 0x20
      11'h54A: dout <= 8'b00100000; // 1354 :  32 - 0x20
      11'h54B: dout <= 8'b00100000; // 1355 :  32 - 0x20
      11'h54C: dout <= 8'b00100000; // 1356 :  32 - 0x20
      11'h54D: dout <= 8'b00100000; // 1357 :  32 - 0x20
      11'h54E: dout <= 8'b00100000; // 1358 :  32 - 0x20
      11'h54F: dout <= 8'b00100000; // 1359 :  32 - 0x20
      11'h550: dout <= 8'b00100000; // 1360 :  32 - 0x20
      11'h551: dout <= 8'b00100000; // 1361 :  32 - 0x20
      11'h552: dout <= 8'b00100000; // 1362 :  32 - 0x20
      11'h553: dout <= 8'b00100000; // 1363 :  32 - 0x20
      11'h554: dout <= 8'b00100000; // 1364 :  32 - 0x20
      11'h555: dout <= 8'b00100000; // 1365 :  32 - 0x20
      11'h556: dout <= 8'b00100000; // 1366 :  32 - 0x20
      11'h557: dout <= 8'b00100000; // 1367 :  32 - 0x20
      11'h558: dout <= 8'b00100000; // 1368 :  32 - 0x20
      11'h559: dout <= 8'b00100000; // 1369 :  32 - 0x20
      11'h55A: dout <= 8'b00100000; // 1370 :  32 - 0x20
      11'h55B: dout <= 8'b00100000; // 1371 :  32 - 0x20
      11'h55C: dout <= 8'b00100000; // 1372 :  32 - 0x20
      11'h55D: dout <= 8'b00100000; // 1373 :  32 - 0x20
      11'h55E: dout <= 8'b00100000; // 1374 :  32 - 0x20
      11'h55F: dout <= 8'b00100000; // 1375 :  32 - 0x20
      11'h560: dout <= 8'b00100000; // 1376 :  32 - 0x20 -- line 0xb
      11'h561: dout <= 8'b00100000; // 1377 :  32 - 0x20
      11'h562: dout <= 8'b00100000; // 1378 :  32 - 0x20
      11'h563: dout <= 8'b00100000; // 1379 :  32 - 0x20
      11'h564: dout <= 8'b00100000; // 1380 :  32 - 0x20
      11'h565: dout <= 8'b00100000; // 1381 :  32 - 0x20
      11'h566: dout <= 8'b00100000; // 1382 :  32 - 0x20
      11'h567: dout <= 8'b00100000; // 1383 :  32 - 0x20
      11'h568: dout <= 8'b00100000; // 1384 :  32 - 0x20
      11'h569: dout <= 8'b00100000; // 1385 :  32 - 0x20
      11'h56A: dout <= 8'b00100000; // 1386 :  32 - 0x20
      11'h56B: dout <= 8'b00100000; // 1387 :  32 - 0x20
      11'h56C: dout <= 8'b00100000; // 1388 :  32 - 0x20
      11'h56D: dout <= 8'b00100000; // 1389 :  32 - 0x20
      11'h56E: dout <= 8'b00100000; // 1390 :  32 - 0x20
      11'h56F: dout <= 8'b00100000; // 1391 :  32 - 0x20
      11'h570: dout <= 8'b00100000; // 1392 :  32 - 0x20
      11'h571: dout <= 8'b00100000; // 1393 :  32 - 0x20
      11'h572: dout <= 8'b00100000; // 1394 :  32 - 0x20
      11'h573: dout <= 8'b00100000; // 1395 :  32 - 0x20
      11'h574: dout <= 8'b00100000; // 1396 :  32 - 0x20
      11'h575: dout <= 8'b00100000; // 1397 :  32 - 0x20
      11'h576: dout <= 8'b00100000; // 1398 :  32 - 0x20
      11'h577: dout <= 8'b00100000; // 1399 :  32 - 0x20
      11'h578: dout <= 8'b00100000; // 1400 :  32 - 0x20
      11'h579: dout <= 8'b00100000; // 1401 :  32 - 0x20
      11'h57A: dout <= 8'b00100000; // 1402 :  32 - 0x20
      11'h57B: dout <= 8'b00100000; // 1403 :  32 - 0x20
      11'h57C: dout <= 8'b00100000; // 1404 :  32 - 0x20
      11'h57D: dout <= 8'b00100000; // 1405 :  32 - 0x20
      11'h57E: dout <= 8'b00100000; // 1406 :  32 - 0x20
      11'h57F: dout <= 8'b00100000; // 1407 :  32 - 0x20
      11'h580: dout <= 8'b00100000; // 1408 :  32 - 0x20 -- line 0xc
      11'h581: dout <= 8'b00100000; // 1409 :  32 - 0x20
      11'h582: dout <= 8'b00100000; // 1410 :  32 - 0x20
      11'h583: dout <= 8'b00100000; // 1411 :  32 - 0x20
      11'h584: dout <= 8'b00100000; // 1412 :  32 - 0x20
      11'h585: dout <= 8'b00100000; // 1413 :  32 - 0x20
      11'h586: dout <= 8'b00100000; // 1414 :  32 - 0x20
      11'h587: dout <= 8'b00100000; // 1415 :  32 - 0x20
      11'h588: dout <= 8'b00100000; // 1416 :  32 - 0x20
      11'h589: dout <= 8'b00100000; // 1417 :  32 - 0x20
      11'h58A: dout <= 8'b00100000; // 1418 :  32 - 0x20
      11'h58B: dout <= 8'b00100000; // 1419 :  32 - 0x20
      11'h58C: dout <= 8'b00100000; // 1420 :  32 - 0x20
      11'h58D: dout <= 8'b00100000; // 1421 :  32 - 0x20
      11'h58E: dout <= 8'b00100000; // 1422 :  32 - 0x20
      11'h58F: dout <= 8'b00100000; // 1423 :  32 - 0x20
      11'h590: dout <= 8'b00100000; // 1424 :  32 - 0x20
      11'h591: dout <= 8'b00100000; // 1425 :  32 - 0x20
      11'h592: dout <= 8'b00100000; // 1426 :  32 - 0x20
      11'h593: dout <= 8'b00100000; // 1427 :  32 - 0x20
      11'h594: dout <= 8'b00100000; // 1428 :  32 - 0x20
      11'h595: dout <= 8'b00100000; // 1429 :  32 - 0x20
      11'h596: dout <= 8'b00100000; // 1430 :  32 - 0x20
      11'h597: dout <= 8'b00100000; // 1431 :  32 - 0x20
      11'h598: dout <= 8'b00100000; // 1432 :  32 - 0x20
      11'h599: dout <= 8'b00100000; // 1433 :  32 - 0x20
      11'h59A: dout <= 8'b00100000; // 1434 :  32 - 0x20
      11'h59B: dout <= 8'b00100000; // 1435 :  32 - 0x20
      11'h59C: dout <= 8'b00100000; // 1436 :  32 - 0x20
      11'h59D: dout <= 8'b00100000; // 1437 :  32 - 0x20
      11'h59E: dout <= 8'b00100000; // 1438 :  32 - 0x20
      11'h59F: dout <= 8'b00100000; // 1439 :  32 - 0x20
      11'h5A0: dout <= 8'b00100000; // 1440 :  32 - 0x20 -- line 0xd
      11'h5A1: dout <= 8'b00100000; // 1441 :  32 - 0x20
      11'h5A2: dout <= 8'b00100000; // 1442 :  32 - 0x20
      11'h5A3: dout <= 8'b00100000; // 1443 :  32 - 0x20
      11'h5A4: dout <= 8'b00100000; // 1444 :  32 - 0x20
      11'h5A5: dout <= 8'b00100000; // 1445 :  32 - 0x20
      11'h5A6: dout <= 8'b00100000; // 1446 :  32 - 0x20
      11'h5A7: dout <= 8'b00100000; // 1447 :  32 - 0x20
      11'h5A8: dout <= 8'b00100000; // 1448 :  32 - 0x20
      11'h5A9: dout <= 8'b00100000; // 1449 :  32 - 0x20
      11'h5AA: dout <= 8'b00100000; // 1450 :  32 - 0x20
      11'h5AB: dout <= 8'b00100000; // 1451 :  32 - 0x20
      11'h5AC: dout <= 8'b00100000; // 1452 :  32 - 0x20
      11'h5AD: dout <= 8'b00100000; // 1453 :  32 - 0x20
      11'h5AE: dout <= 8'b00100000; // 1454 :  32 - 0x20
      11'h5AF: dout <= 8'b00100000; // 1455 :  32 - 0x20
      11'h5B0: dout <= 8'b00100000; // 1456 :  32 - 0x20
      11'h5B1: dout <= 8'b00100000; // 1457 :  32 - 0x20
      11'h5B2: dout <= 8'b00100000; // 1458 :  32 - 0x20
      11'h5B3: dout <= 8'b00100000; // 1459 :  32 - 0x20
      11'h5B4: dout <= 8'b00100000; // 1460 :  32 - 0x20
      11'h5B5: dout <= 8'b00100000; // 1461 :  32 - 0x20
      11'h5B6: dout <= 8'b00100000; // 1462 :  32 - 0x20
      11'h5B7: dout <= 8'b00100000; // 1463 :  32 - 0x20
      11'h5B8: dout <= 8'b00100000; // 1464 :  32 - 0x20
      11'h5B9: dout <= 8'b00100000; // 1465 :  32 - 0x20
      11'h5BA: dout <= 8'b00100000; // 1466 :  32 - 0x20
      11'h5BB: dout <= 8'b00100000; // 1467 :  32 - 0x20
      11'h5BC: dout <= 8'b00100000; // 1468 :  32 - 0x20
      11'h5BD: dout <= 8'b00100000; // 1469 :  32 - 0x20
      11'h5BE: dout <= 8'b00100000; // 1470 :  32 - 0x20
      11'h5BF: dout <= 8'b00100000; // 1471 :  32 - 0x20
      11'h5C0: dout <= 8'b00100000; // 1472 :  32 - 0x20 -- line 0xe
      11'h5C1: dout <= 8'b00100000; // 1473 :  32 - 0x20
      11'h5C2: dout <= 8'b00100000; // 1474 :  32 - 0x20
      11'h5C3: dout <= 8'b00100000; // 1475 :  32 - 0x20
      11'h5C4: dout <= 8'b00100000; // 1476 :  32 - 0x20
      11'h5C5: dout <= 8'b00100000; // 1477 :  32 - 0x20
      11'h5C6: dout <= 8'b00100000; // 1478 :  32 - 0x20
      11'h5C7: dout <= 8'b00100000; // 1479 :  32 - 0x20
      11'h5C8: dout <= 8'b00100000; // 1480 :  32 - 0x20
      11'h5C9: dout <= 8'b00100000; // 1481 :  32 - 0x20
      11'h5CA: dout <= 8'b00100000; // 1482 :  32 - 0x20
      11'h5CB: dout <= 8'b00100000; // 1483 :  32 - 0x20
      11'h5CC: dout <= 8'b00100000; // 1484 :  32 - 0x20
      11'h5CD: dout <= 8'b00100000; // 1485 :  32 - 0x20
      11'h5CE: dout <= 8'b00100000; // 1486 :  32 - 0x20
      11'h5CF: dout <= 8'b00100000; // 1487 :  32 - 0x20
      11'h5D0: dout <= 8'b00100000; // 1488 :  32 - 0x20
      11'h5D1: dout <= 8'b00100000; // 1489 :  32 - 0x20
      11'h5D2: dout <= 8'b00100000; // 1490 :  32 - 0x20
      11'h5D3: dout <= 8'b00100000; // 1491 :  32 - 0x20
      11'h5D4: dout <= 8'b00100000; // 1492 :  32 - 0x20
      11'h5D5: dout <= 8'b00100000; // 1493 :  32 - 0x20
      11'h5D6: dout <= 8'b00100000; // 1494 :  32 - 0x20
      11'h5D7: dout <= 8'b00100000; // 1495 :  32 - 0x20
      11'h5D8: dout <= 8'b00100000; // 1496 :  32 - 0x20
      11'h5D9: dout <= 8'b00100000; // 1497 :  32 - 0x20
      11'h5DA: dout <= 8'b00100000; // 1498 :  32 - 0x20
      11'h5DB: dout <= 8'b00100000; // 1499 :  32 - 0x20
      11'h5DC: dout <= 8'b00100000; // 1500 :  32 - 0x20
      11'h5DD: dout <= 8'b00100000; // 1501 :  32 - 0x20
      11'h5DE: dout <= 8'b00100000; // 1502 :  32 - 0x20
      11'h5DF: dout <= 8'b00100000; // 1503 :  32 - 0x20
      11'h5E0: dout <= 8'b00100000; // 1504 :  32 - 0x20 -- line 0xf
      11'h5E1: dout <= 8'b00100000; // 1505 :  32 - 0x20
      11'h5E2: dout <= 8'b00100000; // 1506 :  32 - 0x20
      11'h5E3: dout <= 8'b00100000; // 1507 :  32 - 0x20
      11'h5E4: dout <= 8'b00100000; // 1508 :  32 - 0x20
      11'h5E5: dout <= 8'b00100000; // 1509 :  32 - 0x20
      11'h5E6: dout <= 8'b00100000; // 1510 :  32 - 0x20
      11'h5E7: dout <= 8'b00100000; // 1511 :  32 - 0x20
      11'h5E8: dout <= 8'b00100000; // 1512 :  32 - 0x20
      11'h5E9: dout <= 8'b00100000; // 1513 :  32 - 0x20
      11'h5EA: dout <= 8'b00100000; // 1514 :  32 - 0x20
      11'h5EB: dout <= 8'b00100000; // 1515 :  32 - 0x20
      11'h5EC: dout <= 8'b00100000; // 1516 :  32 - 0x20
      11'h5ED: dout <= 8'b00100000; // 1517 :  32 - 0x20
      11'h5EE: dout <= 8'b00100000; // 1518 :  32 - 0x20
      11'h5EF: dout <= 8'b00100000; // 1519 :  32 - 0x20
      11'h5F0: dout <= 8'b00100000; // 1520 :  32 - 0x20
      11'h5F1: dout <= 8'b00100000; // 1521 :  32 - 0x20
      11'h5F2: dout <= 8'b00100000; // 1522 :  32 - 0x20
      11'h5F3: dout <= 8'b00100000; // 1523 :  32 - 0x20
      11'h5F4: dout <= 8'b00100000; // 1524 :  32 - 0x20
      11'h5F5: dout <= 8'b00100000; // 1525 :  32 - 0x20
      11'h5F6: dout <= 8'b00100000; // 1526 :  32 - 0x20
      11'h5F7: dout <= 8'b00100000; // 1527 :  32 - 0x20
      11'h5F8: dout <= 8'b00100000; // 1528 :  32 - 0x20
      11'h5F9: dout <= 8'b00100000; // 1529 :  32 - 0x20
      11'h5FA: dout <= 8'b00100000; // 1530 :  32 - 0x20
      11'h5FB: dout <= 8'b00100000; // 1531 :  32 - 0x20
      11'h5FC: dout <= 8'b00100000; // 1532 :  32 - 0x20
      11'h5FD: dout <= 8'b00100000; // 1533 :  32 - 0x20
      11'h5FE: dout <= 8'b00100000; // 1534 :  32 - 0x20
      11'h5FF: dout <= 8'b00100000; // 1535 :  32 - 0x20
      11'h600: dout <= 8'b00100000; // 1536 :  32 - 0x20 -- line 0x10
      11'h601: dout <= 8'b00100000; // 1537 :  32 - 0x20
      11'h602: dout <= 8'b00100000; // 1538 :  32 - 0x20
      11'h603: dout <= 8'b00100000; // 1539 :  32 - 0x20
      11'h604: dout <= 8'b00100000; // 1540 :  32 - 0x20
      11'h605: dout <= 8'b00100000; // 1541 :  32 - 0x20
      11'h606: dout <= 8'b00100000; // 1542 :  32 - 0x20
      11'h607: dout <= 8'b00100000; // 1543 :  32 - 0x20
      11'h608: dout <= 8'b00100000; // 1544 :  32 - 0x20
      11'h609: dout <= 8'b00100000; // 1545 :  32 - 0x20
      11'h60A: dout <= 8'b00100000; // 1546 :  32 - 0x20
      11'h60B: dout <= 8'b00100000; // 1547 :  32 - 0x20
      11'h60C: dout <= 8'b00100000; // 1548 :  32 - 0x20
      11'h60D: dout <= 8'b00100000; // 1549 :  32 - 0x20
      11'h60E: dout <= 8'b00100000; // 1550 :  32 - 0x20
      11'h60F: dout <= 8'b00100000; // 1551 :  32 - 0x20
      11'h610: dout <= 8'b00100000; // 1552 :  32 - 0x20
      11'h611: dout <= 8'b00100000; // 1553 :  32 - 0x20
      11'h612: dout <= 8'b00100000; // 1554 :  32 - 0x20
      11'h613: dout <= 8'b00100000; // 1555 :  32 - 0x20
      11'h614: dout <= 8'b00100000; // 1556 :  32 - 0x20
      11'h615: dout <= 8'b00100000; // 1557 :  32 - 0x20
      11'h616: dout <= 8'b00100000; // 1558 :  32 - 0x20
      11'h617: dout <= 8'b00100000; // 1559 :  32 - 0x20
      11'h618: dout <= 8'b00100000; // 1560 :  32 - 0x20
      11'h619: dout <= 8'b00100000; // 1561 :  32 - 0x20
      11'h61A: dout <= 8'b00100000; // 1562 :  32 - 0x20
      11'h61B: dout <= 8'b00100000; // 1563 :  32 - 0x20
      11'h61C: dout <= 8'b00100000; // 1564 :  32 - 0x20
      11'h61D: dout <= 8'b00100000; // 1565 :  32 - 0x20
      11'h61E: dout <= 8'b00100000; // 1566 :  32 - 0x20
      11'h61F: dout <= 8'b00100000; // 1567 :  32 - 0x20
      11'h620: dout <= 8'b00100000; // 1568 :  32 - 0x20 -- line 0x11
      11'h621: dout <= 8'b00100000; // 1569 :  32 - 0x20
      11'h622: dout <= 8'b00100000; // 1570 :  32 - 0x20
      11'h623: dout <= 8'b00100000; // 1571 :  32 - 0x20
      11'h624: dout <= 8'b00100000; // 1572 :  32 - 0x20
      11'h625: dout <= 8'b00100000; // 1573 :  32 - 0x20
      11'h626: dout <= 8'b00100000; // 1574 :  32 - 0x20
      11'h627: dout <= 8'b00100000; // 1575 :  32 - 0x20
      11'h628: dout <= 8'b00100000; // 1576 :  32 - 0x20
      11'h629: dout <= 8'b00100000; // 1577 :  32 - 0x20
      11'h62A: dout <= 8'b00100000; // 1578 :  32 - 0x20
      11'h62B: dout <= 8'b00100000; // 1579 :  32 - 0x20
      11'h62C: dout <= 8'b00100000; // 1580 :  32 - 0x20
      11'h62D: dout <= 8'b00100000; // 1581 :  32 - 0x20
      11'h62E: dout <= 8'b00100000; // 1582 :  32 - 0x20
      11'h62F: dout <= 8'b00100000; // 1583 :  32 - 0x20
      11'h630: dout <= 8'b00100000; // 1584 :  32 - 0x20
      11'h631: dout <= 8'b00100000; // 1585 :  32 - 0x20
      11'h632: dout <= 8'b00100000; // 1586 :  32 - 0x20
      11'h633: dout <= 8'b00100000; // 1587 :  32 - 0x20
      11'h634: dout <= 8'b00100000; // 1588 :  32 - 0x20
      11'h635: dout <= 8'b00100000; // 1589 :  32 - 0x20
      11'h636: dout <= 8'b00100000; // 1590 :  32 - 0x20
      11'h637: dout <= 8'b00100000; // 1591 :  32 - 0x20
      11'h638: dout <= 8'b00100000; // 1592 :  32 - 0x20
      11'h639: dout <= 8'b00100000; // 1593 :  32 - 0x20
      11'h63A: dout <= 8'b00100000; // 1594 :  32 - 0x20
      11'h63B: dout <= 8'b00100000; // 1595 :  32 - 0x20
      11'h63C: dout <= 8'b00100000; // 1596 :  32 - 0x20
      11'h63D: dout <= 8'b00100000; // 1597 :  32 - 0x20
      11'h63E: dout <= 8'b00100000; // 1598 :  32 - 0x20
      11'h63F: dout <= 8'b00100000; // 1599 :  32 - 0x20
      11'h640: dout <= 8'b00100000; // 1600 :  32 - 0x20 -- line 0x12
      11'h641: dout <= 8'b00100000; // 1601 :  32 - 0x20
      11'h642: dout <= 8'b00100000; // 1602 :  32 - 0x20
      11'h643: dout <= 8'b00100000; // 1603 :  32 - 0x20
      11'h644: dout <= 8'b00100000; // 1604 :  32 - 0x20
      11'h645: dout <= 8'b00100000; // 1605 :  32 - 0x20
      11'h646: dout <= 8'b00100000; // 1606 :  32 - 0x20
      11'h647: dout <= 8'b00100000; // 1607 :  32 - 0x20
      11'h648: dout <= 8'b00100000; // 1608 :  32 - 0x20
      11'h649: dout <= 8'b00100000; // 1609 :  32 - 0x20
      11'h64A: dout <= 8'b00100000; // 1610 :  32 - 0x20
      11'h64B: dout <= 8'b00100000; // 1611 :  32 - 0x20
      11'h64C: dout <= 8'b00100000; // 1612 :  32 - 0x20
      11'h64D: dout <= 8'b00100000; // 1613 :  32 - 0x20
      11'h64E: dout <= 8'b00100000; // 1614 :  32 - 0x20
      11'h64F: dout <= 8'b00100000; // 1615 :  32 - 0x20
      11'h650: dout <= 8'b00100000; // 1616 :  32 - 0x20
      11'h651: dout <= 8'b00100000; // 1617 :  32 - 0x20
      11'h652: dout <= 8'b00100000; // 1618 :  32 - 0x20
      11'h653: dout <= 8'b00100000; // 1619 :  32 - 0x20
      11'h654: dout <= 8'b00100000; // 1620 :  32 - 0x20
      11'h655: dout <= 8'b00100000; // 1621 :  32 - 0x20
      11'h656: dout <= 8'b00100000; // 1622 :  32 - 0x20
      11'h657: dout <= 8'b00100000; // 1623 :  32 - 0x20
      11'h658: dout <= 8'b00100000; // 1624 :  32 - 0x20
      11'h659: dout <= 8'b00100000; // 1625 :  32 - 0x20
      11'h65A: dout <= 8'b00100000; // 1626 :  32 - 0x20
      11'h65B: dout <= 8'b00100000; // 1627 :  32 - 0x20
      11'h65C: dout <= 8'b00100000; // 1628 :  32 - 0x20
      11'h65D: dout <= 8'b00100000; // 1629 :  32 - 0x20
      11'h65E: dout <= 8'b00100000; // 1630 :  32 - 0x20
      11'h65F: dout <= 8'b00100000; // 1631 :  32 - 0x20
      11'h660: dout <= 8'b00100000; // 1632 :  32 - 0x20 -- line 0x13
      11'h661: dout <= 8'b00100000; // 1633 :  32 - 0x20
      11'h662: dout <= 8'b00100000; // 1634 :  32 - 0x20
      11'h663: dout <= 8'b00100000; // 1635 :  32 - 0x20
      11'h664: dout <= 8'b00100000; // 1636 :  32 - 0x20
      11'h665: dout <= 8'b00100000; // 1637 :  32 - 0x20
      11'h666: dout <= 8'b00100000; // 1638 :  32 - 0x20
      11'h667: dout <= 8'b00100000; // 1639 :  32 - 0x20
      11'h668: dout <= 8'b00100000; // 1640 :  32 - 0x20
      11'h669: dout <= 8'b00100000; // 1641 :  32 - 0x20
      11'h66A: dout <= 8'b00100000; // 1642 :  32 - 0x20
      11'h66B: dout <= 8'b00100000; // 1643 :  32 - 0x20
      11'h66C: dout <= 8'b00100000; // 1644 :  32 - 0x20
      11'h66D: dout <= 8'b00100000; // 1645 :  32 - 0x20
      11'h66E: dout <= 8'b00100000; // 1646 :  32 - 0x20
      11'h66F: dout <= 8'b00100000; // 1647 :  32 - 0x20
      11'h670: dout <= 8'b00100000; // 1648 :  32 - 0x20
      11'h671: dout <= 8'b00100000; // 1649 :  32 - 0x20
      11'h672: dout <= 8'b00100000; // 1650 :  32 - 0x20
      11'h673: dout <= 8'b00100000; // 1651 :  32 - 0x20
      11'h674: dout <= 8'b00100000; // 1652 :  32 - 0x20
      11'h675: dout <= 8'b00100000; // 1653 :  32 - 0x20
      11'h676: dout <= 8'b00100000; // 1654 :  32 - 0x20
      11'h677: dout <= 8'b00100000; // 1655 :  32 - 0x20
      11'h678: dout <= 8'b00100000; // 1656 :  32 - 0x20
      11'h679: dout <= 8'b00100000; // 1657 :  32 - 0x20
      11'h67A: dout <= 8'b00100000; // 1658 :  32 - 0x20
      11'h67B: dout <= 8'b00100000; // 1659 :  32 - 0x20
      11'h67C: dout <= 8'b00100000; // 1660 :  32 - 0x20
      11'h67D: dout <= 8'b00100000; // 1661 :  32 - 0x20
      11'h67E: dout <= 8'b00100000; // 1662 :  32 - 0x20
      11'h67F: dout <= 8'b00100000; // 1663 :  32 - 0x20
      11'h680: dout <= 8'b00100000; // 1664 :  32 - 0x20 -- line 0x14
      11'h681: dout <= 8'b00100000; // 1665 :  32 - 0x20
      11'h682: dout <= 8'b00100000; // 1666 :  32 - 0x20
      11'h683: dout <= 8'b00100000; // 1667 :  32 - 0x20
      11'h684: dout <= 8'b00100000; // 1668 :  32 - 0x20
      11'h685: dout <= 8'b00100000; // 1669 :  32 - 0x20
      11'h686: dout <= 8'b00100000; // 1670 :  32 - 0x20
      11'h687: dout <= 8'b00100000; // 1671 :  32 - 0x20
      11'h688: dout <= 8'b00100000; // 1672 :  32 - 0x20
      11'h689: dout <= 8'b00100000; // 1673 :  32 - 0x20
      11'h68A: dout <= 8'b00100000; // 1674 :  32 - 0x20
      11'h68B: dout <= 8'b00100000; // 1675 :  32 - 0x20
      11'h68C: dout <= 8'b00100000; // 1676 :  32 - 0x20
      11'h68D: dout <= 8'b00100000; // 1677 :  32 - 0x20
      11'h68E: dout <= 8'b00100000; // 1678 :  32 - 0x20
      11'h68F: dout <= 8'b00100000; // 1679 :  32 - 0x20
      11'h690: dout <= 8'b00100000; // 1680 :  32 - 0x20
      11'h691: dout <= 8'b00100000; // 1681 :  32 - 0x20
      11'h692: dout <= 8'b00100000; // 1682 :  32 - 0x20
      11'h693: dout <= 8'b00100000; // 1683 :  32 - 0x20
      11'h694: dout <= 8'b00100000; // 1684 :  32 - 0x20
      11'h695: dout <= 8'b00100000; // 1685 :  32 - 0x20
      11'h696: dout <= 8'b00100000; // 1686 :  32 - 0x20
      11'h697: dout <= 8'b00100000; // 1687 :  32 - 0x20
      11'h698: dout <= 8'b00100000; // 1688 :  32 - 0x20
      11'h699: dout <= 8'b00100000; // 1689 :  32 - 0x20
      11'h69A: dout <= 8'b00100000; // 1690 :  32 - 0x20
      11'h69B: dout <= 8'b00100000; // 1691 :  32 - 0x20
      11'h69C: dout <= 8'b00100000; // 1692 :  32 - 0x20
      11'h69D: dout <= 8'b00100000; // 1693 :  32 - 0x20
      11'h69E: dout <= 8'b00100000; // 1694 :  32 - 0x20
      11'h69F: dout <= 8'b00100000; // 1695 :  32 - 0x20
      11'h6A0: dout <= 8'b00100000; // 1696 :  32 - 0x20 -- line 0x15
      11'h6A1: dout <= 8'b00100000; // 1697 :  32 - 0x20
      11'h6A2: dout <= 8'b00100000; // 1698 :  32 - 0x20
      11'h6A3: dout <= 8'b00100000; // 1699 :  32 - 0x20
      11'h6A4: dout <= 8'b00100000; // 1700 :  32 - 0x20
      11'h6A5: dout <= 8'b00100000; // 1701 :  32 - 0x20
      11'h6A6: dout <= 8'b00100000; // 1702 :  32 - 0x20
      11'h6A7: dout <= 8'b00100000; // 1703 :  32 - 0x20
      11'h6A8: dout <= 8'b00100000; // 1704 :  32 - 0x20
      11'h6A9: dout <= 8'b00100000; // 1705 :  32 - 0x20
      11'h6AA: dout <= 8'b00100000; // 1706 :  32 - 0x20
      11'h6AB: dout <= 8'b00100000; // 1707 :  32 - 0x20
      11'h6AC: dout <= 8'b00100000; // 1708 :  32 - 0x20
      11'h6AD: dout <= 8'b00100000; // 1709 :  32 - 0x20
      11'h6AE: dout <= 8'b00100000; // 1710 :  32 - 0x20
      11'h6AF: dout <= 8'b00100000; // 1711 :  32 - 0x20
      11'h6B0: dout <= 8'b00100000; // 1712 :  32 - 0x20
      11'h6B1: dout <= 8'b00100000; // 1713 :  32 - 0x20
      11'h6B2: dout <= 8'b00100000; // 1714 :  32 - 0x20
      11'h6B3: dout <= 8'b00100000; // 1715 :  32 - 0x20
      11'h6B4: dout <= 8'b00100000; // 1716 :  32 - 0x20
      11'h6B5: dout <= 8'b00100000; // 1717 :  32 - 0x20
      11'h6B6: dout <= 8'b00100000; // 1718 :  32 - 0x20
      11'h6B7: dout <= 8'b00100000; // 1719 :  32 - 0x20
      11'h6B8: dout <= 8'b00100000; // 1720 :  32 - 0x20
      11'h6B9: dout <= 8'b00100000; // 1721 :  32 - 0x20
      11'h6BA: dout <= 8'b00100000; // 1722 :  32 - 0x20
      11'h6BB: dout <= 8'b00100000; // 1723 :  32 - 0x20
      11'h6BC: dout <= 8'b00100000; // 1724 :  32 - 0x20
      11'h6BD: dout <= 8'b00100000; // 1725 :  32 - 0x20
      11'h6BE: dout <= 8'b00100000; // 1726 :  32 - 0x20
      11'h6BF: dout <= 8'b00100000; // 1727 :  32 - 0x20
      11'h6C0: dout <= 8'b00100000; // 1728 :  32 - 0x20 -- line 0x16
      11'h6C1: dout <= 8'b00100000; // 1729 :  32 - 0x20
      11'h6C2: dout <= 8'b00100000; // 1730 :  32 - 0x20
      11'h6C3: dout <= 8'b00100000; // 1731 :  32 - 0x20
      11'h6C4: dout <= 8'b00100000; // 1732 :  32 - 0x20
      11'h6C5: dout <= 8'b00100000; // 1733 :  32 - 0x20
      11'h6C6: dout <= 8'b00100000; // 1734 :  32 - 0x20
      11'h6C7: dout <= 8'b00100000; // 1735 :  32 - 0x20
      11'h6C8: dout <= 8'b00100000; // 1736 :  32 - 0x20
      11'h6C9: dout <= 8'b00100000; // 1737 :  32 - 0x20
      11'h6CA: dout <= 8'b00100000; // 1738 :  32 - 0x20
      11'h6CB: dout <= 8'b00100000; // 1739 :  32 - 0x20
      11'h6CC: dout <= 8'b00100000; // 1740 :  32 - 0x20
      11'h6CD: dout <= 8'b00100000; // 1741 :  32 - 0x20
      11'h6CE: dout <= 8'b00100000; // 1742 :  32 - 0x20
      11'h6CF: dout <= 8'b00100000; // 1743 :  32 - 0x20
      11'h6D0: dout <= 8'b00100000; // 1744 :  32 - 0x20
      11'h6D1: dout <= 8'b00100000; // 1745 :  32 - 0x20
      11'h6D2: dout <= 8'b00100000; // 1746 :  32 - 0x20
      11'h6D3: dout <= 8'b00100000; // 1747 :  32 - 0x20
      11'h6D4: dout <= 8'b00100000; // 1748 :  32 - 0x20
      11'h6D5: dout <= 8'b00100000; // 1749 :  32 - 0x20
      11'h6D6: dout <= 8'b00100000; // 1750 :  32 - 0x20
      11'h6D7: dout <= 8'b00100000; // 1751 :  32 - 0x20
      11'h6D8: dout <= 8'b00100000; // 1752 :  32 - 0x20
      11'h6D9: dout <= 8'b00100000; // 1753 :  32 - 0x20
      11'h6DA: dout <= 8'b00100000; // 1754 :  32 - 0x20
      11'h6DB: dout <= 8'b00100000; // 1755 :  32 - 0x20
      11'h6DC: dout <= 8'b00100000; // 1756 :  32 - 0x20
      11'h6DD: dout <= 8'b00100000; // 1757 :  32 - 0x20
      11'h6DE: dout <= 8'b00100000; // 1758 :  32 - 0x20
      11'h6DF: dout <= 8'b00100000; // 1759 :  32 - 0x20
      11'h6E0: dout <= 8'b00100000; // 1760 :  32 - 0x20 -- line 0x17
      11'h6E1: dout <= 8'b00100000; // 1761 :  32 - 0x20
      11'h6E2: dout <= 8'b00100000; // 1762 :  32 - 0x20
      11'h6E3: dout <= 8'b00100000; // 1763 :  32 - 0x20
      11'h6E4: dout <= 8'b00100000; // 1764 :  32 - 0x20
      11'h6E5: dout <= 8'b00100000; // 1765 :  32 - 0x20
      11'h6E6: dout <= 8'b00100000; // 1766 :  32 - 0x20
      11'h6E7: dout <= 8'b00100000; // 1767 :  32 - 0x20
      11'h6E8: dout <= 8'b00100000; // 1768 :  32 - 0x20
      11'h6E9: dout <= 8'b00100000; // 1769 :  32 - 0x20
      11'h6EA: dout <= 8'b00100000; // 1770 :  32 - 0x20
      11'h6EB: dout <= 8'b00100000; // 1771 :  32 - 0x20
      11'h6EC: dout <= 8'b00100000; // 1772 :  32 - 0x20
      11'h6ED: dout <= 8'b00100000; // 1773 :  32 - 0x20
      11'h6EE: dout <= 8'b00100000; // 1774 :  32 - 0x20
      11'h6EF: dout <= 8'b00100000; // 1775 :  32 - 0x20
      11'h6F0: dout <= 8'b00100000; // 1776 :  32 - 0x20
      11'h6F1: dout <= 8'b00100000; // 1777 :  32 - 0x20
      11'h6F2: dout <= 8'b00100000; // 1778 :  32 - 0x20
      11'h6F3: dout <= 8'b00100000; // 1779 :  32 - 0x20
      11'h6F4: dout <= 8'b00100000; // 1780 :  32 - 0x20
      11'h6F5: dout <= 8'b00100000; // 1781 :  32 - 0x20
      11'h6F6: dout <= 8'b00100000; // 1782 :  32 - 0x20
      11'h6F7: dout <= 8'b00100000; // 1783 :  32 - 0x20
      11'h6F8: dout <= 8'b00100000; // 1784 :  32 - 0x20
      11'h6F9: dout <= 8'b00100000; // 1785 :  32 - 0x20
      11'h6FA: dout <= 8'b00100000; // 1786 :  32 - 0x20
      11'h6FB: dout <= 8'b00100000; // 1787 :  32 - 0x20
      11'h6FC: dout <= 8'b00100000; // 1788 :  32 - 0x20
      11'h6FD: dout <= 8'b00100000; // 1789 :  32 - 0x20
      11'h6FE: dout <= 8'b00100000; // 1790 :  32 - 0x20
      11'h6FF: dout <= 8'b00100000; // 1791 :  32 - 0x20
      11'h700: dout <= 8'b00100000; // 1792 :  32 - 0x20 -- line 0x18
      11'h701: dout <= 8'b00100000; // 1793 :  32 - 0x20
      11'h702: dout <= 8'b00100000; // 1794 :  32 - 0x20
      11'h703: dout <= 8'b00100000; // 1795 :  32 - 0x20
      11'h704: dout <= 8'b00100000; // 1796 :  32 - 0x20
      11'h705: dout <= 8'b00100000; // 1797 :  32 - 0x20
      11'h706: dout <= 8'b00100000; // 1798 :  32 - 0x20
      11'h707: dout <= 8'b00100000; // 1799 :  32 - 0x20
      11'h708: dout <= 8'b00100000; // 1800 :  32 - 0x20
      11'h709: dout <= 8'b00100000; // 1801 :  32 - 0x20
      11'h70A: dout <= 8'b00100000; // 1802 :  32 - 0x20
      11'h70B: dout <= 8'b00100000; // 1803 :  32 - 0x20
      11'h70C: dout <= 8'b00100000; // 1804 :  32 - 0x20
      11'h70D: dout <= 8'b00100000; // 1805 :  32 - 0x20
      11'h70E: dout <= 8'b00100000; // 1806 :  32 - 0x20
      11'h70F: dout <= 8'b00100000; // 1807 :  32 - 0x20
      11'h710: dout <= 8'b00100000; // 1808 :  32 - 0x20
      11'h711: dout <= 8'b00100000; // 1809 :  32 - 0x20
      11'h712: dout <= 8'b00100000; // 1810 :  32 - 0x20
      11'h713: dout <= 8'b00100000; // 1811 :  32 - 0x20
      11'h714: dout <= 8'b00100000; // 1812 :  32 - 0x20
      11'h715: dout <= 8'b00100000; // 1813 :  32 - 0x20
      11'h716: dout <= 8'b00100000; // 1814 :  32 - 0x20
      11'h717: dout <= 8'b00100000; // 1815 :  32 - 0x20
      11'h718: dout <= 8'b00100000; // 1816 :  32 - 0x20
      11'h719: dout <= 8'b00100000; // 1817 :  32 - 0x20
      11'h71A: dout <= 8'b00100000; // 1818 :  32 - 0x20
      11'h71B: dout <= 8'b00100000; // 1819 :  32 - 0x20
      11'h71C: dout <= 8'b00100000; // 1820 :  32 - 0x20
      11'h71D: dout <= 8'b00100000; // 1821 :  32 - 0x20
      11'h71E: dout <= 8'b00100000; // 1822 :  32 - 0x20
      11'h71F: dout <= 8'b00100000; // 1823 :  32 - 0x20
      11'h720: dout <= 8'b00100000; // 1824 :  32 - 0x20 -- line 0x19
      11'h721: dout <= 8'b00100000; // 1825 :  32 - 0x20
      11'h722: dout <= 8'b00100000; // 1826 :  32 - 0x20
      11'h723: dout <= 8'b00100000; // 1827 :  32 - 0x20
      11'h724: dout <= 8'b00100000; // 1828 :  32 - 0x20
      11'h725: dout <= 8'b00100000; // 1829 :  32 - 0x20
      11'h726: dout <= 8'b00100000; // 1830 :  32 - 0x20
      11'h727: dout <= 8'b00100000; // 1831 :  32 - 0x20
      11'h728: dout <= 8'b00100000; // 1832 :  32 - 0x20
      11'h729: dout <= 8'b00100000; // 1833 :  32 - 0x20
      11'h72A: dout <= 8'b00100000; // 1834 :  32 - 0x20
      11'h72B: dout <= 8'b00100000; // 1835 :  32 - 0x20
      11'h72C: dout <= 8'b00100000; // 1836 :  32 - 0x20
      11'h72D: dout <= 8'b00100000; // 1837 :  32 - 0x20
      11'h72E: dout <= 8'b00100000; // 1838 :  32 - 0x20
      11'h72F: dout <= 8'b00100000; // 1839 :  32 - 0x20
      11'h730: dout <= 8'b00100000; // 1840 :  32 - 0x20
      11'h731: dout <= 8'b00100000; // 1841 :  32 - 0x20
      11'h732: dout <= 8'b00100000; // 1842 :  32 - 0x20
      11'h733: dout <= 8'b00100000; // 1843 :  32 - 0x20
      11'h734: dout <= 8'b00100000; // 1844 :  32 - 0x20
      11'h735: dout <= 8'b00100000; // 1845 :  32 - 0x20
      11'h736: dout <= 8'b00100000; // 1846 :  32 - 0x20
      11'h737: dout <= 8'b00100000; // 1847 :  32 - 0x20
      11'h738: dout <= 8'b00100000; // 1848 :  32 - 0x20
      11'h739: dout <= 8'b00100000; // 1849 :  32 - 0x20
      11'h73A: dout <= 8'b00100000; // 1850 :  32 - 0x20
      11'h73B: dout <= 8'b00100000; // 1851 :  32 - 0x20
      11'h73C: dout <= 8'b00100000; // 1852 :  32 - 0x20
      11'h73D: dout <= 8'b00100000; // 1853 :  32 - 0x20
      11'h73E: dout <= 8'b00100000; // 1854 :  32 - 0x20
      11'h73F: dout <= 8'b00100000; // 1855 :  32 - 0x20
      11'h740: dout <= 8'b00100000; // 1856 :  32 - 0x20 -- line 0x1a
      11'h741: dout <= 8'b00100000; // 1857 :  32 - 0x20
      11'h742: dout <= 8'b00100000; // 1858 :  32 - 0x20
      11'h743: dout <= 8'b00100000; // 1859 :  32 - 0x20
      11'h744: dout <= 8'b00100000; // 1860 :  32 - 0x20
      11'h745: dout <= 8'b00100000; // 1861 :  32 - 0x20
      11'h746: dout <= 8'b00100000; // 1862 :  32 - 0x20
      11'h747: dout <= 8'b00100000; // 1863 :  32 - 0x20
      11'h748: dout <= 8'b00100000; // 1864 :  32 - 0x20
      11'h749: dout <= 8'b00100000; // 1865 :  32 - 0x20
      11'h74A: dout <= 8'b00100000; // 1866 :  32 - 0x20
      11'h74B: dout <= 8'b00100000; // 1867 :  32 - 0x20
      11'h74C: dout <= 8'b00100000; // 1868 :  32 - 0x20
      11'h74D: dout <= 8'b00100000; // 1869 :  32 - 0x20
      11'h74E: dout <= 8'b00100000; // 1870 :  32 - 0x20
      11'h74F: dout <= 8'b00100000; // 1871 :  32 - 0x20
      11'h750: dout <= 8'b00100000; // 1872 :  32 - 0x20
      11'h751: dout <= 8'b00100000; // 1873 :  32 - 0x20
      11'h752: dout <= 8'b00100000; // 1874 :  32 - 0x20
      11'h753: dout <= 8'b00100000; // 1875 :  32 - 0x20
      11'h754: dout <= 8'b00100000; // 1876 :  32 - 0x20
      11'h755: dout <= 8'b00100000; // 1877 :  32 - 0x20
      11'h756: dout <= 8'b00100000; // 1878 :  32 - 0x20
      11'h757: dout <= 8'b00100000; // 1879 :  32 - 0x20
      11'h758: dout <= 8'b00100000; // 1880 :  32 - 0x20
      11'h759: dout <= 8'b00100000; // 1881 :  32 - 0x20
      11'h75A: dout <= 8'b00100000; // 1882 :  32 - 0x20
      11'h75B: dout <= 8'b00100000; // 1883 :  32 - 0x20
      11'h75C: dout <= 8'b00100000; // 1884 :  32 - 0x20
      11'h75D: dout <= 8'b00100000; // 1885 :  32 - 0x20
      11'h75E: dout <= 8'b00100000; // 1886 :  32 - 0x20
      11'h75F: dout <= 8'b00100000; // 1887 :  32 - 0x20
      11'h760: dout <= 8'b00100000; // 1888 :  32 - 0x20 -- line 0x1b
      11'h761: dout <= 8'b00100000; // 1889 :  32 - 0x20
      11'h762: dout <= 8'b00100000; // 1890 :  32 - 0x20
      11'h763: dout <= 8'b00100000; // 1891 :  32 - 0x20
      11'h764: dout <= 8'b00100000; // 1892 :  32 - 0x20
      11'h765: dout <= 8'b00100000; // 1893 :  32 - 0x20
      11'h766: dout <= 8'b00100000; // 1894 :  32 - 0x20
      11'h767: dout <= 8'b00100000; // 1895 :  32 - 0x20
      11'h768: dout <= 8'b00100000; // 1896 :  32 - 0x20
      11'h769: dout <= 8'b00100000; // 1897 :  32 - 0x20
      11'h76A: dout <= 8'b00100000; // 1898 :  32 - 0x20
      11'h76B: dout <= 8'b00100000; // 1899 :  32 - 0x20
      11'h76C: dout <= 8'b00100000; // 1900 :  32 - 0x20
      11'h76D: dout <= 8'b00100000; // 1901 :  32 - 0x20
      11'h76E: dout <= 8'b00100000; // 1902 :  32 - 0x20
      11'h76F: dout <= 8'b00100000; // 1903 :  32 - 0x20
      11'h770: dout <= 8'b00100000; // 1904 :  32 - 0x20
      11'h771: dout <= 8'b00100000; // 1905 :  32 - 0x20
      11'h772: dout <= 8'b00100000; // 1906 :  32 - 0x20
      11'h773: dout <= 8'b00100000; // 1907 :  32 - 0x20
      11'h774: dout <= 8'b00100000; // 1908 :  32 - 0x20
      11'h775: dout <= 8'b00100000; // 1909 :  32 - 0x20
      11'h776: dout <= 8'b00100000; // 1910 :  32 - 0x20
      11'h777: dout <= 8'b00100000; // 1911 :  32 - 0x20
      11'h778: dout <= 8'b00100000; // 1912 :  32 - 0x20
      11'h779: dout <= 8'b00100000; // 1913 :  32 - 0x20
      11'h77A: dout <= 8'b00100000; // 1914 :  32 - 0x20
      11'h77B: dout <= 8'b00100000; // 1915 :  32 - 0x20
      11'h77C: dout <= 8'b00100000; // 1916 :  32 - 0x20
      11'h77D: dout <= 8'b00100000; // 1917 :  32 - 0x20
      11'h77E: dout <= 8'b00100000; // 1918 :  32 - 0x20
      11'h77F: dout <= 8'b00100000; // 1919 :  32 - 0x20
      11'h780: dout <= 8'b00100000; // 1920 :  32 - 0x20 -- line 0x1c
      11'h781: dout <= 8'b00100000; // 1921 :  32 - 0x20
      11'h782: dout <= 8'b00100000; // 1922 :  32 - 0x20
      11'h783: dout <= 8'b00100000; // 1923 :  32 - 0x20
      11'h784: dout <= 8'b00100000; // 1924 :  32 - 0x20
      11'h785: dout <= 8'b00100000; // 1925 :  32 - 0x20
      11'h786: dout <= 8'b00100000; // 1926 :  32 - 0x20
      11'h787: dout <= 8'b00100000; // 1927 :  32 - 0x20
      11'h788: dout <= 8'b00100000; // 1928 :  32 - 0x20
      11'h789: dout <= 8'b00100000; // 1929 :  32 - 0x20
      11'h78A: dout <= 8'b00100000; // 1930 :  32 - 0x20
      11'h78B: dout <= 8'b00100000; // 1931 :  32 - 0x20
      11'h78C: dout <= 8'b00100000; // 1932 :  32 - 0x20
      11'h78D: dout <= 8'b00100000; // 1933 :  32 - 0x20
      11'h78E: dout <= 8'b00100000; // 1934 :  32 - 0x20
      11'h78F: dout <= 8'b00100000; // 1935 :  32 - 0x20
      11'h790: dout <= 8'b00100000; // 1936 :  32 - 0x20
      11'h791: dout <= 8'b00100000; // 1937 :  32 - 0x20
      11'h792: dout <= 8'b00100000; // 1938 :  32 - 0x20
      11'h793: dout <= 8'b00100000; // 1939 :  32 - 0x20
      11'h794: dout <= 8'b00100000; // 1940 :  32 - 0x20
      11'h795: dout <= 8'b00100000; // 1941 :  32 - 0x20
      11'h796: dout <= 8'b00100000; // 1942 :  32 - 0x20
      11'h797: dout <= 8'b00100000; // 1943 :  32 - 0x20
      11'h798: dout <= 8'b00100000; // 1944 :  32 - 0x20
      11'h799: dout <= 8'b00100000; // 1945 :  32 - 0x20
      11'h79A: dout <= 8'b00100000; // 1946 :  32 - 0x20
      11'h79B: dout <= 8'b00100000; // 1947 :  32 - 0x20
      11'h79C: dout <= 8'b00100000; // 1948 :  32 - 0x20
      11'h79D: dout <= 8'b00100000; // 1949 :  32 - 0x20
      11'h79E: dout <= 8'b00100000; // 1950 :  32 - 0x20
      11'h79F: dout <= 8'b00100000; // 1951 :  32 - 0x20
      11'h7A0: dout <= 8'b00100000; // 1952 :  32 - 0x20 -- line 0x1d
      11'h7A1: dout <= 8'b00100000; // 1953 :  32 - 0x20
      11'h7A2: dout <= 8'b00100000; // 1954 :  32 - 0x20
      11'h7A3: dout <= 8'b00100000; // 1955 :  32 - 0x20
      11'h7A4: dout <= 8'b00100000; // 1956 :  32 - 0x20
      11'h7A5: dout <= 8'b00100000; // 1957 :  32 - 0x20
      11'h7A6: dout <= 8'b00100000; // 1958 :  32 - 0x20
      11'h7A7: dout <= 8'b00100000; // 1959 :  32 - 0x20
      11'h7A8: dout <= 8'b00100000; // 1960 :  32 - 0x20
      11'h7A9: dout <= 8'b00100000; // 1961 :  32 - 0x20
      11'h7AA: dout <= 8'b00100000; // 1962 :  32 - 0x20
      11'h7AB: dout <= 8'b00100000; // 1963 :  32 - 0x20
      11'h7AC: dout <= 8'b00100000; // 1964 :  32 - 0x20
      11'h7AD: dout <= 8'b00100000; // 1965 :  32 - 0x20
      11'h7AE: dout <= 8'b00100000; // 1966 :  32 - 0x20
      11'h7AF: dout <= 8'b00100000; // 1967 :  32 - 0x20
      11'h7B0: dout <= 8'b00100000; // 1968 :  32 - 0x20
      11'h7B1: dout <= 8'b00100000; // 1969 :  32 - 0x20
      11'h7B2: dout <= 8'b00100000; // 1970 :  32 - 0x20
      11'h7B3: dout <= 8'b00100000; // 1971 :  32 - 0x20
      11'h7B4: dout <= 8'b00100000; // 1972 :  32 - 0x20
      11'h7B5: dout <= 8'b00100000; // 1973 :  32 - 0x20
      11'h7B6: dout <= 8'b00100000; // 1974 :  32 - 0x20
      11'h7B7: dout <= 8'b00100000; // 1975 :  32 - 0x20
      11'h7B8: dout <= 8'b00100000; // 1976 :  32 - 0x20
      11'h7B9: dout <= 8'b00100000; // 1977 :  32 - 0x20
      11'h7BA: dout <= 8'b00100000; // 1978 :  32 - 0x20
      11'h7BB: dout <= 8'b00100000; // 1979 :  32 - 0x20
      11'h7BC: dout <= 8'b00100000; // 1980 :  32 - 0x20
      11'h7BD: dout <= 8'b00100000; // 1981 :  32 - 0x20
      11'h7BE: dout <= 8'b00100000; // 1982 :  32 - 0x20
      11'h7BF: dout <= 8'b00100000; // 1983 :  32 - 0x20
        //-- Attribute Table 1----
      11'h7C0: dout <= 8'b01010101; // 1984 :  85 - 0x55
      11'h7C1: dout <= 8'b01010101; // 1985 :  85 - 0x55
      11'h7C2: dout <= 8'b01010101; // 1986 :  85 - 0x55
      11'h7C3: dout <= 8'b01010101; // 1987 :  85 - 0x55
      11'h7C4: dout <= 8'b01010101; // 1988 :  85 - 0x55
      11'h7C5: dout <= 8'b00010001; // 1989 :  17 - 0x11
      11'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b01010101; // 1992 :  85 - 0x55
      11'h7C9: dout <= 8'b01010101; // 1993 :  85 - 0x55
      11'h7CA: dout <= 8'b01010101; // 1994 :  85 - 0x55
      11'h7CB: dout <= 8'b01010101; // 1995 :  85 - 0x55
      11'h7CC: dout <= 8'b01010101; // 1996 :  85 - 0x55
      11'h7CD: dout <= 8'b00010001; // 1997 :  17 - 0x11
      11'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout <= 8'b01010101; // 2000 :  85 - 0x55
      11'h7D1: dout <= 8'b01010101; // 2001 :  85 - 0x55
      11'h7D2: dout <= 8'b01010101; // 2002 :  85 - 0x55
      11'h7D3: dout <= 8'b01010101; // 2003 :  85 - 0x55
      11'h7D4: dout <= 8'b01010101; // 2004 :  85 - 0x55
      11'h7D5: dout <= 8'b00010001; // 2005 :  17 - 0x11
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b01010101; // 2008 :  85 - 0x55
      11'h7D9: dout <= 8'b01010101; // 2009 :  85 - 0x55
      11'h7DA: dout <= 8'b01010101; // 2010 :  85 - 0x55
      11'h7DB: dout <= 8'b01010101; // 2011 :  85 - 0x55
      11'h7DC: dout <= 8'b01010101; // 2012 :  85 - 0x55
      11'h7DD: dout <= 8'b01010001; // 2013 :  81 - 0x51
      11'h7DE: dout <= 8'b01010000; // 2014 :  80 - 0x50
      11'h7DF: dout <= 8'b01010000; // 2015 :  80 - 0x50
      11'h7E0: dout <= 8'b01010101; // 2016 :  85 - 0x55
      11'h7E1: dout <= 8'b01010101; // 2017 :  85 - 0x55
      11'h7E2: dout <= 8'b01010101; // 2018 :  85 - 0x55
      11'h7E3: dout <= 8'b01010101; // 2019 :  85 - 0x55
      11'h7E4: dout <= 8'b01010101; // 2020 :  85 - 0x55
      11'h7E5: dout <= 8'b00010001; // 2021 :  17 - 0x11
      11'h7E6: dout <= 8'b00000101; // 2022 :   5 - 0x5
      11'h7E7: dout <= 8'b00000101; // 2023 :   5 - 0x5
      11'h7E8: dout <= 8'b01010101; // 2024 :  85 - 0x55
      11'h7E9: dout <= 8'b01010101; // 2025 :  85 - 0x55
      11'h7EA: dout <= 8'b01010101; // 2026 :  85 - 0x55
      11'h7EB: dout <= 8'b01010101; // 2027 :  85 - 0x55
      11'h7EC: dout <= 8'b01010101; // 2028 :  85 - 0x55
      11'h7ED: dout <= 8'b00010001; // 2029 :  17 - 0x11
      11'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout <= 8'b01010101; // 2032 :  85 - 0x55
      11'h7F1: dout <= 8'b01010101; // 2033 :  85 - 0x55
      11'h7F2: dout <= 8'b01010101; // 2034 :  85 - 0x55
      11'h7F3: dout <= 8'b01010101; // 2035 :  85 - 0x55
      11'h7F4: dout <= 8'b01010101; // 2036 :  85 - 0x55
      11'h7F5: dout <= 8'b01010101; // 2037 :  85 - 0x55
      11'h7F6: dout <= 8'b01010101; // 2038 :  85 - 0x55
      11'h7F7: dout <= 8'b01010101; // 2039 :  85 - 0x55
      11'h7F8: dout <= 8'b01010101; // 2040 :  85 - 0x55
      11'h7F9: dout <= 8'b01010101; // 2041 :  85 - 0x55
      11'h7FA: dout <= 8'b01010101; // 2042 :  85 - 0x55
      11'h7FB: dout <= 8'b01010101; // 2043 :  85 - 0x55
      11'h7FC: dout <= 8'b01010101; // 2044 :  85 - 0x55
      11'h7FD: dout <= 8'b01010101; // 2045 :  85 - 0x55
      11'h7FE: dout <= 8'b01010101; // 2046 :  85 - 0x55
      11'h7FF: dout <= 8'b01010101; // 2047 :  85 - 0x55
    endcase
  end

endmodule
