//- Autcmatically generated verilog ROM from a NES memory file----
//-   SPRITEs MEMORY (OAM)
// https://wiki.nesdev.com/w/index.php/PPU_OAM


//-  Original memory dump file name: donkeykong_oam.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_OAM_DONKEYKONG
  (
     input     clk,   // clock
     input      [8-1:0] addr,  //256 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
      8'h0: dout <= 8'b01101011; //    0 : 107 - 0x6b -- Sprite 0x0
      8'h1: dout <= 8'b00000110; //    1 :   6 - 0x6
      8'h2: dout <= 8'b01000000; //    2 :  64 - 0x40
      8'h3: dout <= 8'b01110011; //    3 : 115 - 0x73
      8'h4: dout <= 8'b01110011; //    4 : 115 - 0x73 -- Sprite 0x1
      8'h5: dout <= 8'b00000111; //    5 :   7 - 0x7
      8'h6: dout <= 8'b01000000; //    6 :  64 - 0x40
      8'h7: dout <= 8'b01110011; //    7 : 115 - 0x73
      8'h8: dout <= 8'b01101011; //    8 : 107 - 0x6b -- Sprite 0x2
      8'h9: dout <= 8'b00000100; //    9 :   4 - 0x4
      8'hA: dout <= 8'b01000000; //   10 :  64 - 0x40
      8'hB: dout <= 8'b01111011; //   11 : 123 - 0x7b
      8'hC: dout <= 8'b01110011; //   12 : 115 - 0x73 -- Sprite 0x3
      8'hD: dout <= 8'b00000101; //   13 :   5 - 0x5
      8'hE: dout <= 8'b01000000; //   14 :  64 - 0x40
      8'hF: dout <= 8'b01111011; //   15 : 123 - 0x7b
      8'h10: dout <= 8'b10100101; //   16 : 165 - 0xa5 -- Sprite 0x4
      8'h11: dout <= 8'b10011010; //   17 : 154 - 0x9a
      8'h12: dout <= 8'b01000010; //   18 :  66 - 0x42
      8'h13: dout <= 8'b01001011; //   19 :  75 - 0x4b
      8'h14: dout <= 8'b10101101; //   20 : 173 - 0xad -- Sprite 0x5
      8'h15: dout <= 8'b10011011; //   21 : 155 - 0x9b
      8'h16: dout <= 8'b01000010; //   22 :  66 - 0x42
      8'h17: dout <= 8'b01001011; //   23 :  75 - 0x4b
      8'h18: dout <= 8'b10100101; //   24 : 165 - 0xa5 -- Sprite 0x6
      8'h19: dout <= 8'b10011000; //   25 : 152 - 0x98
      8'h1A: dout <= 8'b01000010; //   26 :  66 - 0x42
      8'h1B: dout <= 8'b01010011; //   27 :  83 - 0x53
      8'h1C: dout <= 8'b10101101; //   28 : 173 - 0xad -- Sprite 0x7
      8'h1D: dout <= 8'b10011001; //   29 : 153 - 0x99
      8'h1E: dout <= 8'b01000010; //   30 :  66 - 0x42
      8'h1F: dout <= 8'b01010011; //   31 :  83 - 0x53
      8'h20: dout <= 8'b11000111; //   32 : 199 - 0xc7 -- Sprite 0x8
      8'h21: dout <= 8'b10011110; //   33 : 158 - 0x9e
      8'h22: dout <= 8'b01000010; //   34 :  66 - 0x42
      8'h23: dout <= 8'b01001100; //   35 :  76 - 0x4c
      8'h24: dout <= 8'b11001111; //   36 : 207 - 0xcf -- Sprite 0x9
      8'h25: dout <= 8'b10011111; //   37 : 159 - 0x9f
      8'h26: dout <= 8'b01000010; //   38 :  66 - 0x42
      8'h27: dout <= 8'b01001100; //   39 :  76 - 0x4c
      8'h28: dout <= 8'b11000111; //   40 : 199 - 0xc7 -- Sprite 0xa
      8'h29: dout <= 8'b10011100; //   41 : 156 - 0x9c
      8'h2A: dout <= 8'b01000010; //   42 :  66 - 0x42
      8'h2B: dout <= 8'b01010100; //   43 :  84 - 0x54
      8'h2C: dout <= 8'b11001111; //   44 : 207 - 0xcf -- Sprite 0xb
      8'h2D: dout <= 8'b10011101; //   45 : 157 - 0x9d
      8'h2E: dout <= 8'b01000010; //   46 :  66 - 0x42
      8'h2F: dout <= 8'b01010100; //   47 :  84 - 0x54
      8'h30: dout <= 8'b10001010; //   48 : 138 - 0x8a -- Sprite 0xc
      8'h31: dout <= 8'b10001000; //   49 : 136 - 0x88
      8'h32: dout <= 8'b00000011; //   50 :   3 - 0x3
      8'h33: dout <= 8'b10111010; //   51 : 186 - 0xba
      8'h34: dout <= 8'b10010010; //   52 : 146 - 0x92 -- Sprite 0xd
      8'h35: dout <= 8'b10001001; //   53 : 137 - 0x89
      8'h36: dout <= 8'b00000011; //   54 :   3 - 0x3
      8'h37: dout <= 8'b10111010; //   55 : 186 - 0xba
      8'h38: dout <= 8'b10001010; //   56 : 138 - 0x8a -- Sprite 0xe
      8'h39: dout <= 8'b10001010; //   57 : 138 - 0x8a
      8'h3A: dout <= 8'b00000011; //   58 :   3 - 0x3
      8'h3B: dout <= 8'b11000010; //   59 : 194 - 0xc2
      8'h3C: dout <= 8'b10010010; //   60 : 146 - 0x92 -- Sprite 0xf
      8'h3D: dout <= 8'b10001011; //   61 : 139 - 0x8b
      8'h3E: dout <= 8'b00000011; //   62 :   3 - 0x3
      8'h3F: dout <= 8'b11000010; //   63 : 194 - 0xc2
      8'h40: dout <= 8'b10000111; //   64 : 135 - 0x87 -- Sprite 0x10
      8'h41: dout <= 8'b10001000; //   65 : 136 - 0x88
      8'h42: dout <= 8'b00000011; //   66 :   3 - 0x3
      8'h43: dout <= 8'b11100110; //   67 : 230 - 0xe6
      8'h44: dout <= 8'b10001111; //   68 : 143 - 0x8f -- Sprite 0x11
      8'h45: dout <= 8'b10001001; //   69 : 137 - 0x89
      8'h46: dout <= 8'b00000011; //   70 :   3 - 0x3
      8'h47: dout <= 8'b11100110; //   71 : 230 - 0xe6
      8'h48: dout <= 8'b10000111; //   72 : 135 - 0x87 -- Sprite 0x12
      8'h49: dout <= 8'b10001010; //   73 : 138 - 0x8a
      8'h4A: dout <= 8'b00000011; //   74 :   3 - 0x3
      8'h4B: dout <= 8'b11101110; //   75 : 238 - 0xee
      8'h4C: dout <= 8'b10001111; //   76 : 143 - 0x8f -- Sprite 0x13
      8'h4D: dout <= 8'b10001011; //   77 : 139 - 0x8b
      8'h4E: dout <= 8'b00000011; //   78 :   3 - 0x3
      8'h4F: dout <= 8'b11101110; //   79 : 238 - 0xee
      8'h50: dout <= 8'b01010011; //   80 :  83 - 0x53 -- Sprite 0x14
      8'h51: dout <= 8'b10000000; //   81 : 128 - 0x80
      8'h52: dout <= 8'b00000011; //   82 :   3 - 0x3
      8'h53: dout <= 8'b00110010; //   83 :  50 - 0x32
      8'h54: dout <= 8'b01011011; //   84 :  91 - 0x5b -- Sprite 0x15
      8'h55: dout <= 8'b10000001; //   85 : 129 - 0x81
      8'h56: dout <= 8'b00000011; //   86 :   3 - 0x3
      8'h57: dout <= 8'b00110010; //   87 :  50 - 0x32
      8'h58: dout <= 8'b01010011; //   88 :  83 - 0x53 -- Sprite 0x16
      8'h59: dout <= 8'b10000010; //   89 : 130 - 0x82
      8'h5A: dout <= 8'b00000011; //   90 :   3 - 0x3
      8'h5B: dout <= 8'b00111010; //   91 :  58 - 0x3a
      8'h5C: dout <= 8'b01011011; //   92 :  91 - 0x5b -- Sprite 0x17
      8'h5D: dout <= 8'b10000011; //   93 : 131 - 0x83
      8'h5E: dout <= 8'b00000011; //   94 :   3 - 0x3
      8'h5F: dout <= 8'b00111010; //   95 :  58 - 0x3a
      8'h60: dout <= 8'b01001001; //   96 :  73 - 0x49 -- Sprite 0x18
      8'h61: dout <= 8'b10001000; //   97 : 136 - 0x88
      8'h62: dout <= 8'b00000011; //   98 :   3 - 0x3
      8'h63: dout <= 8'b11011101; //   99 : 221 - 0xdd
      8'h64: dout <= 8'b01010001; //  100 :  81 - 0x51 -- Sprite 0x19
      8'h65: dout <= 8'b10001001; //  101 : 137 - 0x89
      8'h66: dout <= 8'b00000011; //  102 :   3 - 0x3
      8'h67: dout <= 8'b11011101; //  103 : 221 - 0xdd
      8'h68: dout <= 8'b01001001; //  104 :  73 - 0x49 -- Sprite 0x1a
      8'h69: dout <= 8'b10001010; //  105 : 138 - 0x8a
      8'h6A: dout <= 8'b00000011; //  106 :   3 - 0x3
      8'h6B: dout <= 8'b11100101; //  107 : 229 - 0xe5
      8'h6C: dout <= 8'b01010001; //  108 :  81 - 0x51 -- Sprite 0x1b
      8'h6D: dout <= 8'b10001011; //  109 : 139 - 0x8b
      8'h6E: dout <= 8'b00000011; //  110 :   3 - 0x3
      8'h6F: dout <= 8'b11100101; //  111 : 229 - 0xe5
      8'h70: dout <= 8'b00110010; //  112 :  50 - 0x32 -- Sprite 0x1c
      8'h71: dout <= 8'b10000100; //  113 : 132 - 0x84
      8'h72: dout <= 8'b00000011; //  114 :   3 - 0x3
      8'h73: dout <= 8'b01001101; //  115 :  77 - 0x4d
      8'h74: dout <= 8'b00111010; //  116 :  58 - 0x3a -- Sprite 0x1d
      8'h75: dout <= 8'b10000101; //  117 : 133 - 0x85
      8'h76: dout <= 8'b00000011; //  118 :   3 - 0x3
      8'h77: dout <= 8'b01001101; //  119 :  77 - 0x4d
      8'h78: dout <= 8'b00110010; //  120 :  50 - 0x32 -- Sprite 0x1e
      8'h79: dout <= 8'b10000110; //  121 : 134 - 0x86
      8'h7A: dout <= 8'b00000011; //  122 :   3 - 0x3
      8'h7B: dout <= 8'b01010101; //  123 :  85 - 0x55
      8'h7C: dout <= 8'b00111010; //  124 :  58 - 0x3a -- Sprite 0x1f
      8'h7D: dout <= 8'b10000111; //  125 : 135 - 0x87
      8'h7E: dout <= 8'b00000011; //  126 :   3 - 0x3
      8'h7F: dout <= 8'b01010101; //  127 :  85 - 0x55
      8'h80: dout <= 8'b11111111; //  128 : 255 - 0xff -- Sprite 0x20
      8'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      8'h82: dout <= 8'b00000011; //  130 :   3 - 0x3
      8'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      8'h84: dout <= 8'b11111111; //  132 : 255 - 0xff -- Sprite 0x21
      8'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      8'h86: dout <= 8'b00000011; //  134 :   3 - 0x3
      8'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      8'h88: dout <= 8'b11111111; //  136 : 255 - 0xff -- Sprite 0x22
      8'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      8'h8A: dout <= 8'b00000011; //  138 :   3 - 0x3
      8'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      8'h8C: dout <= 8'b11111111; //  140 : 255 - 0xff -- Sprite 0x23
      8'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      8'h8E: dout <= 8'b00000011; //  142 :   3 - 0x3
      8'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      8'h90: dout <= 8'b11111111; //  144 : 255 - 0xff -- Sprite 0x24
      8'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      8'h92: dout <= 8'b00000011; //  146 :   3 - 0x3
      8'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      8'h94: dout <= 8'b11111111; //  148 : 255 - 0xff -- Sprite 0x25
      8'h95: dout <= 8'b00000000; //  149 :   0 - 0x0
      8'h96: dout <= 8'b00000011; //  150 :   3 - 0x3
      8'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      8'h98: dout <= 8'b11111111; //  152 : 255 - 0xff -- Sprite 0x26
      8'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      8'h9A: dout <= 8'b00000011; //  154 :   3 - 0x3
      8'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      8'h9C: dout <= 8'b11111111; //  156 : 255 - 0xff -- Sprite 0x27
      8'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      8'h9E: dout <= 8'b00000011; //  158 :   3 - 0x3
      8'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      8'hA0: dout <= 8'b11111111; //  160 : 255 - 0xff -- Sprite 0x28
      8'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      8'hA2: dout <= 8'b00000011; //  162 :   3 - 0x3
      8'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      8'hA4: dout <= 8'b11111111; //  164 : 255 - 0xff -- Sprite 0x29
      8'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      8'hA6: dout <= 8'b00000011; //  166 :   3 - 0x3
      8'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      8'hA8: dout <= 8'b11111111; //  168 : 255 - 0xff -- Sprite 0x2a
      8'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      8'hAA: dout <= 8'b00000011; //  170 :   3 - 0x3
      8'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      8'hAC: dout <= 8'b11111111; //  172 : 255 - 0xff -- Sprite 0x2b
      8'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      8'hAE: dout <= 8'b00000011; //  174 :   3 - 0x3
      8'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      8'hB0: dout <= 8'b11111111; //  176 : 255 - 0xff -- Sprite 0x2c
      8'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      8'hB2: dout <= 8'b00000011; //  178 :   3 - 0x3
      8'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      8'hB4: dout <= 8'b11111111; //  180 : 255 - 0xff -- Sprite 0x2d
      8'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      8'hB6: dout <= 8'b00000011; //  182 :   3 - 0x3
      8'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      8'hB8: dout <= 8'b11111111; //  184 : 255 - 0xff -- Sprite 0x2e
      8'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      8'hBA: dout <= 8'b00000011; //  186 :   3 - 0x3
      8'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      8'hBC: dout <= 8'b11111111; //  188 : 255 - 0xff -- Sprite 0x2f
      8'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      8'hBE: dout <= 8'b00000011; //  190 :   3 - 0x3
      8'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      8'hC0: dout <= 8'b11111111; //  192 : 255 - 0xff -- Sprite 0x30
      8'hC1: dout <= 8'b11010000; //  193 : 208 - 0xd0
      8'hC2: dout <= 8'b00000001; //  194 :   1 - 0x1
      8'hC3: dout <= 8'b01110100; //  195 : 116 - 0x74
      8'hC4: dout <= 8'b11111111; //  196 : 255 - 0xff -- Sprite 0x31
      8'hC5: dout <= 8'b11010100; //  197 : 212 - 0xd4
      8'hC6: dout <= 8'b00000001; //  198 :   1 - 0x1
      8'hC7: dout <= 8'b01111100; //  199 : 124 - 0x7c
      8'hC8: dout <= 8'b11111111; //  200 : 255 - 0xff -- Sprite 0x32
      8'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      8'hCA: dout <= 8'b00000001; //  202 :   1 - 0x1
      8'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      8'hCC: dout <= 8'b11111111; //  204 : 255 - 0xff -- Sprite 0x33
      8'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      8'hCE: dout <= 8'b00000001; //  206 :   1 - 0x1
      8'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      8'hD0: dout <= 8'b11111111; //  208 : 255 - 0xff -- Sprite 0x34
      8'hD1: dout <= 8'b11110110; //  209 : 246 - 0xf6
      8'hD2: dout <= 8'b00000011; //  210 :   3 - 0x3
      8'hD3: dout <= 8'b10100110; //  211 : 166 - 0xa6
      8'hD4: dout <= 8'b11111111; //  212 : 255 - 0xff -- Sprite 0x35
      8'hD5: dout <= 8'b11110111; //  213 : 247 - 0xf7
      8'hD6: dout <= 8'b00000011; //  214 :   3 - 0x3
      8'hD7: dout <= 8'b10100110; //  215 : 166 - 0xa6
      8'hD8: dout <= 8'b01000110; //  216 :  70 - 0x46 -- Sprite 0x36
      8'hD9: dout <= 8'b11110110; //  217 : 246 - 0xf6
      8'hDA: dout <= 8'b00000011; //  218 :   3 - 0x3
      8'hDB: dout <= 8'b00100000; //  219 :  32 - 0x20
      8'hDC: dout <= 8'b01001110; //  220 :  78 - 0x4e -- Sprite 0x37
      8'hDD: dout <= 8'b11110111; //  221 : 247 - 0xf7
      8'hDE: dout <= 8'b00000011; //  222 :   3 - 0x3
      8'hDF: dout <= 8'b00100000; //  223 :  32 - 0x20
      8'hE0: dout <= 8'b11000000; //  224 : 192 - 0xc0 -- Sprite 0x38
      8'hE1: dout <= 8'b11111110; //  225 : 254 - 0xfe
      8'hE2: dout <= 8'b00000010; //  226 :   2 - 0x2
      8'hE3: dout <= 8'b00100000; //  227 :  32 - 0x20
      8'hE4: dout <= 8'b11000000; //  228 : 192 - 0xc0 -- Sprite 0x39
      8'hE5: dout <= 8'b11111111; //  229 : 255 - 0xff
      8'hE6: dout <= 8'b00000010; //  230 :   2 - 0x2
      8'hE7: dout <= 8'b00101000; //  231 :  40 - 0x28
      8'hE8: dout <= 8'b00011000; //  232 :  24 - 0x18 -- Sprite 0x3a
      8'hE9: dout <= 8'b11010101; //  233 : 213 - 0xd5
      8'hEA: dout <= 8'b00000001; //  234 :   1 - 0x1
      8'hEB: dout <= 8'b01010000; //  235 :  80 - 0x50
      8'hEC: dout <= 8'b00011000; //  236 :  24 - 0x18 -- Sprite 0x3b
      8'hED: dout <= 8'b11010110; //  237 : 214 - 0xd6
      8'hEE: dout <= 8'b00000001; //  238 :   1 - 0x1
      8'hEF: dout <= 8'b01011000; //  239 :  88 - 0x58
      8'hF0: dout <= 8'b00100000; //  240 :  32 - 0x20 -- Sprite 0x3c
      8'hF1: dout <= 8'b11011011; //  241 : 219 - 0xdb
      8'hF2: dout <= 8'b00000001; //  242 :   1 - 0x1
      8'hF3: dout <= 8'b01010000; //  243 :  80 - 0x50
      8'hF4: dout <= 8'b00101000; //  244 :  40 - 0x28 -- Sprite 0x3d
      8'hF5: dout <= 8'b11011100; //  245 : 220 - 0xdc
      8'hF6: dout <= 8'b00000001; //  246 :   1 - 0x1
      8'hF7: dout <= 8'b01010000; //  247 :  80 - 0x50
      8'hF8: dout <= 8'b00100000; //  248 :  32 - 0x20 -- Sprite 0x3e
      8'hF9: dout <= 8'b11011101; //  249 : 221 - 0xdd
      8'hFA: dout <= 8'b00000001; //  250 :   1 - 0x1
      8'hFB: dout <= 8'b01011000; //  251 :  88 - 0x58
      8'hFC: dout <= 8'b00101000; //  252 :  40 - 0x28 -- Sprite 0x3f
      8'hFD: dout <= 8'b11011110; //  253 : 222 - 0xde
      8'hFE: dout <= 8'b00000001; //  254 :   1 - 0x1
      8'hFF: dout <= 8'b01011000; //  255 :  88 - 0x58
    endcase
  end

endmodule
