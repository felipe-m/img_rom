--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: lawnmower_ntable_start.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_LAWN_START is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_LAWN_START;

architecture BEHAVIORAL of ROM_NTABLE_LAWN_START is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "10000100", --    0 -  0x0  :  132 - 0x84 -- line 0x0
    "10000101", --    1 -  0x1  :  133 - 0x85
    "10000100", --    2 -  0x2  :  132 - 0x84
    "10000101", --    3 -  0x3  :  133 - 0x85
    "10000111", --    4 -  0x4  :  135 - 0x87
    "10000101", --    5 -  0x5  :  133 - 0x85
    "10000100", --    6 -  0x6  :  132 - 0x84
    "10000111", --    7 -  0x7  :  135 - 0x87
    "10000100", --    8 -  0x8  :  132 - 0x84
    "10000101", --    9 -  0x9  :  133 - 0x85
    "10000100", --   10 -  0xa  :  132 - 0x84
    "10000101", --   11 -  0xb  :  133 - 0x85
    "10000100", --   12 -  0xc  :  132 - 0x84
    "10000110", --   13 -  0xd  :  134 - 0x86
    "10000100", --   14 -  0xe  :  132 - 0x84
    "10010110", --   15 -  0xf  :  150 - 0x96
    "10000111", --   16 - 0x10  :  135 - 0x87
    "10000101", --   17 - 0x11  :  133 - 0x85
    "10000100", --   18 - 0x12  :  132 - 0x84
    "10010111", --   19 - 0x13  :  151 - 0x97
    "10000100", --   20 - 0x14  :  132 - 0x84
    "10000101", --   21 - 0x15  :  133 - 0x85
    "10000100", --   22 - 0x16  :  132 - 0x84
    "10000101", --   23 - 0x17  :  133 - 0x85
    "10000100", --   24 - 0x18  :  132 - 0x84
    "10000111", --   25 - 0x19  :  135 - 0x87
    "10000100", --   26 - 0x1a  :  132 - 0x84
    "10000101", --   27 - 0x1b  :  133 - 0x85
    "10000110", --   28 - 0x1c  :  134 - 0x86
    "10000101", --   29 - 0x1d  :  133 - 0x85
    "10000100", --   30 - 0x1e  :  132 - 0x84
    "10000101", --   31 - 0x1f  :  133 - 0x85
    "10010100", --   32 - 0x20  :  148 - 0x94 -- line 0x1
    "10000111", --   33 - 0x21  :  135 - 0x87
    "10010100", --   34 - 0x22  :  148 - 0x94
    "10000110", --   35 - 0x23  :  134 - 0x86
    "10010100", --   36 - 0x24  :  148 - 0x94
    "10010101", --   37 - 0x25  :  149 - 0x95
    "10010110", --   38 - 0x26  :  150 - 0x96
    "10010101", --   39 - 0x27  :  149 - 0x95
    "10010100", --   40 - 0x28  :  148 - 0x94
    "10010101", --   41 - 0x29  :  149 - 0x95
    "10010100", --   42 - 0x2a  :  148 - 0x94
    "10010111", --   43 - 0x2b  :  151 - 0x97
    "10010100", --   44 - 0x2c  :  148 - 0x94
    "10010101", --   45 - 0x2d  :  149 - 0x95
    "10010100", --   46 - 0x2e  :  148 - 0x94
    "10010101", --   47 - 0x2f  :  149 - 0x95
    "10010100", --   48 - 0x30  :  148 - 0x94
    "10000110", --   49 - 0x31  :  134 - 0x86
    "10010100", --   50 - 0x32  :  148 - 0x94
    "10010101", --   51 - 0x33  :  149 - 0x95
    "10010100", --   52 - 0x34  :  148 - 0x94
    "10010101", --   53 - 0x35  :  149 - 0x95
    "10010110", --   54 - 0x36  :  150 - 0x96
    "10010101", --   55 - 0x37  :  149 - 0x95
    "10000110", --   56 - 0x38  :  134 - 0x86
    "10010101", --   57 - 0x39  :  149 - 0x95
    "10010100", --   58 - 0x3a  :  148 - 0x94
    "10010111", --   59 - 0x3b  :  151 - 0x97
    "10010100", --   60 - 0x3c  :  148 - 0x94
    "10000111", --   61 - 0x3d  :  135 - 0x87
    "10010100", --   62 - 0x3e  :  148 - 0x94
    "10010101", --   63 - 0x3f  :  149 - 0x95
    "10000010", --   64 - 0x40  :  130 - 0x82 -- line 0x2
    "10000011", --   65 - 0x41  :  131 - 0x83
    "10000010", --   66 - 0x42  :  130 - 0x82
    "10000011", --   67 - 0x43  :  131 - 0x83
    "10000010", --   68 - 0x44  :  130 - 0x82
    "10010001", --   69 - 0x45  :  145 - 0x91
    "10010000", --   70 - 0x46  :  144 - 0x90
    "10000011", --   71 - 0x47  :  131 - 0x83
    "10000010", --   72 - 0x48  :  130 - 0x82
    "10010001", --   73 - 0x49  :  145 - 0x91
    "10010010", --   74 - 0x4a  :  146 - 0x92
    "10000011", --   75 - 0x4b  :  131 - 0x83
    "10000010", --   76 - 0x4c  :  130 - 0x82
    "10000011", --   77 - 0x4d  :  131 - 0x83
    "10000010", --   78 - 0x4e  :  130 - 0x82
    "10000001", --   79 - 0x4f  :  129 - 0x81
    "10000010", --   80 - 0x50  :  130 - 0x82
    "10000011", --   81 - 0x51  :  131 - 0x83
    "10000010", --   82 - 0x52  :  130 - 0x82
    "10000011", --   83 - 0x53  :  131 - 0x83
    "10000010", --   84 - 0x54  :  130 - 0x82
    "10000011", --   85 - 0x55  :  131 - 0x83
    "10000010", --   86 - 0x56  :  130 - 0x82
    "10000011", --   87 - 0x57  :  131 - 0x83
    "10000001", --   88 - 0x58  :  129 - 0x81
    "10000011", --   89 - 0x59  :  131 - 0x83
    "10010000", --   90 - 0x5a  :  144 - 0x90
    "10010011", --   91 - 0x5b  :  147 - 0x93
    "10000010", --   92 - 0x5c  :  130 - 0x82
    "10010000", --   93 - 0x5d  :  144 - 0x90
    "10010010", --   94 - 0x5e  :  146 - 0x92
    "10000011", --   95 - 0x5f  :  131 - 0x83
    "01001001", --   96 - 0x60  :   73 - 0x49 -- line 0x3
    "01001001", --   97 - 0x61  :   73 - 0x49
    "01001001", --   98 - 0x62  :   73 - 0x49
    "01001001", --   99 - 0x63  :   73 - 0x49
    "01001001", --  100 - 0x64  :   73 - 0x49
    "01001001", --  101 - 0x65  :   73 - 0x49
    "01001001", --  102 - 0x66  :   73 - 0x49
    "01001001", --  103 - 0x67  :   73 - 0x49
    "01001001", --  104 - 0x68  :   73 - 0x49
    "01001001", --  105 - 0x69  :   73 - 0x49
    "01001001", --  106 - 0x6a  :   73 - 0x49
    "01001001", --  107 - 0x6b  :   73 - 0x49
    "01001001", --  108 - 0x6c  :   73 - 0x49
    "01001001", --  109 - 0x6d  :   73 - 0x49
    "01001001", --  110 - 0x6e  :   73 - 0x49
    "01001001", --  111 - 0x6f  :   73 - 0x49
    "01001001", --  112 - 0x70  :   73 - 0x49
    "01001001", --  113 - 0x71  :   73 - 0x49
    "01001001", --  114 - 0x72  :   73 - 0x49
    "01001001", --  115 - 0x73  :   73 - 0x49
    "01001001", --  116 - 0x74  :   73 - 0x49
    "01001001", --  117 - 0x75  :   73 - 0x49
    "01001001", --  118 - 0x76  :   73 - 0x49
    "01001001", --  119 - 0x77  :   73 - 0x49
    "01001001", --  120 - 0x78  :   73 - 0x49
    "01001001", --  121 - 0x79  :   73 - 0x49
    "01001001", --  122 - 0x7a  :   73 - 0x49
    "01001001", --  123 - 0x7b  :   73 - 0x49
    "01001001", --  124 - 0x7c  :   73 - 0x49
    "01001001", --  125 - 0x7d  :   73 - 0x49
    "01001001", --  126 - 0x7e  :   73 - 0x49
    "01001001", --  127 - 0x7f  :   73 - 0x49
    "00000000", --  128 - 0x80  :    0 - 0x0 -- line 0x4
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000001", --  132 - 0x84  :    1 - 0x1
    "00000010", --  133 - 0x85  :    2 - 0x2
    "00000010", --  134 - 0x86  :    2 - 0x2
    "00000011", --  135 - 0x87  :    3 - 0x3
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000100", --  139 - 0x8b  :    4 - 0x4
    "00000010", --  140 - 0x8c  :    2 - 0x2
    "00000010", --  141 - 0x8d  :    2 - 0x2
    "00000010", --  142 - 0x8e  :    2 - 0x2
    "00000101", --  143 - 0x8f  :    5 - 0x5
    "00000001", --  144 - 0x90  :    1 - 0x1
    "00000010", --  145 - 0x91  :    2 - 0x2
    "00000010", --  146 - 0x92  :    2 - 0x2
    "00000110", --  147 - 0x93  :    6 - 0x6
    "00000010", --  148 - 0x94  :    2 - 0x2
    "00000010", --  149 - 0x95  :    2 - 0x2
    "00000110", --  150 - 0x96  :    6 - 0x6
    "00000010", --  151 - 0x97  :    2 - 0x2
    "00000010", --  152 - 0x98  :    2 - 0x2
    "00000111", --  153 - 0x99  :    7 - 0x7
    "00000010", --  154 - 0x9a  :    2 - 0x2
    "00000010", --  155 - 0x9b  :    2 - 0x2
    "00000011", --  156 - 0x9c  :    3 - 0x3
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- line 0x5
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00001000", --  164 - 0xa4  :    8 - 0x8
    "00001001", --  165 - 0xa5  :    9 - 0x9
    "00001001", --  166 - 0xa6  :    9 - 0x9
    "00001010", --  167 - 0xa7  :   10 - 0xa
    "00000000", --  168 - 0xa8  :    0 - 0x0
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00001011", --  170 - 0xaa  :   11 - 0xb
    "00001100", --  171 - 0xab  :   12 - 0xc
    "00001001", --  172 - 0xac  :    9 - 0x9
    "00001001", --  173 - 0xad  :    9 - 0x9
    "00001001", --  174 - 0xae  :    9 - 0x9
    "00001101", --  175 - 0xaf  :   13 - 0xd
    "00001110", --  176 - 0xb0  :   14 - 0xe
    "00001001", --  177 - 0xb1  :    9 - 0x9
    "00001001", --  178 - 0xb2  :    9 - 0x9
    "00001111", --  179 - 0xb3  :   15 - 0xf
    "00001001", --  180 - 0xb4  :    9 - 0x9
    "00001001", --  181 - 0xb5  :    9 - 0x9
    "00001111", --  182 - 0xb6  :   15 - 0xf
    "00001001", --  183 - 0xb7  :    9 - 0x9
    "00001001", --  184 - 0xb8  :    9 - 0x9
    "00010000", --  185 - 0xb9  :   16 - 0x10
    "00001001", --  186 - 0xba  :    9 - 0x9
    "00001001", --  187 - 0xbb  :    9 - 0x9
    "00001010", --  188 - 0xbc  :   10 - 0xa
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- line 0x6
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00001000", --  196 - 0xc4  :    8 - 0x8
    "00001001", --  197 - 0xc5  :    9 - 0x9
    "00001001", --  198 - 0xc6  :    9 - 0x9
    "00001010", --  199 - 0xc7  :   10 - 0xa
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00001000", --  202 - 0xca  :    8 - 0x8
    "00001001", --  203 - 0xcb  :    9 - 0x9
    "00001001", --  204 - 0xcc  :    9 - 0x9
    "00010001", --  205 - 0xcd  :   17 - 0x11
    "00001001", --  206 - 0xce  :    9 - 0x9
    "00001001", --  207 - 0xcf  :    9 - 0x9
    "00001111", --  208 - 0xd0  :   15 - 0xf
    "00001001", --  209 - 0xd1  :    9 - 0x9
    "00001001", --  210 - 0xd2  :    9 - 0x9
    "00001111", --  211 - 0xd3  :   15 - 0xf
    "00001001", --  212 - 0xd4  :    9 - 0x9
    "00001001", --  213 - 0xd5  :    9 - 0x9
    "00001111", --  214 - 0xd6  :   15 - 0xf
    "00001001", --  215 - 0xd7  :    9 - 0x9
    "00001001", --  216 - 0xd8  :    9 - 0x9
    "00010010", --  217 - 0xd9  :   18 - 0x12
    "00001001", --  218 - 0xda  :    9 - 0x9
    "00001001", --  219 - 0xdb  :    9 - 0x9
    "00001010", --  220 - 0xdc  :   10 - 0xa
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- line 0x7
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00001000", --  228 - 0xe4  :    8 - 0x8
    "00001001", --  229 - 0xe5  :    9 - 0x9
    "00001001", --  230 - 0xe6  :    9 - 0x9
    "00001010", --  231 - 0xe7  :   10 - 0xa
    "00000000", --  232 - 0xe8  :    0 - 0x0
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00001000", --  234 - 0xea  :    8 - 0x8
    "00001001", --  235 - 0xeb  :    9 - 0x9
    "00001001", --  236 - 0xec  :    9 - 0x9
    "00001111", --  237 - 0xed  :   15 - 0xf
    "00001001", --  238 - 0xee  :    9 - 0x9
    "00001001", --  239 - 0xef  :    9 - 0x9
    "00001111", --  240 - 0xf0  :   15 - 0xf
    "00001001", --  241 - 0xf1  :    9 - 0x9
    "00001001", --  242 - 0xf2  :    9 - 0x9
    "00010011", --  243 - 0xf3  :   19 - 0x13
    "00001001", --  244 - 0xf4  :    9 - 0x9
    "00001001", --  245 - 0xf5  :    9 - 0x9
    "00001111", --  246 - 0xf6  :   15 - 0xf
    "00001001", --  247 - 0xf7  :    9 - 0x9
    "00001001", --  248 - 0xf8  :    9 - 0x9
    "00010100", --  249 - 0xf9  :   20 - 0x14
    "00001001", --  250 - 0xfa  :    9 - 0x9
    "00001001", --  251 - 0xfb  :    9 - 0x9
    "00001010", --  252 - 0xfc  :   10 - 0xa
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- line 0x8
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00001000", --  260 - 0x104  :    8 - 0x8
    "00001001", --  261 - 0x105  :    9 - 0x9
    "00001001", --  262 - 0x106  :    9 - 0x9
    "00001010", --  263 - 0x107  :   10 - 0xa
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00001000", --  266 - 0x10a  :    8 - 0x8
    "00001001", --  267 - 0x10b  :    9 - 0x9
    "00001001", --  268 - 0x10c  :    9 - 0x9
    "00010101", --  269 - 0x10d  :   21 - 0x15
    "00001001", --  270 - 0x10e  :    9 - 0x9
    "00001001", --  271 - 0x10f  :    9 - 0x9
    "00001111", --  272 - 0x110  :   15 - 0xf
    "00001001", --  273 - 0x111  :    9 - 0x9
    "00001001", --  274 - 0x112  :    9 - 0x9
    "00010110", --  275 - 0x113  :   22 - 0x16
    "00001001", --  276 - 0x114  :    9 - 0x9
    "00001001", --  277 - 0x115  :    9 - 0x9
    "00001111", --  278 - 0x116  :   15 - 0xf
    "00001001", --  279 - 0x117  :    9 - 0x9
    "00001001", --  280 - 0x118  :    9 - 0x9
    "00010111", --  281 - 0x119  :   23 - 0x17
    "00001001", --  282 - 0x11a  :    9 - 0x9
    "00001001", --  283 - 0x11b  :    9 - 0x9
    "00001010", --  284 - 0x11c  :   10 - 0xa
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- line 0x9
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00001000", --  292 - 0x124  :    8 - 0x8
    "00001001", --  293 - 0x125  :    9 - 0x9
    "00001001", --  294 - 0x126  :    9 - 0x9
    "00011000", --  295 - 0x127  :   24 - 0x18
    "00000010", --  296 - 0x128  :    2 - 0x2
    "00000010", --  297 - 0x129  :    2 - 0x2
    "00011001", --  298 - 0x12a  :   25 - 0x19
    "00001001", --  299 - 0x12b  :    9 - 0x9
    "00001001", --  300 - 0x12c  :    9 - 0x9
    "00001001", --  301 - 0x12d  :    9 - 0x9
    "00001001", --  302 - 0x12e  :    9 - 0x9
    "00001001", --  303 - 0x12f  :    9 - 0x9
    "00001111", --  304 - 0x130  :   15 - 0xf
    "00001001", --  305 - 0x131  :    9 - 0x9
    "00001001", --  306 - 0x132  :    9 - 0x9
    "00011010", --  307 - 0x133  :   26 - 0x1a
    "00001001", --  308 - 0x134  :    9 - 0x9
    "00001001", --  309 - 0x135  :    9 - 0x9
    "00001111", --  310 - 0x136  :   15 - 0xf
    "00001001", --  311 - 0x137  :    9 - 0x9
    "00001001", --  312 - 0x138  :    9 - 0x9
    "00001111", --  313 - 0x139  :   15 - 0xf
    "00001001", --  314 - 0x13a  :    9 - 0x9
    "00001001", --  315 - 0x13b  :    9 - 0x9
    "00001010", --  316 - 0x13c  :   10 - 0xa
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- line 0xa
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00001000", --  324 - 0x144  :    8 - 0x8
    "00001001", --  325 - 0x145  :    9 - 0x9
    "00001001", --  326 - 0x146  :    9 - 0x9
    "00001001", --  327 - 0x147  :    9 - 0x9
    "00001001", --  328 - 0x148  :    9 - 0x9
    "00001001", --  329 - 0x149  :    9 - 0x9
    "00001111", --  330 - 0x14a  :   15 - 0xf
    "00001001", --  331 - 0x14b  :    9 - 0x9
    "00001001", --  332 - 0x14c  :    9 - 0x9
    "00011011", --  333 - 0x14d  :   27 - 0x1b
    "00001001", --  334 - 0x14e  :    9 - 0x9
    "00001001", --  335 - 0x14f  :    9 - 0x9
    "00001111", --  336 - 0x150  :   15 - 0xf
    "00001001", --  337 - 0x151  :    9 - 0x9
    "00011100", --  338 - 0x152  :   28 - 0x1c
    "00011101", --  339 - 0x153  :   29 - 0x1d
    "00011110", --  340 - 0x154  :   30 - 0x1e
    "00001001", --  341 - 0x155  :    9 - 0x9
    "00001111", --  342 - 0x156  :   15 - 0xf
    "00001001", --  343 - 0x157  :    9 - 0x9
    "00001001", --  344 - 0x158  :    9 - 0x9
    "00001111", --  345 - 0x159  :   15 - 0xf
    "00001001", --  346 - 0x15a  :    9 - 0x9
    "00001001", --  347 - 0x15b  :    9 - 0x9
    "00001010", --  348 - 0x15c  :   10 - 0xa
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- line 0xb
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00011111", --  356 - 0x164  :   31 - 0x1f
    "00100000", --  357 - 0x165  :   32 - 0x20
    "00100000", --  358 - 0x166  :   32 - 0x20
    "00100000", --  359 - 0x167  :   32 - 0x20
    "00100000", --  360 - 0x168  :   32 - 0x20
    "00100000", --  361 - 0x169  :   32 - 0x20
    "00100001", --  362 - 0x16a  :   33 - 0x21
    "00100000", --  363 - 0x16b  :   32 - 0x20
    "00100000", --  364 - 0x16c  :   32 - 0x20
    "00100001", --  365 - 0x16d  :   33 - 0x21
    "00100000", --  366 - 0x16e  :   32 - 0x20
    "00100000", --  367 - 0x16f  :   32 - 0x20
    "00100001", --  368 - 0x170  :   33 - 0x21
    "00100000", --  369 - 0x171  :   32 - 0x20
    "00100010", --  370 - 0x172  :   34 - 0x22
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00100011", --  372 - 0x174  :   35 - 0x23
    "00100000", --  373 - 0x175  :   32 - 0x20
    "00100001", --  374 - 0x176  :   33 - 0x21
    "00100000", --  375 - 0x177  :   32 - 0x20
    "00100000", --  376 - 0x178  :   32 - 0x20
    "00100001", --  377 - 0x179  :   33 - 0x21
    "00100000", --  378 - 0x17a  :   32 - 0x20
    "00100000", --  379 - 0x17b  :   32 - 0x20
    "00100100", --  380 - 0x17c  :   36 - 0x24
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- line 0xc
    "00000001", --  385 - 0x181  :    1 - 0x1
    "00000010", --  386 - 0x182  :    2 - 0x2
    "00100101", --  387 - 0x183  :   37 - 0x25
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00100110", --  389 - 0x185  :   38 - 0x26
    "00000010", --  390 - 0x186  :    2 - 0x2
    "00000011", --  391 - 0x187  :    3 - 0x3
    "00000100", --  392 - 0x188  :    4 - 0x4
    "00000010", --  393 - 0x189  :    2 - 0x2
    "00000010", --  394 - 0x18a  :    2 - 0x2
    "00000010", --  395 - 0x18b  :    2 - 0x2
    "00000101", --  396 - 0x18c  :    5 - 0x5
    "00000001", --  397 - 0x18d  :    1 - 0x1
    "00000010", --  398 - 0x18e  :    2 - 0x2
    "00000010", --  399 - 0x18f  :    2 - 0x2
    "00000110", --  400 - 0x190  :    6 - 0x6
    "00000010", --  401 - 0x191  :    2 - 0x2
    "00000010", --  402 - 0x192  :    2 - 0x2
    "00000110", --  403 - 0x193  :    6 - 0x6
    "00000010", --  404 - 0x194  :    2 - 0x2
    "00000010", --  405 - 0x195  :    2 - 0x2
    "00000010", --  406 - 0x196  :    2 - 0x2
    "00000010", --  407 - 0x197  :    2 - 0x2
    "00000010", --  408 - 0x198  :    2 - 0x2
    "00000110", --  409 - 0x199  :    6 - 0x6
    "00000010", --  410 - 0x19a  :    2 - 0x2
    "00000010", --  411 - 0x19b  :    2 - 0x2
    "00000010", --  412 - 0x19c  :    2 - 0x2
    "00000010", --  413 - 0x19d  :    2 - 0x2
    "00000101", --  414 - 0x19e  :    5 - 0x5
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- line 0xd
    "00001000", --  417 - 0x1a1  :    8 - 0x8
    "00001001", --  418 - 0x1a2  :    9 - 0x9
    "00100111", --  419 - 0x1a3  :   39 - 0x27
    "00101000", --  420 - 0x1a4  :   40 - 0x28
    "00101001", --  421 - 0x1a5  :   41 - 0x29
    "00001001", --  422 - 0x1a6  :    9 - 0x9
    "00101010", --  423 - 0x1a7  :   42 - 0x2a
    "00001100", --  424 - 0x1a8  :   12 - 0xc
    "00001001", --  425 - 0x1a9  :    9 - 0x9
    "00001001", --  426 - 0x1aa  :    9 - 0x9
    "00001001", --  427 - 0x1ab  :    9 - 0x9
    "00001101", --  428 - 0x1ac  :   13 - 0xd
    "00001110", --  429 - 0x1ad  :   14 - 0xe
    "00001001", --  430 - 0x1ae  :    9 - 0x9
    "00001001", --  431 - 0x1af  :    9 - 0x9
    "00001111", --  432 - 0x1b0  :   15 - 0xf
    "00001001", --  433 - 0x1b1  :    9 - 0x9
    "00001001", --  434 - 0x1b2  :    9 - 0x9
    "00001111", --  435 - 0x1b3  :   15 - 0xf
    "00001001", --  436 - 0x1b4  :    9 - 0x9
    "00001001", --  437 - 0x1b5  :    9 - 0x9
    "00001001", --  438 - 0x1b6  :    9 - 0x9
    "00001001", --  439 - 0x1b7  :    9 - 0x9
    "00001001", --  440 - 0x1b8  :    9 - 0x9
    "00001111", --  441 - 0x1b9  :   15 - 0xf
    "00001001", --  442 - 0x1ba  :    9 - 0x9
    "00001001", --  443 - 0x1bb  :    9 - 0x9
    "00001001", --  444 - 0x1bc  :    9 - 0x9
    "00001001", --  445 - 0x1bd  :    9 - 0x9
    "00001101", --  446 - 0x1be  :   13 - 0xd
    "00101011", --  447 - 0x1bf  :   43 - 0x2b
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- line 0xe
    "00001000", --  449 - 0x1c1  :    8 - 0x8
    "00001001", --  450 - 0x1c2  :    9 - 0x9
    "00001001", --  451 - 0x1c3  :    9 - 0x9
    "00101100", --  452 - 0x1c4  :   44 - 0x2c
    "00001001", --  453 - 0x1c5  :    9 - 0x9
    "00001001", --  454 - 0x1c6  :    9 - 0x9
    "00001111", --  455 - 0x1c7  :   15 - 0xf
    "00001001", --  456 - 0x1c8  :    9 - 0x9
    "00001001", --  457 - 0x1c9  :    9 - 0x9
    "00010001", --  458 - 0x1ca  :   17 - 0x11
    "00001001", --  459 - 0x1cb  :    9 - 0x9
    "00001001", --  460 - 0x1cc  :    9 - 0x9
    "00001111", --  461 - 0x1cd  :   15 - 0xf
    "00001001", --  462 - 0x1ce  :    9 - 0x9
    "00001001", --  463 - 0x1cf  :    9 - 0x9
    "00001111", --  464 - 0x1d0  :   15 - 0xf
    "00001001", --  465 - 0x1d1  :    9 - 0x9
    "00001001", --  466 - 0x1d2  :    9 - 0x9
    "00001111", --  467 - 0x1d3  :   15 - 0xf
    "00001001", --  468 - 0x1d4  :    9 - 0x9
    "00001001", --  469 - 0x1d5  :    9 - 0x9
    "00101101", --  470 - 0x1d6  :   45 - 0x2d
    "00100000", --  471 - 0x1d7  :   32 - 0x20
    "00100000", --  472 - 0x1d8  :   32 - 0x20
    "00101110", --  473 - 0x1d9  :   46 - 0x2e
    "00001001", --  474 - 0x1da  :    9 - 0x9
    "00001001", --  475 - 0x1db  :    9 - 0x9
    "00101111", --  476 - 0x1dc  :   47 - 0x2f
    "00001001", --  477 - 0x1dd  :    9 - 0x9
    "00001001", --  478 - 0x1de  :    9 - 0x9
    "00001010", --  479 - 0x1df  :   10 - 0xa
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- line 0xf
    "00001000", --  481 - 0x1e1  :    8 - 0x8
    "00001001", --  482 - 0x1e2  :    9 - 0x9
    "00001001", --  483 - 0x1e3  :    9 - 0x9
    "00110000", --  484 - 0x1e4  :   48 - 0x30
    "00001001", --  485 - 0x1e5  :    9 - 0x9
    "00001001", --  486 - 0x1e6  :    9 - 0x9
    "00001111", --  487 - 0x1e7  :   15 - 0xf
    "00001001", --  488 - 0x1e8  :    9 - 0x9
    "00001001", --  489 - 0x1e9  :    9 - 0x9
    "00001111", --  490 - 0x1ea  :   15 - 0xf
    "00001001", --  491 - 0x1eb  :    9 - 0x9
    "00001001", --  492 - 0x1ec  :    9 - 0x9
    "00001111", --  493 - 0x1ed  :   15 - 0xf
    "00001001", --  494 - 0x1ee  :    9 - 0x9
    "00001001", --  495 - 0x1ef  :    9 - 0x9
    "00010011", --  496 - 0x1f0  :   19 - 0x13
    "00001001", --  497 - 0x1f1  :    9 - 0x9
    "00001001", --  498 - 0x1f2  :    9 - 0x9
    "00001111", --  499 - 0x1f3  :   15 - 0xf
    "00001001", --  500 - 0x1f4  :    9 - 0x9
    "00001001", --  501 - 0x1f5  :    9 - 0x9
    "00110001", --  502 - 0x1f6  :   49 - 0x31
    "00110010", --  503 - 0x1f7  :   50 - 0x32
    "00110011", --  504 - 0x1f8  :   51 - 0x33
    "00001000", --  505 - 0x1f9  :    8 - 0x8
    "00001001", --  506 - 0x1fa  :    9 - 0x9
    "00001001", --  507 - 0x1fb  :    9 - 0x9
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "00001001", --  509 - 0x1fd  :    9 - 0x9
    "00001001", --  510 - 0x1fe  :    9 - 0x9
    "00001010", --  511 - 0x1ff  :   10 - 0xa
    "00000000", --  512 - 0x200  :    0 - 0x0 -- line 0x10
    "00001000", --  513 - 0x201  :    8 - 0x8
    "00001001", --  514 - 0x202  :    9 - 0x9
    "00001001", --  515 - 0x203  :    9 - 0x9
    "00110100", --  516 - 0x204  :   52 - 0x34
    "00001001", --  517 - 0x205  :    9 - 0x9
    "00001001", --  518 - 0x206  :    9 - 0x9
    "00001111", --  519 - 0x207  :   15 - 0xf
    "00001001", --  520 - 0x208  :    9 - 0x9
    "00001001", --  521 - 0x209  :    9 - 0x9
    "00001111", --  522 - 0x20a  :   15 - 0xf
    "00001001", --  523 - 0x20b  :    9 - 0x9
    "00001001", --  524 - 0x20c  :    9 - 0x9
    "00001111", --  525 - 0x20d  :   15 - 0xf
    "00001001", --  526 - 0x20e  :    9 - 0x9
    "00001001", --  527 - 0x20f  :    9 - 0x9
    "00010110", --  528 - 0x210  :   22 - 0x16
    "00001001", --  529 - 0x211  :    9 - 0x9
    "00001001", --  530 - 0x212  :    9 - 0x9
    "00001111", --  531 - 0x213  :   15 - 0xf
    "00001001", --  532 - 0x214  :    9 - 0x9
    "00001001", --  533 - 0x215  :    9 - 0x9
    "00110101", --  534 - 0x216  :   53 - 0x35
    "00110110", --  535 - 0x217  :   54 - 0x36
    "00110111", --  536 - 0x218  :   55 - 0x37
    "00001000", --  537 - 0x219  :    8 - 0x8
    "00001001", --  538 - 0x21a  :    9 - 0x9
    "00001001", --  539 - 0x21b  :    9 - 0x9
    "00111000", --  540 - 0x21c  :   56 - 0x38
    "00001001", --  541 - 0x21d  :    9 - 0x9
    "00111001", --  542 - 0x21e  :   57 - 0x39
    "00001010", --  543 - 0x21f  :   10 - 0xa
    "00000000", --  544 - 0x220  :    0 - 0x0 -- line 0x11
    "00001000", --  545 - 0x221  :    8 - 0x8
    "00001001", --  546 - 0x222  :    9 - 0x9
    "00001001", --  547 - 0x223  :    9 - 0x9
    "00001111", --  548 - 0x224  :   15 - 0xf
    "00001001", --  549 - 0x225  :    9 - 0x9
    "00001001", --  550 - 0x226  :    9 - 0x9
    "00001111", --  551 - 0x227  :   15 - 0xf
    "00001001", --  552 - 0x228  :    9 - 0x9
    "00001001", --  553 - 0x229  :    9 - 0x9
    "00111010", --  554 - 0x22a  :   58 - 0x3a
    "00001001", --  555 - 0x22b  :    9 - 0x9
    "00001001", --  556 - 0x22c  :    9 - 0x9
    "00001111", --  557 - 0x22d  :   15 - 0xf
    "00001001", --  558 - 0x22e  :    9 - 0x9
    "00001001", --  559 - 0x22f  :    9 - 0x9
    "00011010", --  560 - 0x230  :   26 - 0x1a
    "00001001", --  561 - 0x231  :    9 - 0x9
    "00001001", --  562 - 0x232  :    9 - 0x9
    "00001111", --  563 - 0x233  :   15 - 0xf
    "00001001", --  564 - 0x234  :    9 - 0x9
    "00001001", --  565 - 0x235  :    9 - 0x9
    "00111011", --  566 - 0x236  :   59 - 0x3b
    "00111100", --  567 - 0x237  :   60 - 0x3c
    "00111101", --  568 - 0x238  :   61 - 0x3d
    "00011001", --  569 - 0x239  :   25 - 0x19
    "00001001", --  570 - 0x23a  :    9 - 0x9
    "00001001", --  571 - 0x23b  :    9 - 0x9
    "00001001", --  572 - 0x23c  :    9 - 0x9
    "00001001", --  573 - 0x23d  :    9 - 0x9
    "00111110", --  574 - 0x23e  :   62 - 0x3e
    "00111111", --  575 - 0x23f  :   63 - 0x3f
    "00000000", --  576 - 0x240  :    0 - 0x0 -- line 0x12
    "00001000", --  577 - 0x241  :    8 - 0x8
    "00001001", --  578 - 0x242  :    9 - 0x9
    "00001001", --  579 - 0x243  :    9 - 0x9
    "00001111", --  580 - 0x244  :   15 - 0xf
    "00001001", --  581 - 0x245  :    9 - 0x9
    "00001001", --  582 - 0x246  :    9 - 0x9
    "01000000", --  583 - 0x247  :   64 - 0x40
    "01000001", --  584 - 0x248  :   65 - 0x41
    "00001001", --  585 - 0x249  :    9 - 0x9
    "00001001", --  586 - 0x24a  :    9 - 0x9
    "00001001", --  587 - 0x24b  :    9 - 0x9
    "01000010", --  588 - 0x24c  :   66 - 0x42
    "01000011", --  589 - 0x24d  :   67 - 0x43
    "00001001", --  590 - 0x24e  :    9 - 0x9
    "00011100", --  591 - 0x24f  :   28 - 0x1c
    "00011101", --  592 - 0x250  :   29 - 0x1d
    "00011110", --  593 - 0x251  :   30 - 0x1e
    "00001001", --  594 - 0x252  :    9 - 0x9
    "00001111", --  595 - 0x253  :   15 - 0xf
    "00001001", --  596 - 0x254  :    9 - 0x9
    "00001001", --  597 - 0x255  :    9 - 0x9
    "00001001", --  598 - 0x256  :    9 - 0x9
    "00001001", --  599 - 0x257  :    9 - 0x9
    "00001001", --  600 - 0x258  :    9 - 0x9
    "00001111", --  601 - 0x259  :   15 - 0xf
    "00001001", --  602 - 0x25a  :    9 - 0x9
    "00001001", --  603 - 0x25b  :    9 - 0x9
    "00101111", --  604 - 0x25c  :   47 - 0x2f
    "00001001", --  605 - 0x25d  :    9 - 0x9
    "01000100", --  606 - 0x25e  :   68 - 0x44
    "01000101", --  607 - 0x25f  :   69 - 0x45
    "00000000", --  608 - 0x260  :    0 - 0x0 -- line 0x13
    "00011111", --  609 - 0x261  :   31 - 0x1f
    "00100000", --  610 - 0x262  :   32 - 0x20
    "00100000", --  611 - 0x263  :   32 - 0x20
    "00100001", --  612 - 0x264  :   33 - 0x21
    "00100000", --  613 - 0x265  :   32 - 0x20
    "00100000", --  614 - 0x266  :   32 - 0x20
    "00100100", --  615 - 0x267  :   36 - 0x24
    "01000110", --  616 - 0x268  :   70 - 0x46
    "00100000", --  617 - 0x269  :   32 - 0x20
    "00100000", --  618 - 0x26a  :   32 - 0x20
    "00100000", --  619 - 0x26b  :   32 - 0x20
    "01000111", --  620 - 0x26c  :   71 - 0x47
    "01001000", --  621 - 0x26d  :   72 - 0x48
    "00100000", --  622 - 0x26e  :   32 - 0x20
    "00100010", --  623 - 0x26f  :   34 - 0x22
    "00000000", --  624 - 0x270  :    0 - 0x0
    "00100011", --  625 - 0x271  :   35 - 0x23
    "00100000", --  626 - 0x272  :   32 - 0x20
    "00100001", --  627 - 0x273  :   33 - 0x21
    "00100000", --  628 - 0x274  :   32 - 0x20
    "00100000", --  629 - 0x275  :   32 - 0x20
    "00100000", --  630 - 0x276  :   32 - 0x20
    "00100000", --  631 - 0x277  :   32 - 0x20
    "00100000", --  632 - 0x278  :   32 - 0x20
    "00100001", --  633 - 0x279  :   33 - 0x21
    "00100000", --  634 - 0x27a  :   32 - 0x20
    "00100000", --  635 - 0x27b  :   32 - 0x20
    "00100001", --  636 - 0x27c  :   33 - 0x21
    "00100000", --  637 - 0x27d  :   32 - 0x20
    "00100000", --  638 - 0x27e  :   32 - 0x20
    "00100100", --  639 - 0x27f  :   36 - 0x24
    "00000000", --  640 - 0x280  :    0 - 0x0 -- line 0x14
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- line 0x15
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "01010000", --  683 - 0x2ab  :   80 - 0x50
    "01010001", --  684 - 0x2ac  :   81 - 0x51
    "01010010", --  685 - 0x2ad  :   82 - 0x52
    "01010011", --  686 - 0x2ae  :   83 - 0x53
    "01010011", --  687 - 0x2af  :   83 - 0x53
    "00000000", --  688 - 0x2b0  :    0 - 0x0
    "01010011", --  689 - 0x2b1  :   83 - 0x53
    "01010100", --  690 - 0x2b2  :   84 - 0x54
    "01010101", --  691 - 0x2b3  :   85 - 0x55
    "01010001", --  692 - 0x2b4  :   81 - 0x51
    "01010100", --  693 - 0x2b5  :   84 - 0x54
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- line 0x16
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "01100000", --  715 - 0x2cb  :   96 - 0x60
    "01100001", --  716 - 0x2cc  :   97 - 0x61
    "01100010", --  717 - 0x2cd  :   98 - 0x62
    "01100011", --  718 - 0x2ce  :   99 - 0x63
    "01100011", --  719 - 0x2cf  :   99 - 0x63
    "00000000", --  720 - 0x2d0  :    0 - 0x0
    "01100011", --  721 - 0x2d1  :   99 - 0x63
    "01100100", --  722 - 0x2d2  :  100 - 0x64
    "01100101", --  723 - 0x2d3  :  101 - 0x65
    "01100001", --  724 - 0x2d4  :   97 - 0x61
    "01100100", --  725 - 0x2d5  :  100 - 0x64
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- line 0x17
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- line 0x18
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "10010010", --  800 - 0x320  :  146 - 0x92 -- line 0x19
    "10010011", --  801 - 0x321  :  147 - 0x93
    "10010010", --  802 - 0x322  :  146 - 0x92
    "10000011", --  803 - 0x323  :  131 - 0x83
    "10010010", --  804 - 0x324  :  146 - 0x92
    "10010011", --  805 - 0x325  :  147 - 0x93
    "10000010", --  806 - 0x326  :  130 - 0x82
    "10010011", --  807 - 0x327  :  147 - 0x93
    "10010010", --  808 - 0x328  :  146 - 0x92
    "10010010", --  809 - 0x329  :  146 - 0x92
    "10010011", --  810 - 0x32a  :  147 - 0x93
    "10010000", --  811 - 0x32b  :  144 - 0x90
    "10010010", --  812 - 0x32c  :  146 - 0x92
    "10000010", --  813 - 0x32d  :  130 - 0x82
    "10010000", --  814 - 0x32e  :  144 - 0x90
    "10010011", --  815 - 0x32f  :  147 - 0x93
    "10010010", --  816 - 0x330  :  146 - 0x92
    "10010011", --  817 - 0x331  :  147 - 0x93
    "10000011", --  818 - 0x332  :  131 - 0x83
    "10010011", --  819 - 0x333  :  147 - 0x93
    "10010011", --  820 - 0x334  :  147 - 0x93
    "10010000", --  821 - 0x335  :  144 - 0x90
    "10010010", --  822 - 0x336  :  146 - 0x92
    "10010011", --  823 - 0x337  :  147 - 0x93
    "10010010", --  824 - 0x338  :  146 - 0x92
    "01001010", --  825 - 0x339  :   74 - 0x4a
    "01001011", --  826 - 0x33a  :   75 - 0x4b
    "01001100", --  827 - 0x33b  :   76 - 0x4c
    "01001101", --  828 - 0x33c  :   77 - 0x4d
    "01001110", --  829 - 0x33d  :   78 - 0x4e
    "01001111", --  830 - 0x33e  :   79 - 0x4f
    "10010010", --  831 - 0x33f  :  146 - 0x92
    "10000100", --  832 - 0x340  :  132 - 0x84 -- line 0x1a
    "10000101", --  833 - 0x341  :  133 - 0x85
    "10000100", --  834 - 0x342  :  132 - 0x84
    "10000101", --  835 - 0x343  :  133 - 0x85
    "10000100", --  836 - 0x344  :  132 - 0x84
    "10000101", --  837 - 0x345  :  133 - 0x85
    "10000100", --  838 - 0x346  :  132 - 0x84
    "10000101", --  839 - 0x347  :  133 - 0x85
    "10000100", --  840 - 0x348  :  132 - 0x84
    "10000101", --  841 - 0x349  :  133 - 0x85
    "10000100", --  842 - 0x34a  :  132 - 0x84
    "10000101", --  843 - 0x34b  :  133 - 0x85
    "10000100", --  844 - 0x34c  :  132 - 0x84
    "10000101", --  845 - 0x34d  :  133 - 0x85
    "10000100", --  846 - 0x34e  :  132 - 0x84
    "10000101", --  847 - 0x34f  :  133 - 0x85
    "10000100", --  848 - 0x350  :  132 - 0x84
    "10000101", --  849 - 0x351  :  133 - 0x85
    "10000100", --  850 - 0x352  :  132 - 0x84
    "10000101", --  851 - 0x353  :  133 - 0x85
    "10000100", --  852 - 0x354  :  132 - 0x84
    "10000101", --  853 - 0x355  :  133 - 0x85
    "10000100", --  854 - 0x356  :  132 - 0x84
    "10000101", --  855 - 0x357  :  133 - 0x85
    "10000100", --  856 - 0x358  :  132 - 0x84
    "10000101", --  857 - 0x359  :  133 - 0x85
    "10000100", --  858 - 0x35a  :  132 - 0x84
    "10000101", --  859 - 0x35b  :  133 - 0x85
    "10000100", --  860 - 0x35c  :  132 - 0x84
    "10000101", --  861 - 0x35d  :  133 - 0x85
    "10000100", --  862 - 0x35e  :  132 - 0x84
    "10000101", --  863 - 0x35f  :  133 - 0x85
    "10010100", --  864 - 0x360  :  148 - 0x94 -- line 0x1b
    "10010111", --  865 - 0x361  :  151 - 0x97
    "10010100", --  866 - 0x362  :  148 - 0x94
    "10010101", --  867 - 0x363  :  149 - 0x95
    "10010100", --  868 - 0x364  :  148 - 0x94
    "10000111", --  869 - 0x365  :  135 - 0x87
    "10010111", --  870 - 0x366  :  151 - 0x97
    "10010111", --  871 - 0x367  :  151 - 0x97
    "10010100", --  872 - 0x368  :  148 - 0x94
    "10000110", --  873 - 0x369  :  134 - 0x86
    "10010100", --  874 - 0x36a  :  148 - 0x94
    "10010101", --  875 - 0x36b  :  149 - 0x95
    "10010110", --  876 - 0x36c  :  150 - 0x96
    "10010101", --  877 - 0x36d  :  149 - 0x95
    "10010100", --  878 - 0x36e  :  148 - 0x94
    "10010101", --  879 - 0x36f  :  149 - 0x95
    "10000111", --  880 - 0x370  :  135 - 0x87
    "10010111", --  881 - 0x371  :  151 - 0x97
    "10010100", --  882 - 0x372  :  148 - 0x94
    "10000111", --  883 - 0x373  :  135 - 0x87
    "10010110", --  884 - 0x374  :  150 - 0x96
    "10000110", --  885 - 0x375  :  134 - 0x86
    "10010100", --  886 - 0x376  :  148 - 0x94
    "10010101", --  887 - 0x377  :  149 - 0x95
    "10000111", --  888 - 0x378  :  135 - 0x87
    "10010101", --  889 - 0x379  :  149 - 0x95
    "10010100", --  890 - 0x37a  :  148 - 0x94
    "10010111", --  891 - 0x37b  :  151 - 0x97
    "10010100", --  892 - 0x37c  :  148 - 0x94
    "10000110", --  893 - 0x37d  :  134 - 0x86
    "10010100", --  894 - 0x37e  :  148 - 0x94
    "10010101", --  895 - 0x37f  :  149 - 0x95
    "10000100", --  896 - 0x380  :  132 - 0x84 -- line 0x1c
    "10000101", --  897 - 0x381  :  133 - 0x85
    "10010110", --  898 - 0x382  :  150 - 0x96
    "10000101", --  899 - 0x383  :  133 - 0x85
    "10000111", --  900 - 0x384  :  135 - 0x87
    "10010111", --  901 - 0x385  :  151 - 0x97
    "10000100", --  902 - 0x386  :  132 - 0x84
    "10000101", --  903 - 0x387  :  133 - 0x85
    "10000100", --  904 - 0x388  :  132 - 0x84
    "10000101", --  905 - 0x389  :  133 - 0x85
    "10000100", --  906 - 0x38a  :  132 - 0x84
    "10000111", --  907 - 0x38b  :  135 - 0x87
    "10000100", --  908 - 0x38c  :  132 - 0x84
    "10000110", --  909 - 0x38d  :  134 - 0x86
    "10000100", --  910 - 0x38e  :  132 - 0x84
    "10000101", --  911 - 0x38f  :  133 - 0x85
    "10000100", --  912 - 0x390  :  132 - 0x84
    "10000101", --  913 - 0x391  :  133 - 0x85
    "10000100", --  914 - 0x392  :  132 - 0x84
    "10000101", --  915 - 0x393  :  133 - 0x85
    "10000100", --  916 - 0x394  :  132 - 0x84
    "10000101", --  917 - 0x395  :  133 - 0x85
    "10010111", --  918 - 0x396  :  151 - 0x97
    "10000101", --  919 - 0x397  :  133 - 0x85
    "10000100", --  920 - 0x398  :  132 - 0x84
    "10010111", --  921 - 0x399  :  151 - 0x97
    "10000111", --  922 - 0x39a  :  135 - 0x87
    "10000101", --  923 - 0x39b  :  133 - 0x85
    "10000110", --  924 - 0x39c  :  134 - 0x86
    "10000111", --  925 - 0x39d  :  135 - 0x87
    "10000100", --  926 - 0x39e  :  132 - 0x84
    "10000101", --  927 - 0x39f  :  133 - 0x85
    "10010100", --  928 - 0x3a0  :  148 - 0x94 -- line 0x1d
    "10010101", --  929 - 0x3a1  :  149 - 0x95
    "10010100", --  930 - 0x3a2  :  148 - 0x94
    "10010101", --  931 - 0x3a3  :  149 - 0x95
    "10010100", --  932 - 0x3a4  :  148 - 0x94
    "10000110", --  933 - 0x3a5  :  134 - 0x86
    "10010100", --  934 - 0x3a6  :  148 - 0x94
    "10010101", --  935 - 0x3a7  :  149 - 0x95
    "10010100", --  936 - 0x3a8  :  148 - 0x94
    "10010101", --  937 - 0x3a9  :  149 - 0x95
    "10010100", --  938 - 0x3aa  :  148 - 0x94
    "10010101", --  939 - 0x3ab  :  149 - 0x95
    "10010100", --  940 - 0x3ac  :  148 - 0x94
    "10010111", --  941 - 0x3ad  :  151 - 0x97
    "10010110", --  942 - 0x3ae  :  150 - 0x96
    "10010101", --  943 - 0x3af  :  149 - 0x95
    "10010100", --  944 - 0x3b0  :  148 - 0x94
    "10010101", --  945 - 0x3b1  :  149 - 0x95
    "10010100", --  946 - 0x3b2  :  148 - 0x94
    "10010101", --  947 - 0x3b3  :  149 - 0x95
    "10010100", --  948 - 0x3b4  :  148 - 0x94
    "10010101", --  949 - 0x3b5  :  149 - 0x95
    "10010100", --  950 - 0x3b6  :  148 - 0x94
    "10010101", --  951 - 0x3b7  :  149 - 0x95
    "10000110", --  952 - 0x3b8  :  134 - 0x86
    "10010101", --  953 - 0x3b9  :  149 - 0x95
    "10010100", --  954 - 0x3ba  :  148 - 0x94
    "10010101", --  955 - 0x3bb  :  149 - 0x95
    "10010100", --  956 - 0x3bc  :  148 - 0x94
    "10010101", --  957 - 0x3bd  :  149 - 0x95
    "10010100", --  958 - 0x3be  :  148 - 0x94
    "10010101", --  959 - 0x3bf  :  149 - 0x95
        ---- Attribute Table 0----
    "10101010", --  960 - 0x3c0  :  170 - 0xaa
    "10101010", --  961 - 0x3c1  :  170 - 0xaa
    "10101010", --  962 - 0x3c2  :  170 - 0xaa
    "10101010", --  963 - 0x3c3  :  170 - 0xaa
    "10101010", --  964 - 0x3c4  :  170 - 0xaa
    "10101010", --  965 - 0x3c5  :  170 - 0xaa
    "10101010", --  966 - 0x3c6  :  170 - 0xaa
    "10101010", --  967 - 0x3c7  :  170 - 0xaa
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "01010101", --  990 - 0x3de  :   85 - 0x55
    "01010101", --  991 - 0x3df  :   85 - 0x55
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "01010101", --  997 - 0x3e5  :   85 - 0x55
    "01010101", --  998 - 0x3e6  :   85 - 0x55
    "01010101", --  999 - 0x3e7  :   85 - 0x55
    "00000101", -- 1000 - 0x3e8  :    5 - 0x5
    "10000101", -- 1001 - 0x3e9  :  133 - 0x85
    "11101101", -- 1002 - 0x3ea  :  237 - 0xed
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111111", -- 1004 - 0x3ec  :  255 - 0xff
    "00110111", -- 1005 - 0x3ed  :   55 - 0x37
    "00000101", -- 1006 - 0x3ee  :    5 - 0x5
    "00000101", -- 1007 - 0x3ef  :    5 - 0x5
    "10101010", -- 1008 - 0x3f0  :  170 - 0xaa
    "10101010", -- 1009 - 0x3f1  :  170 - 0xaa
    "10101010", -- 1010 - 0x3f2  :  170 - 0xaa
    "10101010", -- 1011 - 0x3f3  :  170 - 0xaa
    "10101010", -- 1012 - 0x3f4  :  170 - 0xaa
    "10101010", -- 1013 - 0x3f5  :  170 - 0xaa
    "10101010", -- 1014 - 0x3f6  :  170 - 0xaa
    "10101010", -- 1015 - 0x3f7  :  170 - 0xaa
    "00001010", -- 1016 - 0x3f8  :   10 - 0xa
    "00001010", -- 1017 - 0x3f9  :   10 - 0xa
    "00001010", -- 1018 - 0x3fa  :   10 - 0xa
    "00001010", -- 1019 - 0x3fb  :   10 - 0xa
    "00001010", -- 1020 - 0x3fc  :   10 - 0xa
    "00001010", -- 1021 - 0x3fd  :   10 - 0xa
    "00001010", -- 1022 - 0x3fe  :   10 - 0xa
    "00001010"  -- 1023 - 0x3ff  :   10 - 0xa
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
