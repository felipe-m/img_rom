//-   Background Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_traspas_patron.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_MARIO_TRASPAS_BG
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table both color planes
      12'h0: dout  = 8'b00111000; //    0 :  56 - 0x38 -- Background 0x0
      12'h1: dout  = 8'b01001100; //    1 :  76 - 0x4c
      12'h2: dout  = 8'b11000110; //    2 : 198 - 0xc6
      12'h3: dout  = 8'b11000110; //    3 : 198 - 0xc6
      12'h4: dout  = 8'b11000110; //    4 : 198 - 0xc6
      12'h5: dout  = 8'b01100100; //    5 : 100 - 0x64
      12'h6: dout  = 8'b00111000; //    6 :  56 - 0x38
      12'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout  = 8'b00011000; //   16 :  24 - 0x18 -- Background 0x1
      12'h11: dout  = 8'b00111000; //   17 :  56 - 0x38
      12'h12: dout  = 8'b00011000; //   18 :  24 - 0x18
      12'h13: dout  = 8'b00011000; //   19 :  24 - 0x18
      12'h14: dout  = 8'b00011000; //   20 :  24 - 0x18
      12'h15: dout  = 8'b00011000; //   21 :  24 - 0x18
      12'h16: dout  = 8'b01111110; //   22 : 126 - 0x7e
      12'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout  = 8'b01111100; //   32 : 124 - 0x7c -- Background 0x2
      12'h21: dout  = 8'b11000110; //   33 : 198 - 0xc6
      12'h22: dout  = 8'b00001110; //   34 :  14 - 0xe
      12'h23: dout  = 8'b00111100; //   35 :  60 - 0x3c
      12'h24: dout  = 8'b01111000; //   36 : 120 - 0x78
      12'h25: dout  = 8'b11100000; //   37 : 224 - 0xe0
      12'h26: dout  = 8'b11111110; //   38 : 254 - 0xfe
      12'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout  = 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout  = 8'b01111110; //   48 : 126 - 0x7e -- Background 0x3
      12'h31: dout  = 8'b00001100; //   49 :  12 - 0xc
      12'h32: dout  = 8'b00011000; //   50 :  24 - 0x18
      12'h33: dout  = 8'b00111100; //   51 :  60 - 0x3c
      12'h34: dout  = 8'b00000110; //   52 :   6 - 0x6
      12'h35: dout  = 8'b11000110; //   53 : 198 - 0xc6
      12'h36: dout  = 8'b01111100; //   54 : 124 - 0x7c
      12'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout  = 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00011100; //   64 :  28 - 0x1c -- Background 0x4
      12'h41: dout  = 8'b00111100; //   65 :  60 - 0x3c
      12'h42: dout  = 8'b01101100; //   66 : 108 - 0x6c
      12'h43: dout  = 8'b11001100; //   67 : 204 - 0xcc
      12'h44: dout  = 8'b11111110; //   68 : 254 - 0xfe
      12'h45: dout  = 8'b00001100; //   69 :  12 - 0xc
      12'h46: dout  = 8'b00001100; //   70 :  12 - 0xc
      12'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- plane 1
      12'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout  = 8'b11111100; //   80 : 252 - 0xfc -- Background 0x5
      12'h51: dout  = 8'b11000000; //   81 : 192 - 0xc0
      12'h52: dout  = 8'b11111100; //   82 : 252 - 0xfc
      12'h53: dout  = 8'b00000110; //   83 :   6 - 0x6
      12'h54: dout  = 8'b00000110; //   84 :   6 - 0x6
      12'h55: dout  = 8'b11000110; //   85 : 198 - 0xc6
      12'h56: dout  = 8'b01111100; //   86 : 124 - 0x7c
      12'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- plane 1
      12'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout  = 8'b00111100; //   96 :  60 - 0x3c -- Background 0x6
      12'h61: dout  = 8'b01100000; //   97 :  96 - 0x60
      12'h62: dout  = 8'b11000000; //   98 : 192 - 0xc0
      12'h63: dout  = 8'b11111100; //   99 : 252 - 0xfc
      12'h64: dout  = 8'b11000110; //  100 : 198 - 0xc6
      12'h65: dout  = 8'b11000110; //  101 : 198 - 0xc6
      12'h66: dout  = 8'b01111100; //  102 : 124 - 0x7c
      12'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout  = 8'b00000000; //  104 :   0 - 0x0 -- plane 1
      12'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout  = 8'b11111110; //  112 : 254 - 0xfe -- Background 0x7
      12'h71: dout  = 8'b11000110; //  113 : 198 - 0xc6
      12'h72: dout  = 8'b00001100; //  114 :  12 - 0xc
      12'h73: dout  = 8'b00011000; //  115 :  24 - 0x18
      12'h74: dout  = 8'b00110000; //  116 :  48 - 0x30
      12'h75: dout  = 8'b00110000; //  117 :  48 - 0x30
      12'h76: dout  = 8'b00110000; //  118 :  48 - 0x30
      12'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- plane 1
      12'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout  = 8'b01111100; //  128 : 124 - 0x7c -- Background 0x8
      12'h81: dout  = 8'b11000110; //  129 : 198 - 0xc6
      12'h82: dout  = 8'b11000110; //  130 : 198 - 0xc6
      12'h83: dout  = 8'b01111100; //  131 : 124 - 0x7c
      12'h84: dout  = 8'b11000110; //  132 : 198 - 0xc6
      12'h85: dout  = 8'b11000110; //  133 : 198 - 0xc6
      12'h86: dout  = 8'b01111100; //  134 : 124 - 0x7c
      12'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout  = 8'b01111100; //  144 : 124 - 0x7c -- Background 0x9
      12'h91: dout  = 8'b11000110; //  145 : 198 - 0xc6
      12'h92: dout  = 8'b11000110; //  146 : 198 - 0xc6
      12'h93: dout  = 8'b01111110; //  147 : 126 - 0x7e
      12'h94: dout  = 8'b00000110; //  148 :   6 - 0x6
      12'h95: dout  = 8'b00001100; //  149 :  12 - 0xc
      12'h96: dout  = 8'b01111000; //  150 : 120 - 0x78
      12'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- plane 1
      12'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout  = 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout  = 8'b00111000; //  160 :  56 - 0x38 -- Background 0xa
      12'hA1: dout  = 8'b01101100; //  161 : 108 - 0x6c
      12'hA2: dout  = 8'b11000110; //  162 : 198 - 0xc6
      12'hA3: dout  = 8'b11000110; //  163 : 198 - 0xc6
      12'hA4: dout  = 8'b11111110; //  164 : 254 - 0xfe
      12'hA5: dout  = 8'b11000110; //  165 : 198 - 0xc6
      12'hA6: dout  = 8'b11000110; //  166 : 198 - 0xc6
      12'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout  = 8'b00000000; //  168 :   0 - 0x0 -- plane 1
      12'hA9: dout  = 8'b00000000; //  169 :   0 - 0x0
      12'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout  = 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout  = 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout  = 8'b11111100; //  176 : 252 - 0xfc -- Background 0xb
      12'hB1: dout  = 8'b11000110; //  177 : 198 - 0xc6
      12'hB2: dout  = 8'b11000110; //  178 : 198 - 0xc6
      12'hB3: dout  = 8'b11111100; //  179 : 252 - 0xfc
      12'hB4: dout  = 8'b11000110; //  180 : 198 - 0xc6
      12'hB5: dout  = 8'b11000110; //  181 : 198 - 0xc6
      12'hB6: dout  = 8'b11111100; //  182 : 252 - 0xfc
      12'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout  = 8'b00000000; //  184 :   0 - 0x0 -- plane 1
      12'hB9: dout  = 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout  = 8'b00000000; //  186 :   0 - 0x0
      12'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout  = 8'b00000000; //  188 :   0 - 0x0
      12'hBD: dout  = 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout  = 8'b00111100; //  192 :  60 - 0x3c -- Background 0xc
      12'hC1: dout  = 8'b01100110; //  193 : 102 - 0x66
      12'hC2: dout  = 8'b11000000; //  194 : 192 - 0xc0
      12'hC3: dout  = 8'b11000000; //  195 : 192 - 0xc0
      12'hC4: dout  = 8'b11000000; //  196 : 192 - 0xc0
      12'hC5: dout  = 8'b01100110; //  197 : 102 - 0x66
      12'hC6: dout  = 8'b00111100; //  198 :  60 - 0x3c
      12'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- plane 1
      12'hC9: dout  = 8'b00000000; //  201 :   0 - 0x0
      12'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout  = 8'b00000000; //  204 :   0 - 0x0
      12'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout  = 8'b11111000; //  208 : 248 - 0xf8 -- Background 0xd
      12'hD1: dout  = 8'b11001100; //  209 : 204 - 0xcc
      12'hD2: dout  = 8'b11000110; //  210 : 198 - 0xc6
      12'hD3: dout  = 8'b11000110; //  211 : 198 - 0xc6
      12'hD4: dout  = 8'b11000110; //  212 : 198 - 0xc6
      12'hD5: dout  = 8'b11001100; //  213 : 204 - 0xcc
      12'hD6: dout  = 8'b11111000; //  214 : 248 - 0xf8
      12'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- plane 1
      12'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout  = 8'b00000000; //  219 :   0 - 0x0
      12'hDC: dout  = 8'b00000000; //  220 :   0 - 0x0
      12'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout  = 8'b11111110; //  224 : 254 - 0xfe -- Background 0xe
      12'hE1: dout  = 8'b11000000; //  225 : 192 - 0xc0
      12'hE2: dout  = 8'b11000000; //  226 : 192 - 0xc0
      12'hE3: dout  = 8'b11111100; //  227 : 252 - 0xfc
      12'hE4: dout  = 8'b11000000; //  228 : 192 - 0xc0
      12'hE5: dout  = 8'b11000000; //  229 : 192 - 0xc0
      12'hE6: dout  = 8'b11111110; //  230 : 254 - 0xfe
      12'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0 -- plane 1
      12'hE9: dout  = 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout  = 8'b00000000; //  234 :   0 - 0x0
      12'hEB: dout  = 8'b00000000; //  235 :   0 - 0x0
      12'hEC: dout  = 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout  = 8'b11111110; //  240 : 254 - 0xfe -- Background 0xf
      12'hF1: dout  = 8'b11000000; //  241 : 192 - 0xc0
      12'hF2: dout  = 8'b11000000; //  242 : 192 - 0xc0
      12'hF3: dout  = 8'b11111100; //  243 : 252 - 0xfc
      12'hF4: dout  = 8'b11000000; //  244 : 192 - 0xc0
      12'hF5: dout  = 8'b11000000; //  245 : 192 - 0xc0
      12'hF6: dout  = 8'b11000000; //  246 : 192 - 0xc0
      12'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout  = 8'b00111110; //  256 :  62 - 0x3e -- Background 0x10
      12'h101: dout  = 8'b01100000; //  257 :  96 - 0x60
      12'h102: dout  = 8'b11000000; //  258 : 192 - 0xc0
      12'h103: dout  = 8'b11001110; //  259 : 206 - 0xce
      12'h104: dout  = 8'b11000110; //  260 : 198 - 0xc6
      12'h105: dout  = 8'b01100110; //  261 : 102 - 0x66
      12'h106: dout  = 8'b00111110; //  262 :  62 - 0x3e
      12'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout  = 8'b11000110; //  272 : 198 - 0xc6 -- Background 0x11
      12'h111: dout  = 8'b11000110; //  273 : 198 - 0xc6
      12'h112: dout  = 8'b11000110; //  274 : 198 - 0xc6
      12'h113: dout  = 8'b11111110; //  275 : 254 - 0xfe
      12'h114: dout  = 8'b11000110; //  276 : 198 - 0xc6
      12'h115: dout  = 8'b11000110; //  277 : 198 - 0xc6
      12'h116: dout  = 8'b11000110; //  278 : 198 - 0xc6
      12'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout  = 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout  = 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout  = 8'b00000000; //  283 :   0 - 0x0
      12'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout  = 8'b00000000; //  285 :   0 - 0x0
      12'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout  = 8'b01111110; //  288 : 126 - 0x7e -- Background 0x12
      12'h121: dout  = 8'b00011000; //  289 :  24 - 0x18
      12'h122: dout  = 8'b00011000; //  290 :  24 - 0x18
      12'h123: dout  = 8'b00011000; //  291 :  24 - 0x18
      12'h124: dout  = 8'b00011000; //  292 :  24 - 0x18
      12'h125: dout  = 8'b00011000; //  293 :  24 - 0x18
      12'h126: dout  = 8'b01111110; //  294 : 126 - 0x7e
      12'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout  = 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout  = 8'b00000000; //  297 :   0 - 0x0
      12'h12A: dout  = 8'b00000000; //  298 :   0 - 0x0
      12'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout  = 8'b00011110; //  304 :  30 - 0x1e -- Background 0x13
      12'h131: dout  = 8'b00000110; //  305 :   6 - 0x6
      12'h132: dout  = 8'b00000110; //  306 :   6 - 0x6
      12'h133: dout  = 8'b00000110; //  307 :   6 - 0x6
      12'h134: dout  = 8'b11000110; //  308 : 198 - 0xc6
      12'h135: dout  = 8'b11000110; //  309 : 198 - 0xc6
      12'h136: dout  = 8'b01111100; //  310 : 124 - 0x7c
      12'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      12'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- plane 1
      12'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b11000110; //  320 : 198 - 0xc6 -- Background 0x14
      12'h141: dout  = 8'b11001100; //  321 : 204 - 0xcc
      12'h142: dout  = 8'b11011000; //  322 : 216 - 0xd8
      12'h143: dout  = 8'b11110000; //  323 : 240 - 0xf0
      12'h144: dout  = 8'b11111000; //  324 : 248 - 0xf8
      12'h145: dout  = 8'b11011100; //  325 : 220 - 0xdc
      12'h146: dout  = 8'b11001110; //  326 : 206 - 0xce
      12'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      12'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- plane 1
      12'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout  = 8'b00000000; //  330 :   0 - 0x0
      12'h14B: dout  = 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout  = 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout  = 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout  = 8'b01100000; //  336 :  96 - 0x60 -- Background 0x15
      12'h151: dout  = 8'b01100000; //  337 :  96 - 0x60
      12'h152: dout  = 8'b01100000; //  338 :  96 - 0x60
      12'h153: dout  = 8'b01100000; //  339 :  96 - 0x60
      12'h154: dout  = 8'b01100000; //  340 :  96 - 0x60
      12'h155: dout  = 8'b01100000; //  341 :  96 - 0x60
      12'h156: dout  = 8'b01111110; //  342 : 126 - 0x7e
      12'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout  = 8'b00000000; //  344 :   0 - 0x0 -- plane 1
      12'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout  = 8'b11000110; //  352 : 198 - 0xc6 -- Background 0x16
      12'h161: dout  = 8'b11101110; //  353 : 238 - 0xee
      12'h162: dout  = 8'b11111110; //  354 : 254 - 0xfe
      12'h163: dout  = 8'b11111110; //  355 : 254 - 0xfe
      12'h164: dout  = 8'b11010110; //  356 : 214 - 0xd6
      12'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      12'h166: dout  = 8'b11000110; //  358 : 198 - 0xc6
      12'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- plane 1
      12'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout  = 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout  = 8'b11000110; //  368 : 198 - 0xc6 -- Background 0x17
      12'h171: dout  = 8'b11100110; //  369 : 230 - 0xe6
      12'h172: dout  = 8'b11110110; //  370 : 246 - 0xf6
      12'h173: dout  = 8'b11111110; //  371 : 254 - 0xfe
      12'h174: dout  = 8'b11011110; //  372 : 222 - 0xde
      12'h175: dout  = 8'b11001110; //  373 : 206 - 0xce
      12'h176: dout  = 8'b11000110; //  374 : 198 - 0xc6
      12'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout  = 8'b00000000; //  376 :   0 - 0x0 -- plane 1
      12'h179: dout  = 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout  = 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout  = 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout  = 8'b00000000; //  380 :   0 - 0x0
      12'h17D: dout  = 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout  = 8'b01111100; //  384 : 124 - 0x7c -- Background 0x18
      12'h181: dout  = 8'b11000110; //  385 : 198 - 0xc6
      12'h182: dout  = 8'b11000110; //  386 : 198 - 0xc6
      12'h183: dout  = 8'b11000110; //  387 : 198 - 0xc6
      12'h184: dout  = 8'b11000110; //  388 : 198 - 0xc6
      12'h185: dout  = 8'b11000110; //  389 : 198 - 0xc6
      12'h186: dout  = 8'b01111100; //  390 : 124 - 0x7c
      12'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      12'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      12'h18D: dout  = 8'b00000000; //  397 :   0 - 0x0
      12'h18E: dout  = 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout  = 8'b11111100; //  400 : 252 - 0xfc -- Background 0x19
      12'h191: dout  = 8'b11000110; //  401 : 198 - 0xc6
      12'h192: dout  = 8'b11000110; //  402 : 198 - 0xc6
      12'h193: dout  = 8'b11000110; //  403 : 198 - 0xc6
      12'h194: dout  = 8'b11111100; //  404 : 252 - 0xfc
      12'h195: dout  = 8'b11000000; //  405 : 192 - 0xc0
      12'h196: dout  = 8'b11000000; //  406 : 192 - 0xc0
      12'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout  = 8'b00000000; //  412 :   0 - 0x0
      12'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout  = 8'b01111100; //  416 : 124 - 0x7c -- Background 0x1a
      12'h1A1: dout  = 8'b11000110; //  417 : 198 - 0xc6
      12'h1A2: dout  = 8'b11000110; //  418 : 198 - 0xc6
      12'h1A3: dout  = 8'b11000110; //  419 : 198 - 0xc6
      12'h1A4: dout  = 8'b11011110; //  420 : 222 - 0xde
      12'h1A5: dout  = 8'b11001100; //  421 : 204 - 0xcc
      12'h1A6: dout  = 8'b01111010; //  422 : 122 - 0x7a
      12'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout  = 8'b00000000; //  424 :   0 - 0x0 -- plane 1
      12'h1A9: dout  = 8'b00000000; //  425 :   0 - 0x0
      12'h1AA: dout  = 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout  = 8'b11111100; //  432 : 252 - 0xfc -- Background 0x1b
      12'h1B1: dout  = 8'b11000110; //  433 : 198 - 0xc6
      12'h1B2: dout  = 8'b11000110; //  434 : 198 - 0xc6
      12'h1B3: dout  = 8'b11001110; //  435 : 206 - 0xce
      12'h1B4: dout  = 8'b11111000; //  436 : 248 - 0xf8
      12'h1B5: dout  = 8'b11011100; //  437 : 220 - 0xdc
      12'h1B6: dout  = 8'b11001110; //  438 : 206 - 0xce
      12'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout  = 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout  = 8'b00000000; //  441 :   0 - 0x0
      12'h1BA: dout  = 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout  = 8'b00000000; //  444 :   0 - 0x0
      12'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout  = 8'b01111000; //  448 : 120 - 0x78 -- Background 0x1c
      12'h1C1: dout  = 8'b11001100; //  449 : 204 - 0xcc
      12'h1C2: dout  = 8'b11000000; //  450 : 192 - 0xc0
      12'h1C3: dout  = 8'b01111100; //  451 : 124 - 0x7c
      12'h1C4: dout  = 8'b00000110; //  452 :   6 - 0x6
      12'h1C5: dout  = 8'b11000110; //  453 : 198 - 0xc6
      12'h1C6: dout  = 8'b01111100; //  454 : 124 - 0x7c
      12'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- plane 1
      12'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b01111110; //  464 : 126 - 0x7e -- Background 0x1d
      12'h1D1: dout  = 8'b00011000; //  465 :  24 - 0x18
      12'h1D2: dout  = 8'b00011000; //  466 :  24 - 0x18
      12'h1D3: dout  = 8'b00011000; //  467 :  24 - 0x18
      12'h1D4: dout  = 8'b00011000; //  468 :  24 - 0x18
      12'h1D5: dout  = 8'b00011000; //  469 :  24 - 0x18
      12'h1D6: dout  = 8'b00011000; //  470 :  24 - 0x18
      12'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- plane 1
      12'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout  = 8'b11000110; //  480 : 198 - 0xc6 -- Background 0x1e
      12'h1E1: dout  = 8'b11000110; //  481 : 198 - 0xc6
      12'h1E2: dout  = 8'b11000110; //  482 : 198 - 0xc6
      12'h1E3: dout  = 8'b11000110; //  483 : 198 - 0xc6
      12'h1E4: dout  = 8'b11000110; //  484 : 198 - 0xc6
      12'h1E5: dout  = 8'b11000110; //  485 : 198 - 0xc6
      12'h1E6: dout  = 8'b01111100; //  486 : 124 - 0x7c
      12'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- plane 1
      12'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout  = 8'b11000110; //  496 : 198 - 0xc6 -- Background 0x1f
      12'h1F1: dout  = 8'b11000110; //  497 : 198 - 0xc6
      12'h1F2: dout  = 8'b11000110; //  498 : 198 - 0xc6
      12'h1F3: dout  = 8'b11101110; //  499 : 238 - 0xee
      12'h1F4: dout  = 8'b01111100; //  500 : 124 - 0x7c
      12'h1F5: dout  = 8'b00111000; //  501 :  56 - 0x38
      12'h1F6: dout  = 8'b00010000; //  502 :  16 - 0x10
      12'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- plane 1
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout  = 8'b11000110; //  512 : 198 - 0xc6 -- Background 0x20
      12'h201: dout  = 8'b11000110; //  513 : 198 - 0xc6
      12'h202: dout  = 8'b11010110; //  514 : 214 - 0xd6
      12'h203: dout  = 8'b11111110; //  515 : 254 - 0xfe
      12'h204: dout  = 8'b11111110; //  516 : 254 - 0xfe
      12'h205: dout  = 8'b11101110; //  517 : 238 - 0xee
      12'h206: dout  = 8'b11000110; //  518 : 198 - 0xc6
      12'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout  = 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout  = 8'b11000110; //  528 : 198 - 0xc6 -- Background 0x21
      12'h211: dout  = 8'b11101110; //  529 : 238 - 0xee
      12'h212: dout  = 8'b01111100; //  530 : 124 - 0x7c
      12'h213: dout  = 8'b00111000; //  531 :  56 - 0x38
      12'h214: dout  = 8'b01111100; //  532 : 124 - 0x7c
      12'h215: dout  = 8'b11101110; //  533 : 238 - 0xee
      12'h216: dout  = 8'b11000110; //  534 : 198 - 0xc6
      12'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout  = 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout  = 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout  = 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout  = 8'b01100110; //  544 : 102 - 0x66 -- Background 0x22
      12'h221: dout  = 8'b01100110; //  545 : 102 - 0x66
      12'h222: dout  = 8'b01100110; //  546 : 102 - 0x66
      12'h223: dout  = 8'b00111100; //  547 :  60 - 0x3c
      12'h224: dout  = 8'b00011000; //  548 :  24 - 0x18
      12'h225: dout  = 8'b00011000; //  549 :  24 - 0x18
      12'h226: dout  = 8'b00011000; //  550 :  24 - 0x18
      12'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- plane 1
      12'h229: dout  = 8'b00000000; //  553 :   0 - 0x0
      12'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      12'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      12'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      12'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout  = 8'b11111110; //  560 : 254 - 0xfe -- Background 0x23
      12'h231: dout  = 8'b00001110; //  561 :  14 - 0xe
      12'h232: dout  = 8'b00011100; //  562 :  28 - 0x1c
      12'h233: dout  = 8'b00111000; //  563 :  56 - 0x38
      12'h234: dout  = 8'b01110000; //  564 : 112 - 0x70
      12'h235: dout  = 8'b11100000; //  565 : 224 - 0xe0
      12'h236: dout  = 8'b11111110; //  566 : 254 - 0xfe
      12'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout  = 8'b00000000; //  568 :   0 - 0x0 -- plane 1
      12'h239: dout  = 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout  = 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Background 0x24
      12'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout  = 8'b00000000; //  579 :   0 - 0x0
      12'h244: dout  = 8'b00000000; //  580 :   0 - 0x0
      12'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      12'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      12'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout  = 8'b00000000; //  584 :   0 - 0x0 -- plane 1
      12'h249: dout  = 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout  = 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b11111111; //  592 : 255 - 0xff -- Background 0x25
      12'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      12'h252: dout  = 8'b11111111; //  594 : 255 - 0xff
      12'h253: dout  = 8'b11111111; //  595 : 255 - 0xff
      12'h254: dout  = 8'b11111111; //  596 : 255 - 0xff
      12'h255: dout  = 8'b11111111; //  597 : 255 - 0xff
      12'h256: dout  = 8'b11111111; //  598 : 255 - 0xff
      12'h257: dout  = 8'b11111111; //  599 : 255 - 0xff
      12'h258: dout  = 8'b00000000; //  600 :   0 - 0x0 -- plane 1
      12'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout  = 8'b00000000; //  605 :   0 - 0x0
      12'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Background 0x26
      12'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      12'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      12'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      12'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      12'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      12'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout  = 8'b11111111; //  616 : 255 - 0xff -- plane 1
      12'h269: dout  = 8'b11111111; //  617 : 255 - 0xff
      12'h26A: dout  = 8'b11111111; //  618 : 255 - 0xff
      12'h26B: dout  = 8'b11111111; //  619 : 255 - 0xff
      12'h26C: dout  = 8'b11111111; //  620 : 255 - 0xff
      12'h26D: dout  = 8'b11111111; //  621 : 255 - 0xff
      12'h26E: dout  = 8'b11111111; //  622 : 255 - 0xff
      12'h26F: dout  = 8'b11111111; //  623 : 255 - 0xff
      12'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Background 0x27
      12'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      12'h272: dout  = 8'b11111111; //  626 : 255 - 0xff
      12'h273: dout  = 8'b11111111; //  627 : 255 - 0xff
      12'h274: dout  = 8'b11111111; //  628 : 255 - 0xff
      12'h275: dout  = 8'b11111111; //  629 : 255 - 0xff
      12'h276: dout  = 8'b11111111; //  630 : 255 - 0xff
      12'h277: dout  = 8'b11111111; //  631 : 255 - 0xff
      12'h278: dout  = 8'b11111111; //  632 : 255 - 0xff -- plane 1
      12'h279: dout  = 8'b11111111; //  633 : 255 - 0xff
      12'h27A: dout  = 8'b11111111; //  634 : 255 - 0xff
      12'h27B: dout  = 8'b11111111; //  635 : 255 - 0xff
      12'h27C: dout  = 8'b11111111; //  636 : 255 - 0xff
      12'h27D: dout  = 8'b11111111; //  637 : 255 - 0xff
      12'h27E: dout  = 8'b11111111; //  638 : 255 - 0xff
      12'h27F: dout  = 8'b11111111; //  639 : 255 - 0xff
      12'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Background 0x28
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout  = 8'b01111110; //  643 : 126 - 0x7e
      12'h284: dout  = 8'b01111110; //  644 : 126 - 0x7e
      12'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Background 0x29
      12'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout  = 8'b01000100; //  658 :  68 - 0x44
      12'h293: dout  = 8'b00101000; //  659 :  40 - 0x28
      12'h294: dout  = 8'b00010000; //  660 :  16 - 0x10
      12'h295: dout  = 8'b00101000; //  661 :  40 - 0x28
      12'h296: dout  = 8'b01000100; //  662 :  68 - 0x44
      12'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- plane 1
      12'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout  = 8'b11111111; //  672 : 255 - 0xff -- Background 0x2a
      12'h2A1: dout  = 8'b11111111; //  673 : 255 - 0xff
      12'h2A2: dout  = 8'b11111111; //  674 : 255 - 0xff
      12'h2A3: dout  = 8'b11111111; //  675 : 255 - 0xff
      12'h2A4: dout  = 8'b11111111; //  676 : 255 - 0xff
      12'h2A5: dout  = 8'b11111111; //  677 : 255 - 0xff
      12'h2A6: dout  = 8'b11111111; //  678 : 255 - 0xff
      12'h2A7: dout  = 8'b11111111; //  679 : 255 - 0xff
      12'h2A8: dout  = 8'b01111111; //  680 : 127 - 0x7f -- plane 1
      12'h2A9: dout  = 8'b01111111; //  681 : 127 - 0x7f
      12'h2AA: dout  = 8'b01111111; //  682 : 127 - 0x7f
      12'h2AB: dout  = 8'b01111111; //  683 : 127 - 0x7f
      12'h2AC: dout  = 8'b01111111; //  684 : 127 - 0x7f
      12'h2AD: dout  = 8'b01111111; //  685 : 127 - 0x7f
      12'h2AE: dout  = 8'b01111111; //  686 : 127 - 0x7f
      12'h2AF: dout  = 8'b01111111; //  687 : 127 - 0x7f
      12'h2B0: dout  = 8'b00011000; //  688 :  24 - 0x18 -- Background 0x2b
      12'h2B1: dout  = 8'b00111100; //  689 :  60 - 0x3c
      12'h2B2: dout  = 8'b00111100; //  690 :  60 - 0x3c
      12'h2B3: dout  = 8'b00111100; //  691 :  60 - 0x3c
      12'h2B4: dout  = 8'b00011000; //  692 :  24 - 0x18
      12'h2B5: dout  = 8'b00011000; //  693 :  24 - 0x18
      12'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout  = 8'b00011000; //  695 :  24 - 0x18
      12'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- plane 1
      12'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b11111111; //  704 : 255 - 0xff -- Background 0x2c
      12'h2C1: dout  = 8'b01111111; //  705 : 127 - 0x7f
      12'h2C2: dout  = 8'b01111111; //  706 : 127 - 0x7f
      12'h2C3: dout  = 8'b01111111; //  707 : 127 - 0x7f
      12'h2C4: dout  = 8'b01111111; //  708 : 127 - 0x7f
      12'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      12'h2C6: dout  = 8'b11100011; //  710 : 227 - 0xe3
      12'h2C7: dout  = 8'b11000001; //  711 : 193 - 0xc1
      12'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- plane 1
      12'h2C9: dout  = 8'b10000000; //  713 : 128 - 0x80
      12'h2CA: dout  = 8'b10000000; //  714 : 128 - 0x80
      12'h2CB: dout  = 8'b10000000; //  715 : 128 - 0x80
      12'h2CC: dout  = 8'b10000000; //  716 : 128 - 0x80
      12'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout  = 8'b00011100; //  718 :  28 - 0x1c
      12'h2CF: dout  = 8'b00111110; //  719 :  62 - 0x3e
      12'h2D0: dout  = 8'b10000000; //  720 : 128 - 0x80 -- Background 0x2d
      12'h2D1: dout  = 8'b10000000; //  721 : 128 - 0x80
      12'h2D2: dout  = 8'b10000000; //  722 : 128 - 0x80
      12'h2D3: dout  = 8'b11000001; //  723 : 193 - 0xc1
      12'h2D4: dout  = 8'b11100011; //  724 : 227 - 0xe3
      12'h2D5: dout  = 8'b11111111; //  725 : 255 - 0xff
      12'h2D6: dout  = 8'b11111111; //  726 : 255 - 0xff
      12'h2D7: dout  = 8'b11111111; //  727 : 255 - 0xff
      12'h2D8: dout  = 8'b01111111; //  728 : 127 - 0x7f -- plane 1
      12'h2D9: dout  = 8'b01111111; //  729 : 127 - 0x7f
      12'h2DA: dout  = 8'b01111111; //  730 : 127 - 0x7f
      12'h2DB: dout  = 8'b00111110; //  731 :  62 - 0x3e
      12'h2DC: dout  = 8'b00011100; //  732 :  28 - 0x1c
      12'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      12'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      12'h2DF: dout  = 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout  = 8'b00111000; //  736 :  56 - 0x38 -- Background 0x2e
      12'h2E1: dout  = 8'b01111100; //  737 : 124 - 0x7c
      12'h2E2: dout  = 8'b01111100; //  738 : 124 - 0x7c
      12'h2E3: dout  = 8'b01111100; //  739 : 124 - 0x7c
      12'h2E4: dout  = 8'b01111100; //  740 : 124 - 0x7c
      12'h2E5: dout  = 8'b01111100; //  741 : 124 - 0x7c
      12'h2E6: dout  = 8'b00111000; //  742 :  56 - 0x38
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b00001000; //  744 :   8 - 0x8 -- plane 1
      12'h2E9: dout  = 8'b00000100; //  745 :   4 - 0x4
      12'h2EA: dout  = 8'b00000100; //  746 :   4 - 0x4
      12'h2EB: dout  = 8'b00000100; //  747 :   4 - 0x4
      12'h2EC: dout  = 8'b00000100; //  748 :   4 - 0x4
      12'h2ED: dout  = 8'b00000100; //  749 :   4 - 0x4
      12'h2EE: dout  = 8'b00001000; //  750 :   8 - 0x8
      12'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout  = 8'b00000011; //  752 :   3 - 0x3 -- Background 0x2f
      12'h2F1: dout  = 8'b00000110; //  753 :   6 - 0x6
      12'h2F2: dout  = 8'b00001100; //  754 :  12 - 0xc
      12'h2F3: dout  = 8'b00001100; //  755 :  12 - 0xc
      12'h2F4: dout  = 8'b00001000; //  756 :   8 - 0x8
      12'h2F5: dout  = 8'b00001000; //  757 :   8 - 0x8
      12'h2F6: dout  = 8'b00000100; //  758 :   4 - 0x4
      12'h2F7: dout  = 8'b00000011; //  759 :   3 - 0x3
      12'h2F8: dout  = 8'b00000011; //  760 :   3 - 0x3 -- plane 1
      12'h2F9: dout  = 8'b00000101; //  761 :   5 - 0x5
      12'h2FA: dout  = 8'b00001011; //  762 :  11 - 0xb
      12'h2FB: dout  = 8'b00001011; //  763 :  11 - 0xb
      12'h2FC: dout  = 8'b00001111; //  764 :  15 - 0xf
      12'h2FD: dout  = 8'b00001111; //  765 :  15 - 0xf
      12'h2FE: dout  = 8'b00000111; //  766 :   7 - 0x7
      12'h2FF: dout  = 8'b00000011; //  767 :   3 - 0x3
      12'h300: dout  = 8'b00000001; //  768 :   1 - 0x1 -- Background 0x30
      12'h301: dout  = 8'b00000010; //  769 :   2 - 0x2
      12'h302: dout  = 8'b00000100; //  770 :   4 - 0x4
      12'h303: dout  = 8'b00001000; //  771 :   8 - 0x8
      12'h304: dout  = 8'b00010000; //  772 :  16 - 0x10
      12'h305: dout  = 8'b00100000; //  773 :  32 - 0x20
      12'h306: dout  = 8'b01000000; //  774 :  64 - 0x40
      12'h307: dout  = 8'b10000000; //  775 : 128 - 0x80
      12'h308: dout  = 8'b00000001; //  776 :   1 - 0x1 -- plane 1
      12'h309: dout  = 8'b00000011; //  777 :   3 - 0x3
      12'h30A: dout  = 8'b00000111; //  778 :   7 - 0x7
      12'h30B: dout  = 8'b00001111; //  779 :  15 - 0xf
      12'h30C: dout  = 8'b00011111; //  780 :  31 - 0x1f
      12'h30D: dout  = 8'b00111111; //  781 :  63 - 0x3f
      12'h30E: dout  = 8'b01111111; //  782 : 127 - 0x7f
      12'h30F: dout  = 8'b11111111; //  783 : 255 - 0xff
      12'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Background 0x31
      12'h311: dout  = 8'b00000000; //  785 :   0 - 0x0
      12'h312: dout  = 8'b00000000; //  786 :   0 - 0x0
      12'h313: dout  = 8'b00000000; //  787 :   0 - 0x0
      12'h314: dout  = 8'b00000000; //  788 :   0 - 0x0
      12'h315: dout  = 8'b00000111; //  789 :   7 - 0x7
      12'h316: dout  = 8'b00111000; //  790 :  56 - 0x38
      12'h317: dout  = 8'b11000000; //  791 : 192 - 0xc0
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout  = 8'b00000111; //  797 :   7 - 0x7
      12'h31E: dout  = 8'b00111111; //  798 :  63 - 0x3f
      12'h31F: dout  = 8'b11111111; //  799 : 255 - 0xff
      12'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Background 0x32
      12'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout  = 8'b00000000; //  802 :   0 - 0x0
      12'h323: dout  = 8'b00000000; //  803 :   0 - 0x0
      12'h324: dout  = 8'b00000000; //  804 :   0 - 0x0
      12'h325: dout  = 8'b11100000; //  805 : 224 - 0xe0
      12'h326: dout  = 8'b00011100; //  806 :  28 - 0x1c
      12'h327: dout  = 8'b00000011; //  807 :   3 - 0x3
      12'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout  = 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout  = 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout  = 8'b11100000; //  813 : 224 - 0xe0
      12'h32E: dout  = 8'b11111100; //  814 : 252 - 0xfc
      12'h32F: dout  = 8'b11111111; //  815 : 255 - 0xff
      12'h330: dout  = 8'b10000000; //  816 : 128 - 0x80 -- Background 0x33
      12'h331: dout  = 8'b01000000; //  817 :  64 - 0x40
      12'h332: dout  = 8'b00100000; //  818 :  32 - 0x20
      12'h333: dout  = 8'b00010000; //  819 :  16 - 0x10
      12'h334: dout  = 8'b00001000; //  820 :   8 - 0x8
      12'h335: dout  = 8'b00000100; //  821 :   4 - 0x4
      12'h336: dout  = 8'b00000010; //  822 :   2 - 0x2
      12'h337: dout  = 8'b00000001; //  823 :   1 - 0x1
      12'h338: dout  = 8'b10000000; //  824 : 128 - 0x80 -- plane 1
      12'h339: dout  = 8'b11000000; //  825 : 192 - 0xc0
      12'h33A: dout  = 8'b11100000; //  826 : 224 - 0xe0
      12'h33B: dout  = 8'b11110000; //  827 : 240 - 0xf0
      12'h33C: dout  = 8'b11111000; //  828 : 248 - 0xf8
      12'h33D: dout  = 8'b11111100; //  829 : 252 - 0xfc
      12'h33E: dout  = 8'b11111110; //  830 : 254 - 0xfe
      12'h33F: dout  = 8'b11111111; //  831 : 255 - 0xff
      12'h340: dout  = 8'b00000100; //  832 :   4 - 0x4 -- Background 0x34
      12'h341: dout  = 8'b00001110; //  833 :  14 - 0xe
      12'h342: dout  = 8'b00001110; //  834 :  14 - 0xe
      12'h343: dout  = 8'b00001110; //  835 :  14 - 0xe
      12'h344: dout  = 8'b01101110; //  836 : 110 - 0x6e
      12'h345: dout  = 8'b01100100; //  837 : 100 - 0x64
      12'h346: dout  = 8'b01100000; //  838 :  96 - 0x60
      12'h347: dout  = 8'b01100000; //  839 :  96 - 0x60
      12'h348: dout  = 8'b11111111; //  840 : 255 - 0xff -- plane 1
      12'h349: dout  = 8'b11111111; //  841 : 255 - 0xff
      12'h34A: dout  = 8'b11111111; //  842 : 255 - 0xff
      12'h34B: dout  = 8'b11111111; //  843 : 255 - 0xff
      12'h34C: dout  = 8'b11111111; //  844 : 255 - 0xff
      12'h34D: dout  = 8'b11111111; //  845 : 255 - 0xff
      12'h34E: dout  = 8'b11111111; //  846 : 255 - 0xff
      12'h34F: dout  = 8'b11111111; //  847 : 255 - 0xff
      12'h350: dout  = 8'b00000111; //  848 :   7 - 0x7 -- Background 0x35
      12'h351: dout  = 8'b00001111; //  849 :  15 - 0xf
      12'h352: dout  = 8'b00011111; //  850 :  31 - 0x1f
      12'h353: dout  = 8'b00011111; //  851 :  31 - 0x1f
      12'h354: dout  = 8'b01111111; //  852 : 127 - 0x7f
      12'h355: dout  = 8'b11111111; //  853 : 255 - 0xff
      12'h356: dout  = 8'b11111111; //  854 : 255 - 0xff
      12'h357: dout  = 8'b01111111; //  855 : 127 - 0x7f
      12'h358: dout  = 8'b00000111; //  856 :   7 - 0x7 -- plane 1
      12'h359: dout  = 8'b00001000; //  857 :   8 - 0x8
      12'h35A: dout  = 8'b00010000; //  858 :  16 - 0x10
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b01100000; //  860 :  96 - 0x60
      12'h35D: dout  = 8'b10000000; //  861 : 128 - 0x80
      12'h35E: dout  = 8'b10000000; //  862 : 128 - 0x80
      12'h35F: dout  = 8'b01000000; //  863 :  64 - 0x40
      12'h360: dout  = 8'b00000011; //  864 :   3 - 0x3 -- Background 0x36
      12'h361: dout  = 8'b00000111; //  865 :   7 - 0x7
      12'h362: dout  = 8'b00011111; //  866 :  31 - 0x1f
      12'h363: dout  = 8'b00111111; //  867 :  63 - 0x3f
      12'h364: dout  = 8'b00111111; //  868 :  63 - 0x3f
      12'h365: dout  = 8'b00111111; //  869 :  63 - 0x3f
      12'h366: dout  = 8'b01111001; //  870 : 121 - 0x79
      12'h367: dout  = 8'b11110111; //  871 : 247 - 0xf7
      12'h368: dout  = 8'b00000011; //  872 :   3 - 0x3 -- plane 1
      12'h369: dout  = 8'b00000100; //  873 :   4 - 0x4
      12'h36A: dout  = 8'b00011000; //  874 :  24 - 0x18
      12'h36B: dout  = 8'b00100000; //  875 :  32 - 0x20
      12'h36C: dout  = 8'b00100000; //  876 :  32 - 0x20
      12'h36D: dout  = 8'b00100000; //  877 :  32 - 0x20
      12'h36E: dout  = 8'b01000110; //  878 :  70 - 0x46
      12'h36F: dout  = 8'b10001000; //  879 : 136 - 0x88
      12'h370: dout  = 8'b11000000; //  880 : 192 - 0xc0 -- Background 0x37
      12'h371: dout  = 8'b11100000; //  881 : 224 - 0xe0
      12'h372: dout  = 8'b11110000; //  882 : 240 - 0xf0
      12'h373: dout  = 8'b11110100; //  883 : 244 - 0xf4
      12'h374: dout  = 8'b11111110; //  884 : 254 - 0xfe
      12'h375: dout  = 8'b10111111; //  885 : 191 - 0xbf
      12'h376: dout  = 8'b11011111; //  886 : 223 - 0xdf
      12'h377: dout  = 8'b11111111; //  887 : 255 - 0xff
      12'h378: dout  = 8'b11000000; //  888 : 192 - 0xc0 -- plane 1
      12'h379: dout  = 8'b00100000; //  889 :  32 - 0x20
      12'h37A: dout  = 8'b00010000; //  890 :  16 - 0x10
      12'h37B: dout  = 8'b00010100; //  891 :  20 - 0x14
      12'h37C: dout  = 8'b00001010; //  892 :  10 - 0xa
      12'h37D: dout  = 8'b01000001; //  893 :  65 - 0x41
      12'h37E: dout  = 8'b00100001; //  894 :  33 - 0x21
      12'h37F: dout  = 8'b00000001; //  895 :   1 - 0x1
      12'h380: dout  = 8'b10010000; //  896 : 144 - 0x90 -- Background 0x38
      12'h381: dout  = 8'b10111000; //  897 : 184 - 0xb8
      12'h382: dout  = 8'b11111000; //  898 : 248 - 0xf8
      12'h383: dout  = 8'b11111010; //  899 : 250 - 0xfa
      12'h384: dout  = 8'b11111111; //  900 : 255 - 0xff
      12'h385: dout  = 8'b11111111; //  901 : 255 - 0xff
      12'h386: dout  = 8'b11111111; //  902 : 255 - 0xff
      12'h387: dout  = 8'b11111110; //  903 : 254 - 0xfe
      12'h388: dout  = 8'b10010000; //  904 : 144 - 0x90 -- plane 1
      12'h389: dout  = 8'b10101000; //  905 : 168 - 0xa8
      12'h38A: dout  = 8'b01001000; //  906 :  72 - 0x48
      12'h38B: dout  = 8'b00001010; //  907 :  10 - 0xa
      12'h38C: dout  = 8'b00000101; //  908 :   5 - 0x5
      12'h38D: dout  = 8'b00000001; //  909 :   1 - 0x1
      12'h38E: dout  = 8'b00000001; //  910 :   1 - 0x1
      12'h38F: dout  = 8'b00000010; //  911 :   2 - 0x2
      12'h390: dout  = 8'b00111011; //  912 :  59 - 0x3b -- Background 0x39
      12'h391: dout  = 8'b00011101; //  913 :  29 - 0x1d
      12'h392: dout  = 8'b00001110; //  914 :  14 - 0xe
      12'h393: dout  = 8'b00001111; //  915 :  15 - 0xf
      12'h394: dout  = 8'b00000111; //  916 :   7 - 0x7
      12'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b00100100; //  920 :  36 - 0x24 -- plane 1
      12'h399: dout  = 8'b00010010; //  921 :  18 - 0x12
      12'h39A: dout  = 8'b00001001; //  922 :   9 - 0x9
      12'h39B: dout  = 8'b00001000; //  923 :   8 - 0x8
      12'h39C: dout  = 8'b00000111; //  924 :   7 - 0x7
      12'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b11111111; //  928 : 255 - 0xff -- Background 0x3a
      12'h3A1: dout  = 8'b10111111; //  929 : 191 - 0xbf
      12'h3A2: dout  = 8'b00011100; //  930 :  28 - 0x1c
      12'h3A3: dout  = 8'b11000000; //  931 : 192 - 0xc0
      12'h3A4: dout  = 8'b11110011; //  932 : 243 - 0xf3
      12'h3A5: dout  = 8'b11111111; //  933 : 255 - 0xff
      12'h3A6: dout  = 8'b01111110; //  934 : 126 - 0x7e
      12'h3A7: dout  = 8'b00011100; //  935 :  28 - 0x1c
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout  = 8'b01000000; //  937 :  64 - 0x40
      12'h3AA: dout  = 8'b11100011; //  938 : 227 - 0xe3
      12'h3AB: dout  = 8'b00111111; //  939 :  63 - 0x3f
      12'h3AC: dout  = 8'b00001100; //  940 :  12 - 0xc
      12'h3AD: dout  = 8'b10000001; //  941 : 129 - 0x81
      12'h3AE: dout  = 8'b01100010; //  942 :  98 - 0x62
      12'h3AF: dout  = 8'b00011100; //  943 :  28 - 0x1c
      12'h3B0: dout  = 8'b10111111; //  944 : 191 - 0xbf -- Background 0x3b
      12'h3B1: dout  = 8'b01111111; //  945 : 127 - 0x7f
      12'h3B2: dout  = 8'b00111101; //  946 :  61 - 0x3d
      12'h3B3: dout  = 8'b10000011; //  947 : 131 - 0x83
      12'h3B4: dout  = 8'b11000111; //  948 : 199 - 0xc7
      12'h3B5: dout  = 8'b11111111; //  949 : 255 - 0xff
      12'h3B6: dout  = 8'b11111111; //  950 : 255 - 0xff
      12'h3B7: dout  = 8'b00111100; //  951 :  60 - 0x3c
      12'h3B8: dout  = 8'b01000000; //  952 :  64 - 0x40 -- plane 1
      12'h3B9: dout  = 8'b10000000; //  953 : 128 - 0x80
      12'h3BA: dout  = 8'b11000010; //  954 : 194 - 0xc2
      12'h3BB: dout  = 8'b01111100; //  955 : 124 - 0x7c
      12'h3BC: dout  = 8'b00111000; //  956 :  56 - 0x38
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b11000011; //  958 : 195 - 0xc3
      12'h3BF: dout  = 8'b00111100; //  959 :  60 - 0x3c
      12'h3C0: dout  = 8'b11111100; //  960 : 252 - 0xfc -- Background 0x3c
      12'h3C1: dout  = 8'b11111110; //  961 : 254 - 0xfe
      12'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout  = 8'b11111110; //  963 : 254 - 0xfe
      12'h3C4: dout  = 8'b11111110; //  964 : 254 - 0xfe
      12'h3C5: dout  = 8'b11111000; //  965 : 248 - 0xf8
      12'h3C6: dout  = 8'b01100000; //  966 :  96 - 0x60
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b00000100; //  968 :   4 - 0x4 -- plane 1
      12'h3C9: dout  = 8'b00000010; //  969 :   2 - 0x2
      12'h3CA: dout  = 8'b00000001; //  970 :   1 - 0x1
      12'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout  = 8'b00000110; //  972 :   6 - 0x6
      12'h3CD: dout  = 8'b10011000; //  973 : 152 - 0x98
      12'h3CE: dout  = 8'b01100000; //  974 :  96 - 0x60
      12'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout  = 8'b11000000; //  976 : 192 - 0xc0 -- Background 0x3d
      12'h3D1: dout  = 8'b00100000; //  977 :  32 - 0x20
      12'h3D2: dout  = 8'b00010000; //  978 :  16 - 0x10
      12'h3D3: dout  = 8'b00010000; //  979 :  16 - 0x10
      12'h3D4: dout  = 8'b00010000; //  980 :  16 - 0x10
      12'h3D5: dout  = 8'b00010000; //  981 :  16 - 0x10
      12'h3D6: dout  = 8'b00100000; //  982 :  32 - 0x20
      12'h3D7: dout  = 8'b11000000; //  983 : 192 - 0xc0
      12'h3D8: dout  = 8'b11000000; //  984 : 192 - 0xc0 -- plane 1
      12'h3D9: dout  = 8'b11100000; //  985 : 224 - 0xe0
      12'h3DA: dout  = 8'b11110000; //  986 : 240 - 0xf0
      12'h3DB: dout  = 8'b11110000; //  987 : 240 - 0xf0
      12'h3DC: dout  = 8'b11110000; //  988 : 240 - 0xf0
      12'h3DD: dout  = 8'b11110000; //  989 : 240 - 0xf0
      12'h3DE: dout  = 8'b11100000; //  990 : 224 - 0xe0
      12'h3DF: dout  = 8'b11000000; //  991 : 192 - 0xc0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Background 0x3e
      12'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00111111; //  996 :  63 - 0x3f
      12'h3E5: dout  = 8'b01111111; //  997 : 127 - 0x7f
      12'h3E6: dout  = 8'b11100000; //  998 : 224 - 0xe0
      12'h3E7: dout  = 8'b11000000; //  999 : 192 - 0xc0
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00011100; // 1006 :  28 - 0x1c
      12'h3EF: dout  = 8'b00111110; // 1007 :  62 - 0x3e
      12'h3F0: dout  = 8'b10001000; // 1008 : 136 - 0x88 -- Background 0x3f
      12'h3F1: dout  = 8'b10011100; // 1009 : 156 - 0x9c
      12'h3F2: dout  = 8'b10001000; // 1010 : 136 - 0x88
      12'h3F3: dout  = 8'b10000000; // 1011 : 128 - 0x80
      12'h3F4: dout  = 8'b10000000; // 1012 : 128 - 0x80
      12'h3F5: dout  = 8'b10000000; // 1013 : 128 - 0x80
      12'h3F6: dout  = 8'b10000000; // 1014 : 128 - 0x80
      12'h3F7: dout  = 8'b10000000; // 1015 : 128 - 0x80
      12'h3F8: dout  = 8'b01111111; // 1016 : 127 - 0x7f -- plane 1
      12'h3F9: dout  = 8'b01111111; // 1017 : 127 - 0x7f
      12'h3FA: dout  = 8'b01111111; // 1018 : 127 - 0x7f
      12'h3FB: dout  = 8'b00111110; // 1019 :  62 - 0x3e
      12'h3FC: dout  = 8'b00011100; // 1020 :  28 - 0x1c
      12'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout  = 8'b11111110; // 1024 : 254 - 0xfe -- Background 0x40
      12'h401: dout  = 8'b11111110; // 1025 : 254 - 0xfe
      12'h402: dout  = 8'b11111110; // 1026 : 254 - 0xfe
      12'h403: dout  = 8'b11111110; // 1027 : 254 - 0xfe
      12'h404: dout  = 8'b11111110; // 1028 : 254 - 0xfe
      12'h405: dout  = 8'b11111110; // 1029 : 254 - 0xfe
      12'h406: dout  = 8'b11111110; // 1030 : 254 - 0xfe
      12'h407: dout  = 8'b11111110; // 1031 : 254 - 0xfe
      12'h408: dout  = 8'b11111111; // 1032 : 255 - 0xff -- plane 1
      12'h409: dout  = 8'b11111111; // 1033 : 255 - 0xff
      12'h40A: dout  = 8'b11111111; // 1034 : 255 - 0xff
      12'h40B: dout  = 8'b11111111; // 1035 : 255 - 0xff
      12'h40C: dout  = 8'b11111111; // 1036 : 255 - 0xff
      12'h40D: dout  = 8'b11111111; // 1037 : 255 - 0xff
      12'h40E: dout  = 8'b11111111; // 1038 : 255 - 0xff
      12'h40F: dout  = 8'b11111111; // 1039 : 255 - 0xff
      12'h410: dout  = 8'b00001000; // 1040 :   8 - 0x8 -- Background 0x41
      12'h411: dout  = 8'b00010100; // 1041 :  20 - 0x14
      12'h412: dout  = 8'b00100100; // 1042 :  36 - 0x24
      12'h413: dout  = 8'b11000100; // 1043 : 196 - 0xc4
      12'h414: dout  = 8'b00000011; // 1044 :   3 - 0x3
      12'h415: dout  = 8'b01000000; // 1045 :  64 - 0x40
      12'h416: dout  = 8'b10100001; // 1046 : 161 - 0xa1
      12'h417: dout  = 8'b00100110; // 1047 :  38 - 0x26
      12'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout  = 8'b00001000; // 1049 :   8 - 0x8
      12'h41A: dout  = 8'b00011000; // 1050 :  24 - 0x18
      12'h41B: dout  = 8'b00111000; // 1051 :  56 - 0x38
      12'h41C: dout  = 8'b11111100; // 1052 : 252 - 0xfc
      12'h41D: dout  = 8'b10111111; // 1053 : 191 - 0xbf
      12'h41E: dout  = 8'b01011110; // 1054 :  94 - 0x5e
      12'h41F: dout  = 8'b11011001; // 1055 : 217 - 0xd9
      12'h420: dout  = 8'b11111111; // 1056 : 255 - 0xff -- Background 0x42
      12'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      12'h422: dout  = 8'b11111111; // 1058 : 255 - 0xff
      12'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      12'h424: dout  = 8'b01111111; // 1060 : 127 - 0x7f
      12'h425: dout  = 8'b01111111; // 1061 : 127 - 0x7f
      12'h426: dout  = 8'b01111111; // 1062 : 127 - 0x7f
      12'h427: dout  = 8'b01111111; // 1063 : 127 - 0x7f
      12'h428: dout  = 8'b10000001; // 1064 : 129 - 0x81 -- plane 1
      12'h429: dout  = 8'b10000001; // 1065 : 129 - 0x81
      12'h42A: dout  = 8'b10000001; // 1066 : 129 - 0x81
      12'h42B: dout  = 8'b10000001; // 1067 : 129 - 0x81
      12'h42C: dout  = 8'b10000001; // 1068 : 129 - 0x81
      12'h42D: dout  = 8'b10000001; // 1069 : 129 - 0x81
      12'h42E: dout  = 8'b10000001; // 1070 : 129 - 0x81
      12'h42F: dout  = 8'b10000001; // 1071 : 129 - 0x81
      12'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Background 0x43
      12'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      12'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      12'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      12'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      12'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      12'h436: dout  = 8'b11111111; // 1078 : 255 - 0xff
      12'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      12'h438: dout  = 8'b00000001; // 1080 :   1 - 0x1 -- plane 1
      12'h439: dout  = 8'b00000001; // 1081 :   1 - 0x1
      12'h43A: dout  = 8'b00000001; // 1082 :   1 - 0x1
      12'h43B: dout  = 8'b00000001; // 1083 :   1 - 0x1
      12'h43C: dout  = 8'b00000001; // 1084 :   1 - 0x1
      12'h43D: dout  = 8'b00000001; // 1085 :   1 - 0x1
      12'h43E: dout  = 8'b00000001; // 1086 :   1 - 0x1
      12'h43F: dout  = 8'b00000001; // 1087 :   1 - 0x1
      12'h440: dout  = 8'b01111111; // 1088 : 127 - 0x7f -- Background 0x44
      12'h441: dout  = 8'b10000000; // 1089 : 128 - 0x80
      12'h442: dout  = 8'b10000000; // 1090 : 128 - 0x80
      12'h443: dout  = 8'b10011000; // 1091 : 152 - 0x98
      12'h444: dout  = 8'b10011100; // 1092 : 156 - 0x9c
      12'h445: dout  = 8'b10001100; // 1093 : 140 - 0x8c
      12'h446: dout  = 8'b10000000; // 1094 : 128 - 0x80
      12'h447: dout  = 8'b10000000; // 1095 : 128 - 0x80
      12'h448: dout  = 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout  = 8'b01111111; // 1097 : 127 - 0x7f
      12'h44A: dout  = 8'b01111111; // 1098 : 127 - 0x7f
      12'h44B: dout  = 8'b01100111; // 1099 : 103 - 0x67
      12'h44C: dout  = 8'b01100111; // 1100 : 103 - 0x67
      12'h44D: dout  = 8'b01111111; // 1101 : 127 - 0x7f
      12'h44E: dout  = 8'b01111111; // 1102 : 127 - 0x7f
      12'h44F: dout  = 8'b01111111; // 1103 : 127 - 0x7f
      12'h450: dout  = 8'b11111111; // 1104 : 255 - 0xff -- Background 0x45
      12'h451: dout  = 8'b00000001; // 1105 :   1 - 0x1
      12'h452: dout  = 8'b00000001; // 1106 :   1 - 0x1
      12'h453: dout  = 8'b11111111; // 1107 : 255 - 0xff
      12'h454: dout  = 8'b00010000; // 1108 :  16 - 0x10
      12'h455: dout  = 8'b00010000; // 1109 :  16 - 0x10
      12'h456: dout  = 8'b00010000; // 1110 :  16 - 0x10
      12'h457: dout  = 8'b11111111; // 1111 : 255 - 0xff
      12'h458: dout  = 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout  = 8'b11111111; // 1113 : 255 - 0xff
      12'h45A: dout  = 8'b11111111; // 1114 : 255 - 0xff
      12'h45B: dout  = 8'b11111111; // 1115 : 255 - 0xff
      12'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      12'h45D: dout  = 8'b11111111; // 1117 : 255 - 0xff
      12'h45E: dout  = 8'b11111111; // 1118 : 255 - 0xff
      12'h45F: dout  = 8'b11111111; // 1119 : 255 - 0xff
      12'h460: dout  = 8'b10000000; // 1120 : 128 - 0x80 -- Background 0x46
      12'h461: dout  = 8'b10000000; // 1121 : 128 - 0x80
      12'h462: dout  = 8'b10000000; // 1122 : 128 - 0x80
      12'h463: dout  = 8'b10000000; // 1123 : 128 - 0x80
      12'h464: dout  = 8'b10000000; // 1124 : 128 - 0x80
      12'h465: dout  = 8'b10000000; // 1125 : 128 - 0x80
      12'h466: dout  = 8'b10000000; // 1126 : 128 - 0x80
      12'h467: dout  = 8'b10000000; // 1127 : 128 - 0x80
      12'h468: dout  = 8'b01111111; // 1128 : 127 - 0x7f -- plane 1
      12'h469: dout  = 8'b01111111; // 1129 : 127 - 0x7f
      12'h46A: dout  = 8'b01111111; // 1130 : 127 - 0x7f
      12'h46B: dout  = 8'b01111111; // 1131 : 127 - 0x7f
      12'h46C: dout  = 8'b01111111; // 1132 : 127 - 0x7f
      12'h46D: dout  = 8'b01111111; // 1133 : 127 - 0x7f
      12'h46E: dout  = 8'b01111111; // 1134 : 127 - 0x7f
      12'h46F: dout  = 8'b01111111; // 1135 : 127 - 0x7f
      12'h470: dout  = 8'b00000001; // 1136 :   1 - 0x1 -- Background 0x47
      12'h471: dout  = 8'b00000001; // 1137 :   1 - 0x1
      12'h472: dout  = 8'b00000001; // 1138 :   1 - 0x1
      12'h473: dout  = 8'b11111111; // 1139 : 255 - 0xff
      12'h474: dout  = 8'b00010000; // 1140 :  16 - 0x10
      12'h475: dout  = 8'b00010000; // 1141 :  16 - 0x10
      12'h476: dout  = 8'b00010000; // 1142 :  16 - 0x10
      12'h477: dout  = 8'b11111111; // 1143 : 255 - 0xff
      12'h478: dout  = 8'b11111111; // 1144 : 255 - 0xff -- plane 1
      12'h479: dout  = 8'b11111111; // 1145 : 255 - 0xff
      12'h47A: dout  = 8'b11111111; // 1146 : 255 - 0xff
      12'h47B: dout  = 8'b11111111; // 1147 : 255 - 0xff
      12'h47C: dout  = 8'b11111111; // 1148 : 255 - 0xff
      12'h47D: dout  = 8'b11111111; // 1149 : 255 - 0xff
      12'h47E: dout  = 8'b11111111; // 1150 : 255 - 0xff
      12'h47F: dout  = 8'b11111111; // 1151 : 255 - 0xff
      12'h480: dout  = 8'b11111111; // 1152 : 255 - 0xff -- Background 0x48
      12'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout  = 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      12'h48A: dout  = 8'b11111111; // 1162 : 255 - 0xff
      12'h48B: dout  = 8'b11111111; // 1163 : 255 - 0xff
      12'h48C: dout  = 8'b11111111; // 1164 : 255 - 0xff
      12'h48D: dout  = 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout  = 8'b11111111; // 1166 : 255 - 0xff
      12'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      12'h490: dout  = 8'b11111110; // 1168 : 254 - 0xfe -- Background 0x49
      12'h491: dout  = 8'b00000001; // 1169 :   1 - 0x1
      12'h492: dout  = 8'b00000001; // 1170 :   1 - 0x1
      12'h493: dout  = 8'b00011001; // 1171 :  25 - 0x19
      12'h494: dout  = 8'b00011101; // 1172 :  29 - 0x1d
      12'h495: dout  = 8'b00001101; // 1173 :  13 - 0xd
      12'h496: dout  = 8'b00000001; // 1174 :   1 - 0x1
      12'h497: dout  = 8'b00000001; // 1175 :   1 - 0x1
      12'h498: dout  = 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout  = 8'b11111111; // 1177 : 255 - 0xff
      12'h49A: dout  = 8'b11111111; // 1178 : 255 - 0xff
      12'h49B: dout  = 8'b11100111; // 1179 : 231 - 0xe7
      12'h49C: dout  = 8'b11100111; // 1180 : 231 - 0xe7
      12'h49D: dout  = 8'b11111111; // 1181 : 255 - 0xff
      12'h49E: dout  = 8'b11111111; // 1182 : 255 - 0xff
      12'h49F: dout  = 8'b11111111; // 1183 : 255 - 0xff
      12'h4A0: dout  = 8'b00000001; // 1184 :   1 - 0x1 -- Background 0x4a
      12'h4A1: dout  = 8'b00000001; // 1185 :   1 - 0x1
      12'h4A2: dout  = 8'b00000001; // 1186 :   1 - 0x1
      12'h4A3: dout  = 8'b00000001; // 1187 :   1 - 0x1
      12'h4A4: dout  = 8'b00000001; // 1188 :   1 - 0x1
      12'h4A5: dout  = 8'b00000001; // 1189 :   1 - 0x1
      12'h4A6: dout  = 8'b00000001; // 1190 :   1 - 0x1
      12'h4A7: dout  = 8'b00000001; // 1191 :   1 - 0x1
      12'h4A8: dout  = 8'b11111111; // 1192 : 255 - 0xff -- plane 1
      12'h4A9: dout  = 8'b11111111; // 1193 : 255 - 0xff
      12'h4AA: dout  = 8'b11111111; // 1194 : 255 - 0xff
      12'h4AB: dout  = 8'b11111111; // 1195 : 255 - 0xff
      12'h4AC: dout  = 8'b11111111; // 1196 : 255 - 0xff
      12'h4AD: dout  = 8'b11111111; // 1197 : 255 - 0xff
      12'h4AE: dout  = 8'b11111111; // 1198 : 255 - 0xff
      12'h4AF: dout  = 8'b11111111; // 1199 : 255 - 0xff
      12'h4B0: dout  = 8'b00111111; // 1200 :  63 - 0x3f -- Background 0x4b
      12'h4B1: dout  = 8'b01111111; // 1201 : 127 - 0x7f
      12'h4B2: dout  = 8'b01111111; // 1202 : 127 - 0x7f
      12'h4B3: dout  = 8'b11111111; // 1203 : 255 - 0xff
      12'h4B4: dout  = 8'b11111111; // 1204 : 255 - 0xff
      12'h4B5: dout  = 8'b11111111; // 1205 : 255 - 0xff
      12'h4B6: dout  = 8'b11111111; // 1206 : 255 - 0xff
      12'h4B7: dout  = 8'b11111111; // 1207 : 255 - 0xff
      12'h4B8: dout  = 8'b00111111; // 1208 :  63 - 0x3f -- plane 1
      12'h4B9: dout  = 8'b01100000; // 1209 :  96 - 0x60
      12'h4BA: dout  = 8'b01000000; // 1210 :  64 - 0x40
      12'h4BB: dout  = 8'b11000000; // 1211 : 192 - 0xc0
      12'h4BC: dout  = 8'b10000000; // 1212 : 128 - 0x80
      12'h4BD: dout  = 8'b10000000; // 1213 : 128 - 0x80
      12'h4BE: dout  = 8'b10000000; // 1214 : 128 - 0x80
      12'h4BF: dout  = 8'b10000000; // 1215 : 128 - 0x80
      12'h4C0: dout  = 8'b11111111; // 1216 : 255 - 0xff -- Background 0x4c
      12'h4C1: dout  = 8'b11111111; // 1217 : 255 - 0xff
      12'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout  = 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout  = 8'b11111111; // 1220 : 255 - 0xff
      12'h4C5: dout  = 8'b11111111; // 1221 : 255 - 0xff
      12'h4C6: dout  = 8'b01111110; // 1222 : 126 - 0x7e
      12'h4C7: dout  = 8'b00111100; // 1223 :  60 - 0x3c
      12'h4C8: dout  = 8'b10000000; // 1224 : 128 - 0x80 -- plane 1
      12'h4C9: dout  = 8'b10000000; // 1225 : 128 - 0x80
      12'h4CA: dout  = 8'b10000000; // 1226 : 128 - 0x80
      12'h4CB: dout  = 8'b10000000; // 1227 : 128 - 0x80
      12'h4CC: dout  = 8'b10000000; // 1228 : 128 - 0x80
      12'h4CD: dout  = 8'b10000001; // 1229 : 129 - 0x81
      12'h4CE: dout  = 8'b01000010; // 1230 :  66 - 0x42
      12'h4CF: dout  = 8'b00111100; // 1231 :  60 - 0x3c
      12'h4D0: dout  = 8'b11111111; // 1232 : 255 - 0xff -- Background 0x4d
      12'h4D1: dout  = 8'b11111111; // 1233 : 255 - 0xff
      12'h4D2: dout  = 8'b11111111; // 1234 : 255 - 0xff
      12'h4D3: dout  = 8'b11111111; // 1235 : 255 - 0xff
      12'h4D4: dout  = 8'b11111111; // 1236 : 255 - 0xff
      12'h4D5: dout  = 8'b11111111; // 1237 : 255 - 0xff
      12'h4D6: dout  = 8'b11111111; // 1238 : 255 - 0xff
      12'h4D7: dout  = 8'b11111111; // 1239 : 255 - 0xff
      12'h4D8: dout  = 8'b11111111; // 1240 : 255 - 0xff -- plane 1
      12'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout  = 8'b11111111; // 1248 : 255 - 0xff -- Background 0x4e
      12'h4E1: dout  = 8'b11111111; // 1249 : 255 - 0xff
      12'h4E2: dout  = 8'b11111111; // 1250 : 255 - 0xff
      12'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      12'h4E4: dout  = 8'b11111111; // 1252 : 255 - 0xff
      12'h4E5: dout  = 8'b11111111; // 1253 : 255 - 0xff
      12'h4E6: dout  = 8'b11111110; // 1254 : 254 - 0xfe
      12'h4E7: dout  = 8'b01111100; // 1255 : 124 - 0x7c
      12'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout  = 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout  = 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout  = 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout  = 8'b00000001; // 1261 :   1 - 0x1
      12'h4EE: dout  = 8'b10000010; // 1262 : 130 - 0x82
      12'h4EF: dout  = 8'b01111100; // 1263 : 124 - 0x7c
      12'h4F0: dout  = 8'b11111111; // 1264 : 255 - 0xff -- Background 0x4f
      12'h4F1: dout  = 8'b11111111; // 1265 : 255 - 0xff
      12'h4F2: dout  = 8'b11111111; // 1266 : 255 - 0xff
      12'h4F3: dout  = 8'b11111111; // 1267 : 255 - 0xff
      12'h4F4: dout  = 8'b11111111; // 1268 : 255 - 0xff
      12'h4F5: dout  = 8'b11111111; // 1269 : 255 - 0xff
      12'h4F6: dout  = 8'b11111110; // 1270 : 254 - 0xfe
      12'h4F7: dout  = 8'b01111100; // 1271 : 124 - 0x7c
      12'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout  = 8'b00000001; // 1277 :   1 - 0x1
      12'h4FE: dout  = 8'b10000011; // 1278 : 131 - 0x83
      12'h4FF: dout  = 8'b11111111; // 1279 : 255 - 0xff
      12'h500: dout  = 8'b11111000; // 1280 : 248 - 0xf8 -- Background 0x50
      12'h501: dout  = 8'b11111100; // 1281 : 252 - 0xfc
      12'h502: dout  = 8'b11111110; // 1282 : 254 - 0xfe
      12'h503: dout  = 8'b11111110; // 1283 : 254 - 0xfe
      12'h504: dout  = 8'b11111111; // 1284 : 255 - 0xff
      12'h505: dout  = 8'b11111111; // 1285 : 255 - 0xff
      12'h506: dout  = 8'b11111111; // 1286 : 255 - 0xff
      12'h507: dout  = 8'b11111111; // 1287 : 255 - 0xff
      12'h508: dout  = 8'b11111000; // 1288 : 248 - 0xf8 -- plane 1
      12'h509: dout  = 8'b00000100; // 1289 :   4 - 0x4
      12'h50A: dout  = 8'b00000010; // 1290 :   2 - 0x2
      12'h50B: dout  = 8'b00000010; // 1291 :   2 - 0x2
      12'h50C: dout  = 8'b00000001; // 1292 :   1 - 0x1
      12'h50D: dout  = 8'b00000001; // 1293 :   1 - 0x1
      12'h50E: dout  = 8'b00000001; // 1294 :   1 - 0x1
      12'h50F: dout  = 8'b00000001; // 1295 :   1 - 0x1
      12'h510: dout  = 8'b11111111; // 1296 : 255 - 0xff -- Background 0x51
      12'h511: dout  = 8'b11111111; // 1297 : 255 - 0xff
      12'h512: dout  = 8'b11111111; // 1298 : 255 - 0xff
      12'h513: dout  = 8'b11111111; // 1299 : 255 - 0xff
      12'h514: dout  = 8'b11111111; // 1300 : 255 - 0xff
      12'h515: dout  = 8'b11111111; // 1301 : 255 - 0xff
      12'h516: dout  = 8'b01111110; // 1302 : 126 - 0x7e
      12'h517: dout  = 8'b00111100; // 1303 :  60 - 0x3c
      12'h518: dout  = 8'b00000001; // 1304 :   1 - 0x1 -- plane 1
      12'h519: dout  = 8'b00000001; // 1305 :   1 - 0x1
      12'h51A: dout  = 8'b00000001; // 1306 :   1 - 0x1
      12'h51B: dout  = 8'b00000001; // 1307 :   1 - 0x1
      12'h51C: dout  = 8'b00000001; // 1308 :   1 - 0x1
      12'h51D: dout  = 8'b10000001; // 1309 : 129 - 0x81
      12'h51E: dout  = 8'b01000010; // 1310 :  66 - 0x42
      12'h51F: dout  = 8'b00111100; // 1311 :  60 - 0x3c
      12'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Background 0x52
      12'h521: dout  = 8'b00001000; // 1313 :   8 - 0x8
      12'h522: dout  = 8'b00001000; // 1314 :   8 - 0x8
      12'h523: dout  = 8'b00001000; // 1315 :   8 - 0x8
      12'h524: dout  = 8'b00010000; // 1316 :  16 - 0x10
      12'h525: dout  = 8'b00010000; // 1317 :  16 - 0x10
      12'h526: dout  = 8'b00010000; // 1318 :  16 - 0x10
      12'h527: dout  = 8'b00000000; // 1319 :   0 - 0x0
      12'h528: dout  = 8'b11111111; // 1320 : 255 - 0xff -- plane 1
      12'h529: dout  = 8'b11111111; // 1321 : 255 - 0xff
      12'h52A: dout  = 8'b11111111; // 1322 : 255 - 0xff
      12'h52B: dout  = 8'b11111111; // 1323 : 255 - 0xff
      12'h52C: dout  = 8'b11111111; // 1324 : 255 - 0xff
      12'h52D: dout  = 8'b11111111; // 1325 : 255 - 0xff
      12'h52E: dout  = 8'b11111111; // 1326 : 255 - 0xff
      12'h52F: dout  = 8'b11111111; // 1327 : 255 - 0xff
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Background 0x53
      12'h531: dout  = 8'b01111111; // 1329 : 127 - 0x7f
      12'h532: dout  = 8'b01111111; // 1330 : 127 - 0x7f
      12'h533: dout  = 8'b01111000; // 1331 : 120 - 0x78
      12'h534: dout  = 8'b01110011; // 1332 : 115 - 0x73
      12'h535: dout  = 8'b01110011; // 1333 : 115 - 0x73
      12'h536: dout  = 8'b01110011; // 1334 : 115 - 0x73
      12'h537: dout  = 8'b01111111; // 1335 : 127 - 0x7f
      12'h538: dout  = 8'b01111111; // 1336 : 127 - 0x7f -- plane 1
      12'h539: dout  = 8'b10000000; // 1337 : 128 - 0x80
      12'h53A: dout  = 8'b10100000; // 1338 : 160 - 0xa0
      12'h53B: dout  = 8'b10000111; // 1339 : 135 - 0x87
      12'h53C: dout  = 8'b10001111; // 1340 : 143 - 0x8f
      12'h53D: dout  = 8'b10001110; // 1341 : 142 - 0x8e
      12'h53E: dout  = 8'b10001110; // 1342 : 142 - 0x8e
      12'h53F: dout  = 8'b10000110; // 1343 : 134 - 0x86
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Background 0x54
      12'h541: dout  = 8'b11111111; // 1345 : 255 - 0xff
      12'h542: dout  = 8'b11111111; // 1346 : 255 - 0xff
      12'h543: dout  = 8'b00111111; // 1347 :  63 - 0x3f
      12'h544: dout  = 8'b10011111; // 1348 : 159 - 0x9f
      12'h545: dout  = 8'b10011111; // 1349 : 159 - 0x9f
      12'h546: dout  = 8'b10011111; // 1350 : 159 - 0x9f
      12'h547: dout  = 8'b00011111; // 1351 :  31 - 0x1f
      12'h548: dout  = 8'b11111110; // 1352 : 254 - 0xfe -- plane 1
      12'h549: dout  = 8'b00000001; // 1353 :   1 - 0x1
      12'h54A: dout  = 8'b00000101; // 1354 :   5 - 0x5
      12'h54B: dout  = 8'b11000001; // 1355 : 193 - 0xc1
      12'h54C: dout  = 8'b11100001; // 1356 : 225 - 0xe1
      12'h54D: dout  = 8'b01110001; // 1357 : 113 - 0x71
      12'h54E: dout  = 8'b01110001; // 1358 : 113 - 0x71
      12'h54F: dout  = 8'b11110001; // 1359 : 241 - 0xf1
      12'h550: dout  = 8'b01111110; // 1360 : 126 - 0x7e -- Background 0x55
      12'h551: dout  = 8'b01111110; // 1361 : 126 - 0x7e
      12'h552: dout  = 8'b01111111; // 1362 : 127 - 0x7f
      12'h553: dout  = 8'b01111110; // 1363 : 126 - 0x7e
      12'h554: dout  = 8'b01111110; // 1364 : 126 - 0x7e
      12'h555: dout  = 8'b01111111; // 1365 : 127 - 0x7f
      12'h556: dout  = 8'b01111111; // 1366 : 127 - 0x7f
      12'h557: dout  = 8'b11111111; // 1367 : 255 - 0xff
      12'h558: dout  = 8'b10000001; // 1368 : 129 - 0x81 -- plane 1
      12'h559: dout  = 8'b10000001; // 1369 : 129 - 0x81
      12'h55A: dout  = 8'b10000000; // 1370 : 128 - 0x80
      12'h55B: dout  = 8'b10000001; // 1371 : 129 - 0x81
      12'h55C: dout  = 8'b10000001; // 1372 : 129 - 0x81
      12'h55D: dout  = 8'b10100000; // 1373 : 160 - 0xa0
      12'h55E: dout  = 8'b10000000; // 1374 : 128 - 0x80
      12'h55F: dout  = 8'b11111111; // 1375 : 255 - 0xff
      12'h560: dout  = 8'b01111111; // 1376 : 127 - 0x7f -- Background 0x56
      12'h561: dout  = 8'b01111111; // 1377 : 127 - 0x7f
      12'h562: dout  = 8'b11111111; // 1378 : 255 - 0xff
      12'h563: dout  = 8'b01111111; // 1379 : 127 - 0x7f
      12'h564: dout  = 8'b01111111; // 1380 : 127 - 0x7f
      12'h565: dout  = 8'b11111111; // 1381 : 255 - 0xff
      12'h566: dout  = 8'b11111111; // 1382 : 255 - 0xff
      12'h567: dout  = 8'b11111111; // 1383 : 255 - 0xff
      12'h568: dout  = 8'b11110001; // 1384 : 241 - 0xf1 -- plane 1
      12'h569: dout  = 8'b11000001; // 1385 : 193 - 0xc1
      12'h56A: dout  = 8'b11000001; // 1386 : 193 - 0xc1
      12'h56B: dout  = 8'b10000001; // 1387 : 129 - 0x81
      12'h56C: dout  = 8'b11000001; // 1388 : 193 - 0xc1
      12'h56D: dout  = 8'b11000101; // 1389 : 197 - 0xc5
      12'h56E: dout  = 8'b00000001; // 1390 :   1 - 0x1
      12'h56F: dout  = 8'b11111111; // 1391 : 255 - 0xff
      12'h570: dout  = 8'b01111111; // 1392 : 127 - 0x7f -- Background 0x57
      12'h571: dout  = 8'b10000000; // 1393 : 128 - 0x80
      12'h572: dout  = 8'b10100000; // 1394 : 160 - 0xa0
      12'h573: dout  = 8'b10000000; // 1395 : 128 - 0x80
      12'h574: dout  = 8'b10000000; // 1396 : 128 - 0x80
      12'h575: dout  = 8'b10000000; // 1397 : 128 - 0x80
      12'h576: dout  = 8'b10000000; // 1398 : 128 - 0x80
      12'h577: dout  = 8'b10000000; // 1399 : 128 - 0x80
      12'h578: dout  = 8'b01111111; // 1400 : 127 - 0x7f -- plane 1
      12'h579: dout  = 8'b11111111; // 1401 : 255 - 0xff
      12'h57A: dout  = 8'b11111111; // 1402 : 255 - 0xff
      12'h57B: dout  = 8'b11111111; // 1403 : 255 - 0xff
      12'h57C: dout  = 8'b11111111; // 1404 : 255 - 0xff
      12'h57D: dout  = 8'b11111111; // 1405 : 255 - 0xff
      12'h57E: dout  = 8'b11111111; // 1406 : 255 - 0xff
      12'h57F: dout  = 8'b11111111; // 1407 : 255 - 0xff
      12'h580: dout  = 8'b11111110; // 1408 : 254 - 0xfe -- Background 0x58
      12'h581: dout  = 8'b00000001; // 1409 :   1 - 0x1
      12'h582: dout  = 8'b00000101; // 1410 :   5 - 0x5
      12'h583: dout  = 8'b00000001; // 1411 :   1 - 0x1
      12'h584: dout  = 8'b00000001; // 1412 :   1 - 0x1
      12'h585: dout  = 8'b00000001; // 1413 :   1 - 0x1
      12'h586: dout  = 8'b00000001; // 1414 :   1 - 0x1
      12'h587: dout  = 8'b00000001; // 1415 :   1 - 0x1
      12'h588: dout  = 8'b11111110; // 1416 : 254 - 0xfe -- plane 1
      12'h589: dout  = 8'b11111111; // 1417 : 255 - 0xff
      12'h58A: dout  = 8'b11111111; // 1418 : 255 - 0xff
      12'h58B: dout  = 8'b11111111; // 1419 : 255 - 0xff
      12'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      12'h58D: dout  = 8'b11111111; // 1421 : 255 - 0xff
      12'h58E: dout  = 8'b11111111; // 1422 : 255 - 0xff
      12'h58F: dout  = 8'b11111111; // 1423 : 255 - 0xff
      12'h590: dout  = 8'b10000000; // 1424 : 128 - 0x80 -- Background 0x59
      12'h591: dout  = 8'b10000000; // 1425 : 128 - 0x80
      12'h592: dout  = 8'b10000000; // 1426 : 128 - 0x80
      12'h593: dout  = 8'b10000000; // 1427 : 128 - 0x80
      12'h594: dout  = 8'b10000000; // 1428 : 128 - 0x80
      12'h595: dout  = 8'b10100000; // 1429 : 160 - 0xa0
      12'h596: dout  = 8'b10000000; // 1430 : 128 - 0x80
      12'h597: dout  = 8'b01111111; // 1431 : 127 - 0x7f
      12'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff -- plane 1
      12'h599: dout  = 8'b11111111; // 1433 : 255 - 0xff
      12'h59A: dout  = 8'b11111111; // 1434 : 255 - 0xff
      12'h59B: dout  = 8'b11111111; // 1435 : 255 - 0xff
      12'h59C: dout  = 8'b11111111; // 1436 : 255 - 0xff
      12'h59D: dout  = 8'b11111111; // 1437 : 255 - 0xff
      12'h59E: dout  = 8'b11111111; // 1438 : 255 - 0xff
      12'h59F: dout  = 8'b01111111; // 1439 : 127 - 0x7f
      12'h5A0: dout  = 8'b00000001; // 1440 :   1 - 0x1 -- Background 0x5a
      12'h5A1: dout  = 8'b00000001; // 1441 :   1 - 0x1
      12'h5A2: dout  = 8'b00000001; // 1442 :   1 - 0x1
      12'h5A3: dout  = 8'b00000001; // 1443 :   1 - 0x1
      12'h5A4: dout  = 8'b00000001; // 1444 :   1 - 0x1
      12'h5A5: dout  = 8'b00000101; // 1445 :   5 - 0x5
      12'h5A6: dout  = 8'b00000001; // 1446 :   1 - 0x1
      12'h5A7: dout  = 8'b11111110; // 1447 : 254 - 0xfe
      12'h5A8: dout  = 8'b11111111; // 1448 : 255 - 0xff -- plane 1
      12'h5A9: dout  = 8'b11111111; // 1449 : 255 - 0xff
      12'h5AA: dout  = 8'b11111111; // 1450 : 255 - 0xff
      12'h5AB: dout  = 8'b11111111; // 1451 : 255 - 0xff
      12'h5AC: dout  = 8'b11111111; // 1452 : 255 - 0xff
      12'h5AD: dout  = 8'b11111111; // 1453 : 255 - 0xff
      12'h5AE: dout  = 8'b11111111; // 1454 : 255 - 0xff
      12'h5AF: dout  = 8'b11111110; // 1455 : 254 - 0xfe
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Background 0x5b
      12'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout  = 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout  = 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout  = 8'b11111100; // 1460 : 252 - 0xfc
      12'h5B5: dout  = 8'b11111110; // 1461 : 254 - 0xfe
      12'h5B6: dout  = 8'b00000111; // 1462 :   7 - 0x7
      12'h5B7: dout  = 8'b00000011; // 1463 :   3 - 0x3
      12'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout  = 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout  = 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout  = 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout  = 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout  = 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout  = 8'b00111000; // 1470 :  56 - 0x38
      12'h5BF: dout  = 8'b01111100; // 1471 : 124 - 0x7c
      12'h5C0: dout  = 8'b00010001; // 1472 :  17 - 0x11 -- Background 0x5c
      12'h5C1: dout  = 8'b00111001; // 1473 :  57 - 0x39
      12'h5C2: dout  = 8'b00010001; // 1474 :  17 - 0x11
      12'h5C3: dout  = 8'b00000001; // 1475 :   1 - 0x1
      12'h5C4: dout  = 8'b00000001; // 1476 :   1 - 0x1
      12'h5C5: dout  = 8'b00000001; // 1477 :   1 - 0x1
      12'h5C6: dout  = 8'b00000001; // 1478 :   1 - 0x1
      12'h5C7: dout  = 8'b00000001; // 1479 :   1 - 0x1
      12'h5C8: dout  = 8'b11111110; // 1480 : 254 - 0xfe -- plane 1
      12'h5C9: dout  = 8'b11111110; // 1481 : 254 - 0xfe
      12'h5CA: dout  = 8'b11111110; // 1482 : 254 - 0xfe
      12'h5CB: dout  = 8'b01111100; // 1483 : 124 - 0x7c
      12'h5CC: dout  = 8'b00111000; // 1484 :  56 - 0x38
      12'h5CD: dout  = 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout  = 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b11101111; // 1488 : 239 - 0xef -- Background 0x5d
      12'h5D1: dout  = 8'b00101000; // 1489 :  40 - 0x28
      12'h5D2: dout  = 8'b00101000; // 1490 :  40 - 0x28
      12'h5D3: dout  = 8'b00101000; // 1491 :  40 - 0x28
      12'h5D4: dout  = 8'b00101000; // 1492 :  40 - 0x28
      12'h5D5: dout  = 8'b00101000; // 1493 :  40 - 0x28
      12'h5D6: dout  = 8'b11101111; // 1494 : 239 - 0xef
      12'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout  = 8'b00100000; // 1496 :  32 - 0x20 -- plane 1
      12'h5D9: dout  = 8'b11100111; // 1497 : 231 - 0xe7
      12'h5DA: dout  = 8'b11100111; // 1498 : 231 - 0xe7
      12'h5DB: dout  = 8'b11100111; // 1499 : 231 - 0xe7
      12'h5DC: dout  = 8'b11100111; // 1500 : 231 - 0xe7
      12'h5DD: dout  = 8'b11100111; // 1501 : 231 - 0xe7
      12'h5DE: dout  = 8'b11101111; // 1502 : 239 - 0xef
      12'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout  = 8'b11111110; // 1504 : 254 - 0xfe -- Background 0x5e
      12'h5E1: dout  = 8'b10000010; // 1505 : 130 - 0x82
      12'h5E2: dout  = 8'b10000010; // 1506 : 130 - 0x82
      12'h5E3: dout  = 8'b10000010; // 1507 : 130 - 0x82
      12'h5E4: dout  = 8'b10000010; // 1508 : 130 - 0x82
      12'h5E5: dout  = 8'b10000010; // 1509 : 130 - 0x82
      12'h5E6: dout  = 8'b11111110; // 1510 : 254 - 0xfe
      12'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout  = 8'b00000010; // 1512 :   2 - 0x2 -- plane 1
      12'h5E9: dout  = 8'b01111110; // 1513 : 126 - 0x7e
      12'h5EA: dout  = 8'b01111110; // 1514 : 126 - 0x7e
      12'h5EB: dout  = 8'b01111110; // 1515 : 126 - 0x7e
      12'h5EC: dout  = 8'b01111110; // 1516 : 126 - 0x7e
      12'h5ED: dout  = 8'b01111110; // 1517 : 126 - 0x7e
      12'h5EE: dout  = 8'b11111110; // 1518 : 254 - 0xfe
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b10000000; // 1520 : 128 - 0x80 -- Background 0x5f
      12'h5F1: dout  = 8'b10000000; // 1521 : 128 - 0x80
      12'h5F2: dout  = 8'b10000000; // 1522 : 128 - 0x80
      12'h5F3: dout  = 8'b10011000; // 1523 : 152 - 0x98
      12'h5F4: dout  = 8'b10011100; // 1524 : 156 - 0x9c
      12'h5F5: dout  = 8'b10001100; // 1525 : 140 - 0x8c
      12'h5F6: dout  = 8'b10000000; // 1526 : 128 - 0x80
      12'h5F7: dout  = 8'b01111111; // 1527 : 127 - 0x7f
      12'h5F8: dout  = 8'b01111111; // 1528 : 127 - 0x7f -- plane 1
      12'h5F9: dout  = 8'b01111111; // 1529 : 127 - 0x7f
      12'h5FA: dout  = 8'b01111111; // 1530 : 127 - 0x7f
      12'h5FB: dout  = 8'b01100111; // 1531 : 103 - 0x67
      12'h5FC: dout  = 8'b01100111; // 1532 : 103 - 0x67
      12'h5FD: dout  = 8'b01111111; // 1533 : 127 - 0x7f
      12'h5FE: dout  = 8'b01111111; // 1534 : 127 - 0x7f
      12'h5FF: dout  = 8'b01111111; // 1535 : 127 - 0x7f
      12'h600: dout  = 8'b11111111; // 1536 : 255 - 0xff -- Background 0x60
      12'h601: dout  = 8'b11111111; // 1537 : 255 - 0xff
      12'h602: dout  = 8'b10000011; // 1538 : 131 - 0x83
      12'h603: dout  = 8'b11110011; // 1539 : 243 - 0xf3
      12'h604: dout  = 8'b11110011; // 1540 : 243 - 0xf3
      12'h605: dout  = 8'b11110011; // 1541 : 243 - 0xf3
      12'h606: dout  = 8'b11110011; // 1542 : 243 - 0xf3
      12'h607: dout  = 8'b11110011; // 1543 : 243 - 0xf3
      12'h608: dout  = 8'b11111111; // 1544 : 255 - 0xff -- plane 1
      12'h609: dout  = 8'b10000000; // 1545 : 128 - 0x80
      12'h60A: dout  = 8'b11111100; // 1546 : 252 - 0xfc
      12'h60B: dout  = 8'b10001100; // 1547 : 140 - 0x8c
      12'h60C: dout  = 8'b10001100; // 1548 : 140 - 0x8c
      12'h60D: dout  = 8'b10001100; // 1549 : 140 - 0x8c
      12'h60E: dout  = 8'b10001100; // 1550 : 140 - 0x8c
      12'h60F: dout  = 8'b10001100; // 1551 : 140 - 0x8c
      12'h610: dout  = 8'b11111111; // 1552 : 255 - 0xff -- Background 0x61
      12'h611: dout  = 8'b11111111; // 1553 : 255 - 0xff
      12'h612: dout  = 8'b11110000; // 1554 : 240 - 0xf0
      12'h613: dout  = 8'b11110110; // 1555 : 246 - 0xf6
      12'h614: dout  = 8'b11110110; // 1556 : 246 - 0xf6
      12'h615: dout  = 8'b11110110; // 1557 : 246 - 0xf6
      12'h616: dout  = 8'b11110110; // 1558 : 246 - 0xf6
      12'h617: dout  = 8'b11110110; // 1559 : 246 - 0xf6
      12'h618: dout  = 8'b11111111; // 1560 : 255 - 0xff -- plane 1
      12'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout  = 8'b00001111; // 1562 :  15 - 0xf
      12'h61B: dout  = 8'b00001001; // 1563 :   9 - 0x9
      12'h61C: dout  = 8'b00001001; // 1564 :   9 - 0x9
      12'h61D: dout  = 8'b00001001; // 1565 :   9 - 0x9
      12'h61E: dout  = 8'b00001001; // 1566 :   9 - 0x9
      12'h61F: dout  = 8'b00001001; // 1567 :   9 - 0x9
      12'h620: dout  = 8'b11111111; // 1568 : 255 - 0xff -- Background 0x62
      12'h621: dout  = 8'b11111111; // 1569 : 255 - 0xff
      12'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout  = 8'b11111111; // 1576 : 255 - 0xff -- plane 1
      12'h629: dout  = 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout  = 8'b11111111; // 1578 : 255 - 0xff
      12'h62B: dout  = 8'b11111111; // 1579 : 255 - 0xff
      12'h62C: dout  = 8'b11111111; // 1580 : 255 - 0xff
      12'h62D: dout  = 8'b11111111; // 1581 : 255 - 0xff
      12'h62E: dout  = 8'b11111111; // 1582 : 255 - 0xff
      12'h62F: dout  = 8'b11111111; // 1583 : 255 - 0xff
      12'h630: dout  = 8'b11111111; // 1584 : 255 - 0xff -- Background 0x63
      12'h631: dout  = 8'b11111111; // 1585 : 255 - 0xff
      12'h632: dout  = 8'b00000001; // 1586 :   1 - 0x1
      12'h633: dout  = 8'b01010111; // 1587 :  87 - 0x57
      12'h634: dout  = 8'b00101111; // 1588 :  47 - 0x2f
      12'h635: dout  = 8'b01010111; // 1589 :  87 - 0x57
      12'h636: dout  = 8'b00101111; // 1590 :  47 - 0x2f
      12'h637: dout  = 8'b01010111; // 1591 :  87 - 0x57
      12'h638: dout  = 8'b11111111; // 1592 : 255 - 0xff -- plane 1
      12'h639: dout  = 8'b00000001; // 1593 :   1 - 0x1
      12'h63A: dout  = 8'b11111111; // 1594 : 255 - 0xff
      12'h63B: dout  = 8'b10101001; // 1595 : 169 - 0xa9
      12'h63C: dout  = 8'b11010001; // 1596 : 209 - 0xd1
      12'h63D: dout  = 8'b10101001; // 1597 : 169 - 0xa9
      12'h63E: dout  = 8'b11010001; // 1598 : 209 - 0xd1
      12'h63F: dout  = 8'b10101001; // 1599 : 169 - 0xa9
      12'h640: dout  = 8'b11110011; // 1600 : 243 - 0xf3 -- Background 0x64
      12'h641: dout  = 8'b11110011; // 1601 : 243 - 0xf3
      12'h642: dout  = 8'b11110011; // 1602 : 243 - 0xf3
      12'h643: dout  = 8'b11110011; // 1603 : 243 - 0xf3
      12'h644: dout  = 8'b11110011; // 1604 : 243 - 0xf3
      12'h645: dout  = 8'b11110011; // 1605 : 243 - 0xf3
      12'h646: dout  = 8'b11111111; // 1606 : 255 - 0xff
      12'h647: dout  = 8'b00111111; // 1607 :  63 - 0x3f
      12'h648: dout  = 8'b10001100; // 1608 : 140 - 0x8c -- plane 1
      12'h649: dout  = 8'b10001100; // 1609 : 140 - 0x8c
      12'h64A: dout  = 8'b10001100; // 1610 : 140 - 0x8c
      12'h64B: dout  = 8'b10001100; // 1611 : 140 - 0x8c
      12'h64C: dout  = 8'b10001100; // 1612 : 140 - 0x8c
      12'h64D: dout  = 8'b10001100; // 1613 : 140 - 0x8c
      12'h64E: dout  = 8'b11111111; // 1614 : 255 - 0xff
      12'h64F: dout  = 8'b00111111; // 1615 :  63 - 0x3f
      12'h650: dout  = 8'b11110110; // 1616 : 246 - 0xf6 -- Background 0x65
      12'h651: dout  = 8'b11110110; // 1617 : 246 - 0xf6
      12'h652: dout  = 8'b11110110; // 1618 : 246 - 0xf6
      12'h653: dout  = 8'b11110110; // 1619 : 246 - 0xf6
      12'h654: dout  = 8'b11110110; // 1620 : 246 - 0xf6
      12'h655: dout  = 8'b11110110; // 1621 : 246 - 0xf6
      12'h656: dout  = 8'b11111111; // 1622 : 255 - 0xff
      12'h657: dout  = 8'b11111111; // 1623 : 255 - 0xff
      12'h658: dout  = 8'b00001001; // 1624 :   9 - 0x9 -- plane 1
      12'h659: dout  = 8'b00001001; // 1625 :   9 - 0x9
      12'h65A: dout  = 8'b00001001; // 1626 :   9 - 0x9
      12'h65B: dout  = 8'b00001001; // 1627 :   9 - 0x9
      12'h65C: dout  = 8'b00001001; // 1628 :   9 - 0x9
      12'h65D: dout  = 8'b00001001; // 1629 :   9 - 0x9
      12'h65E: dout  = 8'b11111111; // 1630 : 255 - 0xff
      12'h65F: dout  = 8'b11111111; // 1631 : 255 - 0xff
      12'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Background 0x66
      12'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout  = 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout  = 8'b11111111; // 1638 : 255 - 0xff
      12'h667: dout  = 8'b11111111; // 1639 : 255 - 0xff
      12'h668: dout  = 8'b11111111; // 1640 : 255 - 0xff -- plane 1
      12'h669: dout  = 8'b11111111; // 1641 : 255 - 0xff
      12'h66A: dout  = 8'b11111111; // 1642 : 255 - 0xff
      12'h66B: dout  = 8'b11111111; // 1643 : 255 - 0xff
      12'h66C: dout  = 8'b11111111; // 1644 : 255 - 0xff
      12'h66D: dout  = 8'b11111111; // 1645 : 255 - 0xff
      12'h66E: dout  = 8'b11111111; // 1646 : 255 - 0xff
      12'h66F: dout  = 8'b11111111; // 1647 : 255 - 0xff
      12'h670: dout  = 8'b00101111; // 1648 :  47 - 0x2f -- Background 0x67
      12'h671: dout  = 8'b01010111; // 1649 :  87 - 0x57
      12'h672: dout  = 8'b00101111; // 1650 :  47 - 0x2f
      12'h673: dout  = 8'b01010111; // 1651 :  87 - 0x57
      12'h674: dout  = 8'b00101111; // 1652 :  47 - 0x2f
      12'h675: dout  = 8'b01010111; // 1653 :  87 - 0x57
      12'h676: dout  = 8'b11111111; // 1654 : 255 - 0xff
      12'h677: dout  = 8'b11111100; // 1655 : 252 - 0xfc
      12'h678: dout  = 8'b11010001; // 1656 : 209 - 0xd1 -- plane 1
      12'h679: dout  = 8'b10101001; // 1657 : 169 - 0xa9
      12'h67A: dout  = 8'b11010001; // 1658 : 209 - 0xd1
      12'h67B: dout  = 8'b10101001; // 1659 : 169 - 0xa9
      12'h67C: dout  = 8'b11010001; // 1660 : 209 - 0xd1
      12'h67D: dout  = 8'b10101001; // 1661 : 169 - 0xa9
      12'h67E: dout  = 8'b11111111; // 1662 : 255 - 0xff
      12'h67F: dout  = 8'b11111100; // 1663 : 252 - 0xfc
      12'h680: dout  = 8'b00111100; // 1664 :  60 - 0x3c -- Background 0x68
      12'h681: dout  = 8'b00111100; // 1665 :  60 - 0x3c
      12'h682: dout  = 8'b00111100; // 1666 :  60 - 0x3c
      12'h683: dout  = 8'b00111100; // 1667 :  60 - 0x3c
      12'h684: dout  = 8'b00111100; // 1668 :  60 - 0x3c
      12'h685: dout  = 8'b00111100; // 1669 :  60 - 0x3c
      12'h686: dout  = 8'b00111100; // 1670 :  60 - 0x3c
      12'h687: dout  = 8'b00111100; // 1671 :  60 - 0x3c
      12'h688: dout  = 8'b00100011; // 1672 :  35 - 0x23 -- plane 1
      12'h689: dout  = 8'b00100011; // 1673 :  35 - 0x23
      12'h68A: dout  = 8'b00100011; // 1674 :  35 - 0x23
      12'h68B: dout  = 8'b00100011; // 1675 :  35 - 0x23
      12'h68C: dout  = 8'b00100011; // 1676 :  35 - 0x23
      12'h68D: dout  = 8'b00100011; // 1677 :  35 - 0x23
      12'h68E: dout  = 8'b00100011; // 1678 :  35 - 0x23
      12'h68F: dout  = 8'b00100011; // 1679 :  35 - 0x23
      12'h690: dout  = 8'b11111011; // 1680 : 251 - 0xfb -- Background 0x69
      12'h691: dout  = 8'b11111011; // 1681 : 251 - 0xfb
      12'h692: dout  = 8'b11111011; // 1682 : 251 - 0xfb
      12'h693: dout  = 8'b11111011; // 1683 : 251 - 0xfb
      12'h694: dout  = 8'b11111011; // 1684 : 251 - 0xfb
      12'h695: dout  = 8'b11111011; // 1685 : 251 - 0xfb
      12'h696: dout  = 8'b11111011; // 1686 : 251 - 0xfb
      12'h697: dout  = 8'b11111011; // 1687 : 251 - 0xfb
      12'h698: dout  = 8'b00000100; // 1688 :   4 - 0x4 -- plane 1
      12'h699: dout  = 8'b00000100; // 1689 :   4 - 0x4
      12'h69A: dout  = 8'b00000100; // 1690 :   4 - 0x4
      12'h69B: dout  = 8'b00000100; // 1691 :   4 - 0x4
      12'h69C: dout  = 8'b00000100; // 1692 :   4 - 0x4
      12'h69D: dout  = 8'b00000100; // 1693 :   4 - 0x4
      12'h69E: dout  = 8'b00000100; // 1694 :   4 - 0x4
      12'h69F: dout  = 8'b00000100; // 1695 :   4 - 0x4
      12'h6A0: dout  = 8'b10111100; // 1696 : 188 - 0xbc -- Background 0x6a
      12'h6A1: dout  = 8'b01011100; // 1697 :  92 - 0x5c
      12'h6A2: dout  = 8'b10111100; // 1698 : 188 - 0xbc
      12'h6A3: dout  = 8'b01011100; // 1699 :  92 - 0x5c
      12'h6A4: dout  = 8'b10111100; // 1700 : 188 - 0xbc
      12'h6A5: dout  = 8'b01011100; // 1701 :  92 - 0x5c
      12'h6A6: dout  = 8'b10111100; // 1702 : 188 - 0xbc
      12'h6A7: dout  = 8'b01011100; // 1703 :  92 - 0x5c
      12'h6A8: dout  = 8'b01000100; // 1704 :  68 - 0x44 -- plane 1
      12'h6A9: dout  = 8'b10100100; // 1705 : 164 - 0xa4
      12'h6AA: dout  = 8'b01000100; // 1706 :  68 - 0x44
      12'h6AB: dout  = 8'b10100100; // 1707 : 164 - 0xa4
      12'h6AC: dout  = 8'b01000100; // 1708 :  68 - 0x44
      12'h6AD: dout  = 8'b10100100; // 1709 : 164 - 0xa4
      12'h6AE: dout  = 8'b01000100; // 1710 :  68 - 0x44
      12'h6AF: dout  = 8'b10100100; // 1711 : 164 - 0xa4
      12'h6B0: dout  = 8'b00011111; // 1712 :  31 - 0x1f -- Background 0x6b
      12'h6B1: dout  = 8'b00100000; // 1713 :  32 - 0x20
      12'h6B2: dout  = 8'b01000000; // 1714 :  64 - 0x40
      12'h6B3: dout  = 8'b01000000; // 1715 :  64 - 0x40
      12'h6B4: dout  = 8'b10000000; // 1716 : 128 - 0x80
      12'h6B5: dout  = 8'b10000000; // 1717 : 128 - 0x80
      12'h6B6: dout  = 8'b10000000; // 1718 : 128 - 0x80
      12'h6B7: dout  = 8'b10000001; // 1719 : 129 - 0x81
      12'h6B8: dout  = 8'b00011111; // 1720 :  31 - 0x1f -- plane 1
      12'h6B9: dout  = 8'b00111111; // 1721 :  63 - 0x3f
      12'h6BA: dout  = 8'b01111111; // 1722 : 127 - 0x7f
      12'h6BB: dout  = 8'b01111111; // 1723 : 127 - 0x7f
      12'h6BC: dout  = 8'b11111111; // 1724 : 255 - 0xff
      12'h6BD: dout  = 8'b11111111; // 1725 : 255 - 0xff
      12'h6BE: dout  = 8'b11111111; // 1726 : 255 - 0xff
      12'h6BF: dout  = 8'b11111110; // 1727 : 254 - 0xfe
      12'h6C0: dout  = 8'b11111111; // 1728 : 255 - 0xff -- Background 0x6c
      12'h6C1: dout  = 8'b10000000; // 1729 : 128 - 0x80
      12'h6C2: dout  = 8'b10000000; // 1730 : 128 - 0x80
      12'h6C3: dout  = 8'b11000000; // 1731 : 192 - 0xc0
      12'h6C4: dout  = 8'b11111111; // 1732 : 255 - 0xff
      12'h6C5: dout  = 8'b11111111; // 1733 : 255 - 0xff
      12'h6C6: dout  = 8'b11111110; // 1734 : 254 - 0xfe
      12'h6C7: dout  = 8'b11111110; // 1735 : 254 - 0xfe
      12'h6C8: dout  = 8'b11111111; // 1736 : 255 - 0xff -- plane 1
      12'h6C9: dout  = 8'b01111111; // 1737 : 127 - 0x7f
      12'h6CA: dout  = 8'b01111111; // 1738 : 127 - 0x7f
      12'h6CB: dout  = 8'b00111111; // 1739 :  63 - 0x3f
      12'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout  = 8'b00000001; // 1742 :   1 - 0x1
      12'h6CF: dout  = 8'b00000001; // 1743 :   1 - 0x1
      12'h6D0: dout  = 8'b11111111; // 1744 : 255 - 0xff -- Background 0x6d
      12'h6D1: dout  = 8'b01111111; // 1745 : 127 - 0x7f
      12'h6D2: dout  = 8'b01111111; // 1746 : 127 - 0x7f
      12'h6D3: dout  = 8'b11111111; // 1747 : 255 - 0xff
      12'h6D4: dout  = 8'b11111111; // 1748 : 255 - 0xff
      12'h6D5: dout  = 8'b00000111; // 1749 :   7 - 0x7
      12'h6D6: dout  = 8'b00000011; // 1750 :   3 - 0x3
      12'h6D7: dout  = 8'b00000011; // 1751 :   3 - 0x3
      12'h6D8: dout  = 8'b11111111; // 1752 : 255 - 0xff -- plane 1
      12'h6D9: dout  = 8'b10000000; // 1753 : 128 - 0x80
      12'h6DA: dout  = 8'b10000000; // 1754 : 128 - 0x80
      12'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout  = 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout  = 8'b11111000; // 1757 : 248 - 0xf8
      12'h6DE: dout  = 8'b11111100; // 1758 : 252 - 0xfc
      12'h6DF: dout  = 8'b11111100; // 1759 : 252 - 0xfc
      12'h6E0: dout  = 8'b11111111; // 1760 : 255 - 0xff -- Background 0x6e
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout  = 8'b10000001; // 1765 : 129 - 0x81
      12'h6E6: dout  = 8'b11000011; // 1766 : 195 - 0xc3
      12'h6E7: dout  = 8'b11111111; // 1767 : 255 - 0xff
      12'h6E8: dout  = 8'b11111111; // 1768 : 255 - 0xff -- plane 1
      12'h6E9: dout  = 8'b11111111; // 1769 : 255 - 0xff
      12'h6EA: dout  = 8'b11111111; // 1770 : 255 - 0xff
      12'h6EB: dout  = 8'b11111111; // 1771 : 255 - 0xff
      12'h6EC: dout  = 8'b11111111; // 1772 : 255 - 0xff
      12'h6ED: dout  = 8'b01111110; // 1773 : 126 - 0x7e
      12'h6EE: dout  = 8'b00111100; // 1774 :  60 - 0x3c
      12'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout  = 8'b11111000; // 1776 : 248 - 0xf8 -- Background 0x6f
      12'h6F1: dout  = 8'b11111100; // 1777 : 252 - 0xfc
      12'h6F2: dout  = 8'b11111110; // 1778 : 254 - 0xfe
      12'h6F3: dout  = 8'b11111110; // 1779 : 254 - 0xfe
      12'h6F4: dout  = 8'b11100011; // 1780 : 227 - 0xe3
      12'h6F5: dout  = 8'b11000001; // 1781 : 193 - 0xc1
      12'h6F6: dout  = 8'b10000001; // 1782 : 129 - 0x81
      12'h6F7: dout  = 8'b10000001; // 1783 : 129 - 0x81
      12'h6F8: dout  = 8'b11111000; // 1784 : 248 - 0xf8 -- plane 1
      12'h6F9: dout  = 8'b00000100; // 1785 :   4 - 0x4
      12'h6FA: dout  = 8'b00000010; // 1786 :   2 - 0x2
      12'h6FB: dout  = 8'b00000010; // 1787 :   2 - 0x2
      12'h6FC: dout  = 8'b00011101; // 1788 :  29 - 0x1d
      12'h6FD: dout  = 8'b00111111; // 1789 :  63 - 0x3f
      12'h6FE: dout  = 8'b01111111; // 1790 : 127 - 0x7f
      12'h6FF: dout  = 8'b01111111; // 1791 : 127 - 0x7f
      12'h700: dout  = 8'b10000011; // 1792 : 131 - 0x83 -- Background 0x70
      12'h701: dout  = 8'b11111111; // 1793 : 255 - 0xff
      12'h702: dout  = 8'b11111111; // 1794 : 255 - 0xff
      12'h703: dout  = 8'b11111111; // 1795 : 255 - 0xff
      12'h704: dout  = 8'b11111111; // 1796 : 255 - 0xff
      12'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout  = 8'b01111111; // 1798 : 127 - 0x7f
      12'h707: dout  = 8'b00011111; // 1799 :  31 - 0x1f
      12'h708: dout  = 8'b11111100; // 1800 : 252 - 0xfc -- plane 1
      12'h709: dout  = 8'b10000000; // 1801 : 128 - 0x80
      12'h70A: dout  = 8'b10000000; // 1802 : 128 - 0x80
      12'h70B: dout  = 8'b10000000; // 1803 : 128 - 0x80
      12'h70C: dout  = 8'b10000000; // 1804 : 128 - 0x80
      12'h70D: dout  = 8'b10000000; // 1805 : 128 - 0x80
      12'h70E: dout  = 8'b01100000; // 1806 :  96 - 0x60
      12'h70F: dout  = 8'b00011111; // 1807 :  31 - 0x1f
      12'h710: dout  = 8'b11111100; // 1808 : 252 - 0xfc -- Background 0x71
      12'h711: dout  = 8'b11111100; // 1809 : 252 - 0xfc
      12'h712: dout  = 8'b11111100; // 1810 : 252 - 0xfc
      12'h713: dout  = 8'b11111100; // 1811 : 252 - 0xfc
      12'h714: dout  = 8'b11111110; // 1812 : 254 - 0xfe
      12'h715: dout  = 8'b11111110; // 1813 : 254 - 0xfe
      12'h716: dout  = 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout  = 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout  = 8'b00000011; // 1816 :   3 - 0x3 -- plane 1
      12'h719: dout  = 8'b00000011; // 1817 :   3 - 0x3
      12'h71A: dout  = 8'b00000011; // 1818 :   3 - 0x3
      12'h71B: dout  = 8'b00000011; // 1819 :   3 - 0x3
      12'h71C: dout  = 8'b00000001; // 1820 :   1 - 0x1
      12'h71D: dout  = 8'b00000001; // 1821 :   1 - 0x1
      12'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout  = 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout  = 8'b00000001; // 1824 :   1 - 0x1 -- Background 0x72
      12'h721: dout  = 8'b00000001; // 1825 :   1 - 0x1
      12'h722: dout  = 8'b00000001; // 1826 :   1 - 0x1
      12'h723: dout  = 8'b00000001; // 1827 :   1 - 0x1
      12'h724: dout  = 8'b00000011; // 1828 :   3 - 0x3
      12'h725: dout  = 8'b00000011; // 1829 :   3 - 0x3
      12'h726: dout  = 8'b00000111; // 1830 :   7 - 0x7
      12'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout  = 8'b11111110; // 1832 : 254 - 0xfe -- plane 1
      12'h729: dout  = 8'b11111110; // 1833 : 254 - 0xfe
      12'h72A: dout  = 8'b11111110; // 1834 : 254 - 0xfe
      12'h72B: dout  = 8'b11111110; // 1835 : 254 - 0xfe
      12'h72C: dout  = 8'b11111100; // 1836 : 252 - 0xfc
      12'h72D: dout  = 8'b11111100; // 1837 : 252 - 0xfc
      12'h72E: dout  = 8'b11111000; // 1838 : 248 - 0xf8
      12'h72F: dout  = 8'b11111111; // 1839 : 255 - 0xff
      12'h730: dout  = 8'b11111111; // 1840 : 255 - 0xff -- Background 0x73
      12'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout  = 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout  = 8'b11111111; // 1843 : 255 - 0xff
      12'h734: dout  = 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout  = 8'b11111111; // 1845 : 255 - 0xff
      12'h736: dout  = 8'b11111111; // 1846 : 255 - 0xff
      12'h737: dout  = 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- plane 1
      12'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout  = 8'b11111111; // 1855 : 255 - 0xff
      12'h740: dout  = 8'b10000001; // 1856 : 129 - 0x81 -- Background 0x74
      12'h741: dout  = 8'b11000001; // 1857 : 193 - 0xc1
      12'h742: dout  = 8'b11100011; // 1858 : 227 - 0xe3
      12'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout  = 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout  = 8'b11111110; // 1863 : 254 - 0xfe
      12'h748: dout  = 8'b01111111; // 1864 : 127 - 0x7f -- plane 1
      12'h749: dout  = 8'b00111111; // 1865 :  63 - 0x3f
      12'h74A: dout  = 8'b00011101; // 1866 :  29 - 0x1d
      12'h74B: dout  = 8'b00000001; // 1867 :   1 - 0x1
      12'h74C: dout  = 8'b00000001; // 1868 :   1 - 0x1
      12'h74D: dout  = 8'b00000001; // 1869 :   1 - 0x1
      12'h74E: dout  = 8'b00000011; // 1870 :   3 - 0x3
      12'h74F: dout  = 8'b11111110; // 1871 : 254 - 0xfe
      12'h750: dout  = 8'b11111111; // 1872 : 255 - 0xff -- Background 0x75
      12'h751: dout  = 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout  = 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout  = 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout  = 8'b11111011; // 1877 : 251 - 0xfb
      12'h756: dout  = 8'b10110101; // 1878 : 181 - 0xb5
      12'h757: dout  = 8'b11001110; // 1879 : 206 - 0xce
      12'h758: dout  = 8'b10000000; // 1880 : 128 - 0x80 -- plane 1
      12'h759: dout  = 8'b10000000; // 1881 : 128 - 0x80
      12'h75A: dout  = 8'b10000000; // 1882 : 128 - 0x80
      12'h75B: dout  = 8'b10000000; // 1883 : 128 - 0x80
      12'h75C: dout  = 8'b10000000; // 1884 : 128 - 0x80
      12'h75D: dout  = 8'b10000100; // 1885 : 132 - 0x84
      12'h75E: dout  = 8'b11001010; // 1886 : 202 - 0xca
      12'h75F: dout  = 8'b10110001; // 1887 : 177 - 0xb1
      12'h760: dout  = 8'b11111111; // 1888 : 255 - 0xff -- Background 0x76
      12'h761: dout  = 8'b11111111; // 1889 : 255 - 0xff
      12'h762: dout  = 8'b11111111; // 1890 : 255 - 0xff
      12'h763: dout  = 8'b11111111; // 1891 : 255 - 0xff
      12'h764: dout  = 8'b11111111; // 1892 : 255 - 0xff
      12'h765: dout  = 8'b11011111; // 1893 : 223 - 0xdf
      12'h766: dout  = 8'b10101101; // 1894 : 173 - 0xad
      12'h767: dout  = 8'b01110011; // 1895 : 115 - 0x73
      12'h768: dout  = 8'b00000001; // 1896 :   1 - 0x1 -- plane 1
      12'h769: dout  = 8'b00000001; // 1897 :   1 - 0x1
      12'h76A: dout  = 8'b00000001; // 1898 :   1 - 0x1
      12'h76B: dout  = 8'b00000001; // 1899 :   1 - 0x1
      12'h76C: dout  = 8'b00000001; // 1900 :   1 - 0x1
      12'h76D: dout  = 8'b00100001; // 1901 :  33 - 0x21
      12'h76E: dout  = 8'b01010011; // 1902 :  83 - 0x53
      12'h76F: dout  = 8'b10001101; // 1903 : 141 - 0x8d
      12'h770: dout  = 8'b01110111; // 1904 : 119 - 0x77 -- Background 0x77
      12'h771: dout  = 8'b01110111; // 1905 : 119 - 0x77
      12'h772: dout  = 8'b01110111; // 1906 : 119 - 0x77
      12'h773: dout  = 8'b01110111; // 1907 : 119 - 0x77
      12'h774: dout  = 8'b01110111; // 1908 : 119 - 0x77
      12'h775: dout  = 8'b01110111; // 1909 : 119 - 0x77
      12'h776: dout  = 8'b01110111; // 1910 : 119 - 0x77
      12'h777: dout  = 8'b01110111; // 1911 : 119 - 0x77
      12'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- plane 1
      12'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout  = 8'b01110111; // 1916 : 119 - 0x77
      12'h77D: dout  = 8'b11111111; // 1917 : 255 - 0xff
      12'h77E: dout  = 8'b11111111; // 1918 : 255 - 0xff
      12'h77F: dout  = 8'b11111111; // 1919 : 255 - 0xff
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Background 0x78
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- plane 1
      12'h789: dout  = 8'b11111111; // 1929 : 255 - 0xff
      12'h78A: dout  = 8'b11111111; // 1930 : 255 - 0xff
      12'h78B: dout  = 8'b11111111; // 1931 : 255 - 0xff
      12'h78C: dout  = 8'b11111111; // 1932 : 255 - 0xff
      12'h78D: dout  = 8'b11111111; // 1933 : 255 - 0xff
      12'h78E: dout  = 8'b11111111; // 1934 : 255 - 0xff
      12'h78F: dout  = 8'b11111111; // 1935 : 255 - 0xff
      12'h790: dout  = 8'b01110111; // 1936 : 119 - 0x77 -- Background 0x79
      12'h791: dout  = 8'b01110111; // 1937 : 119 - 0x77
      12'h792: dout  = 8'b01110111; // 1938 : 119 - 0x77
      12'h793: dout  = 8'b01110111; // 1939 : 119 - 0x77
      12'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout  = 8'b11111111; // 1944 : 255 - 0xff -- plane 1
      12'h799: dout  = 8'b11111111; // 1945 : 255 - 0xff
      12'h79A: dout  = 8'b11111111; // 1946 : 255 - 0xff
      12'h79B: dout  = 8'b01110111; // 1947 : 119 - 0x77
      12'h79C: dout  = 8'b01110111; // 1948 : 119 - 0x77
      12'h79D: dout  = 8'b01110111; // 1949 : 119 - 0x77
      12'h79E: dout  = 8'b01110111; // 1950 : 119 - 0x77
      12'h79F: dout  = 8'b01110111; // 1951 : 119 - 0x77
      12'h7A0: dout  = 8'b00000001; // 1952 :   1 - 0x1 -- Background 0x7a
      12'h7A1: dout  = 8'b00000001; // 1953 :   1 - 0x1
      12'h7A2: dout  = 8'b00000001; // 1954 :   1 - 0x1
      12'h7A3: dout  = 8'b00011001; // 1955 :  25 - 0x19
      12'h7A4: dout  = 8'b00011101; // 1956 :  29 - 0x1d
      12'h7A5: dout  = 8'b00001101; // 1957 :  13 - 0xd
      12'h7A6: dout  = 8'b00000001; // 1958 :   1 - 0x1
      12'h7A7: dout  = 8'b11111110; // 1959 : 254 - 0xfe
      12'h7A8: dout  = 8'b11111111; // 1960 : 255 - 0xff -- plane 1
      12'h7A9: dout  = 8'b11111111; // 1961 : 255 - 0xff
      12'h7AA: dout  = 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout  = 8'b11100111; // 1963 : 231 - 0xe7
      12'h7AC: dout  = 8'b11100111; // 1964 : 231 - 0xe7
      12'h7AD: dout  = 8'b11111111; // 1965 : 255 - 0xff
      12'h7AE: dout  = 8'b11111111; // 1966 : 255 - 0xff
      12'h7AF: dout  = 8'b11111110; // 1967 : 254 - 0xfe
      12'h7B0: dout  = 8'b00100000; // 1968 :  32 - 0x20 -- Background 0x7b
      12'h7B1: dout  = 8'b01111000; // 1969 : 120 - 0x78
      12'h7B2: dout  = 8'b01111111; // 1970 : 127 - 0x7f
      12'h7B3: dout  = 8'b11111110; // 1971 : 254 - 0xfe
      12'h7B4: dout  = 8'b11111110; // 1972 : 254 - 0xfe
      12'h7B5: dout  = 8'b11111110; // 1973 : 254 - 0xfe
      12'h7B6: dout  = 8'b11111110; // 1974 : 254 - 0xfe
      12'h7B7: dout  = 8'b11111110; // 1975 : 254 - 0xfe
      12'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- plane 1
      12'h7B9: dout  = 8'b00100001; // 1977 :  33 - 0x21
      12'h7BA: dout  = 8'b00100001; // 1978 :  33 - 0x21
      12'h7BB: dout  = 8'b01000001; // 1979 :  65 - 0x41
      12'h7BC: dout  = 8'b01000001; // 1980 :  65 - 0x41
      12'h7BD: dout  = 8'b01000001; // 1981 :  65 - 0x41
      12'h7BE: dout  = 8'b01000001; // 1982 :  65 - 0x41
      12'h7BF: dout  = 8'b01000001; // 1983 :  65 - 0x41
      12'h7C0: dout  = 8'b00000100; // 1984 :   4 - 0x4 -- Background 0x7c
      12'h7C1: dout  = 8'b10011010; // 1985 : 154 - 0x9a
      12'h7C2: dout  = 8'b11111010; // 1986 : 250 - 0xfa
      12'h7C3: dout  = 8'b11111101; // 1987 : 253 - 0xfd
      12'h7C4: dout  = 8'b11111101; // 1988 : 253 - 0xfd
      12'h7C5: dout  = 8'b11111101; // 1989 : 253 - 0xfd
      12'h7C6: dout  = 8'b11111101; // 1990 : 253 - 0xfd
      12'h7C7: dout  = 8'b11111101; // 1991 : 253 - 0xfd
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout  = 8'b10000000; // 1993 : 128 - 0x80
      12'h7CA: dout  = 8'b10000000; // 1994 : 128 - 0x80
      12'h7CB: dout  = 8'b10000000; // 1995 : 128 - 0x80
      12'h7CC: dout  = 8'b10000000; // 1996 : 128 - 0x80
      12'h7CD: dout  = 8'b10000000; // 1997 : 128 - 0x80
      12'h7CE: dout  = 8'b10000000; // 1998 : 128 - 0x80
      12'h7CF: dout  = 8'b10000000; // 1999 : 128 - 0x80
      12'h7D0: dout  = 8'b01111110; // 2000 : 126 - 0x7e -- Background 0x7d
      12'h7D1: dout  = 8'b00111000; // 2001 :  56 - 0x38
      12'h7D2: dout  = 8'b00100001; // 2002 :  33 - 0x21
      12'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout  = 8'b00000001; // 2004 :   1 - 0x1
      12'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout  = 8'b00000001; // 2006 :   1 - 0x1
      12'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout  = 8'b00100001; // 2008 :  33 - 0x21 -- plane 1
      12'h7D9: dout  = 8'b00100001; // 2009 :  33 - 0x21
      12'h7DA: dout  = 8'b00000001; // 2010 :   1 - 0x1
      12'h7DB: dout  = 8'b00000001; // 2011 :   1 - 0x1
      12'h7DC: dout  = 8'b00000001; // 2012 :   1 - 0x1
      12'h7DD: dout  = 8'b00000001; // 2013 :   1 - 0x1
      12'h7DE: dout  = 8'b00000001; // 2014 :   1 - 0x1
      12'h7DF: dout  = 8'b00000001; // 2015 :   1 - 0x1
      12'h7E0: dout  = 8'b11111010; // 2016 : 250 - 0xfa -- Background 0x7e
      12'h7E1: dout  = 8'b10001010; // 2017 : 138 - 0x8a
      12'h7E2: dout  = 8'b10000100; // 2018 : 132 - 0x84
      12'h7E3: dout  = 8'b10000000; // 2019 : 128 - 0x80
      12'h7E4: dout  = 8'b10000000; // 2020 : 128 - 0x80
      12'h7E5: dout  = 8'b10000000; // 2021 : 128 - 0x80
      12'h7E6: dout  = 8'b10000000; // 2022 : 128 - 0x80
      12'h7E7: dout  = 8'b10000000; // 2023 : 128 - 0x80
      12'h7E8: dout  = 8'b10000000; // 2024 : 128 - 0x80 -- plane 1
      12'h7E9: dout  = 8'b10000000; // 2025 : 128 - 0x80
      12'h7EA: dout  = 8'b10000000; // 2026 : 128 - 0x80
      12'h7EB: dout  = 8'b10000000; // 2027 : 128 - 0x80
      12'h7EC: dout  = 8'b10000000; // 2028 : 128 - 0x80
      12'h7ED: dout  = 8'b10000000; // 2029 : 128 - 0x80
      12'h7EE: dout  = 8'b10000000; // 2030 : 128 - 0x80
      12'h7EF: dout  = 8'b10000000; // 2031 : 128 - 0x80
      12'h7F0: dout  = 8'b00000010; // 2032 :   2 - 0x2 -- Background 0x7f
      12'h7F1: dout  = 8'b00000100; // 2033 :   4 - 0x4
      12'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout  = 8'b00010000; // 2035 :  16 - 0x10
      12'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout  = 8'b01000000; // 2037 :  64 - 0x40
      12'h7F6: dout  = 8'b10000000; // 2038 : 128 - 0x80
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000001; // 2040 :   1 - 0x1 -- plane 1
      12'h7F9: dout  = 8'b00000001; // 2041 :   1 - 0x1
      12'h7FA: dout  = 8'b00000110; // 2042 :   6 - 0x6
      12'h7FB: dout  = 8'b00001000; // 2043 :   8 - 0x8
      12'h7FC: dout  = 8'b00011000; // 2044 :  24 - 0x18
      12'h7FD: dout  = 8'b00100000; // 2045 :  32 - 0x20
      12'h7FE: dout  = 8'b00100000; // 2046 :  32 - 0x20
      12'h7FF: dout  = 8'b11000000; // 2047 : 192 - 0xc0
      12'h800: dout  = 8'b00001011; // 2048 :  11 - 0xb -- Background 0x80
      12'h801: dout  = 8'b00001011; // 2049 :  11 - 0xb
      12'h802: dout  = 8'b00111011; // 2050 :  59 - 0x3b
      12'h803: dout  = 8'b00001011; // 2051 :  11 - 0xb
      12'h804: dout  = 8'b11111011; // 2052 : 251 - 0xfb
      12'h805: dout  = 8'b00001011; // 2053 :  11 - 0xb
      12'h806: dout  = 8'b00001011; // 2054 :  11 - 0xb
      12'h807: dout  = 8'b00001010; // 2055 :  10 - 0xa
      12'h808: dout  = 8'b00000100; // 2056 :   4 - 0x4 -- plane 1
      12'h809: dout  = 8'b00000100; // 2057 :   4 - 0x4
      12'h80A: dout  = 8'b11000100; // 2058 : 196 - 0xc4
      12'h80B: dout  = 8'b11110100; // 2059 : 244 - 0xf4
      12'h80C: dout  = 8'b11110100; // 2060 : 244 - 0xf4
      12'h80D: dout  = 8'b00000100; // 2061 :   4 - 0x4
      12'h80E: dout  = 8'b00000100; // 2062 :   4 - 0x4
      12'h80F: dout  = 8'b00000101; // 2063 :   5 - 0x5
      12'h810: dout  = 8'b10010000; // 2064 : 144 - 0x90 -- Background 0x81
      12'h811: dout  = 8'b00010000; // 2065 :  16 - 0x10
      12'h812: dout  = 8'b00011111; // 2066 :  31 - 0x1f
      12'h813: dout  = 8'b00010000; // 2067 :  16 - 0x10
      12'h814: dout  = 8'b00011111; // 2068 :  31 - 0x1f
      12'h815: dout  = 8'b00010000; // 2069 :  16 - 0x10
      12'h816: dout  = 8'b00010000; // 2070 :  16 - 0x10
      12'h817: dout  = 8'b10010000; // 2071 : 144 - 0x90
      12'h818: dout  = 8'b01110000; // 2072 : 112 - 0x70 -- plane 1
      12'h819: dout  = 8'b11110000; // 2073 : 240 - 0xf0
      12'h81A: dout  = 8'b11110000; // 2074 : 240 - 0xf0
      12'h81B: dout  = 8'b11111111; // 2075 : 255 - 0xff
      12'h81C: dout  = 8'b11111111; // 2076 : 255 - 0xff
      12'h81D: dout  = 8'b11110000; // 2077 : 240 - 0xf0
      12'h81E: dout  = 8'b11110000; // 2078 : 240 - 0xf0
      12'h81F: dout  = 8'b01110000; // 2079 : 112 - 0x70
      12'h820: dout  = 8'b00111111; // 2080 :  63 - 0x3f -- Background 0x82
      12'h821: dout  = 8'b01111000; // 2081 : 120 - 0x78
      12'h822: dout  = 8'b11100111; // 2082 : 231 - 0xe7
      12'h823: dout  = 8'b11001111; // 2083 : 207 - 0xcf
      12'h824: dout  = 8'b01011000; // 2084 :  88 - 0x58
      12'h825: dout  = 8'b01011000; // 2085 :  88 - 0x58
      12'h826: dout  = 8'b01010000; // 2086 :  80 - 0x50
      12'h827: dout  = 8'b10010000; // 2087 : 144 - 0x90
      12'h828: dout  = 8'b11000000; // 2088 : 192 - 0xc0 -- plane 1
      12'h829: dout  = 8'b10000111; // 2089 : 135 - 0x87
      12'h82A: dout  = 8'b00011000; // 2090 :  24 - 0x18
      12'h82B: dout  = 8'b10110000; // 2091 : 176 - 0xb0
      12'h82C: dout  = 8'b11100111; // 2092 : 231 - 0xe7
      12'h82D: dout  = 8'b11100111; // 2093 : 231 - 0xe7
      12'h82E: dout  = 8'b11101111; // 2094 : 239 - 0xef
      12'h82F: dout  = 8'b11101111; // 2095 : 239 - 0xef
      12'h830: dout  = 8'b10110000; // 2096 : 176 - 0xb0 -- Background 0x83
      12'h831: dout  = 8'b11111100; // 2097 : 252 - 0xfc
      12'h832: dout  = 8'b11100010; // 2098 : 226 - 0xe2
      12'h833: dout  = 8'b11000001; // 2099 : 193 - 0xc1
      12'h834: dout  = 8'b11000001; // 2100 : 193 - 0xc1
      12'h835: dout  = 8'b10000011; // 2101 : 131 - 0x83
      12'h836: dout  = 8'b10001111; // 2102 : 143 - 0x8f
      12'h837: dout  = 8'b01111110; // 2103 : 126 - 0x7e
      12'h838: dout  = 8'b01101111; // 2104 : 111 - 0x6f -- plane 1
      12'h839: dout  = 8'b01000011; // 2105 :  67 - 0x43
      12'h83A: dout  = 8'b01011101; // 2106 :  93 - 0x5d
      12'h83B: dout  = 8'b00111111; // 2107 :  63 - 0x3f
      12'h83C: dout  = 8'b00111111; // 2108 :  63 - 0x3f
      12'h83D: dout  = 8'b01111111; // 2109 : 127 - 0x7f
      12'h83E: dout  = 8'b01111111; // 2110 : 127 - 0x7f
      12'h83F: dout  = 8'b11111111; // 2111 : 255 - 0xff
      12'h840: dout  = 8'b11111110; // 2112 : 254 - 0xfe -- Background 0x84
      12'h841: dout  = 8'b00000011; // 2113 :   3 - 0x3
      12'h842: dout  = 8'b00001111; // 2114 :  15 - 0xf
      12'h843: dout  = 8'b10010001; // 2115 : 145 - 0x91
      12'h844: dout  = 8'b01110000; // 2116 : 112 - 0x70
      12'h845: dout  = 8'b01100000; // 2117 :  96 - 0x60
      12'h846: dout  = 8'b00100000; // 2118 :  32 - 0x20
      12'h847: dout  = 8'b00110001; // 2119 :  49 - 0x31
      12'h848: dout  = 8'b00000011; // 2120 :   3 - 0x3 -- plane 1
      12'h849: dout  = 8'b11111111; // 2121 : 255 - 0xff
      12'h84A: dout  = 8'b11110001; // 2122 : 241 - 0xf1
      12'h84B: dout  = 8'b01101110; // 2123 : 110 - 0x6e
      12'h84C: dout  = 8'b11001111; // 2124 : 207 - 0xcf
      12'h84D: dout  = 8'b11011111; // 2125 : 223 - 0xdf
      12'h84E: dout  = 8'b11111111; // 2126 : 255 - 0xff
      12'h84F: dout  = 8'b11111111; // 2127 : 255 - 0xff
      12'h850: dout  = 8'b00111111; // 2128 :  63 - 0x3f -- Background 0x85
      12'h851: dout  = 8'b00111111; // 2129 :  63 - 0x3f
      12'h852: dout  = 8'b00011101; // 2130 :  29 - 0x1d
      12'h853: dout  = 8'b00111001; // 2131 :  57 - 0x39
      12'h854: dout  = 8'b01111011; // 2132 : 123 - 0x7b
      12'h855: dout  = 8'b11110011; // 2133 : 243 - 0xf3
      12'h856: dout  = 8'b10000110; // 2134 : 134 - 0x86
      12'h857: dout  = 8'b11111110; // 2135 : 254 - 0xfe
      12'h858: dout  = 8'b11111101; // 2136 : 253 - 0xfd -- plane 1
      12'h859: dout  = 8'b11111011; // 2137 : 251 - 0xfb
      12'h85A: dout  = 8'b11111011; // 2138 : 251 - 0xfb
      12'h85B: dout  = 8'b11110111; // 2139 : 247 - 0xf7
      12'h85C: dout  = 8'b11110111; // 2140 : 247 - 0xf7
      12'h85D: dout  = 8'b00001111; // 2141 :  15 - 0xf
      12'h85E: dout  = 8'b01111111; // 2142 : 127 - 0x7f
      12'h85F: dout  = 8'b11111111; // 2143 : 255 - 0xff
      12'h860: dout  = 8'b11111111; // 2144 : 255 - 0xff -- Background 0x86
      12'h861: dout  = 8'b11111111; // 2145 : 255 - 0xff
      12'h862: dout  = 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout  = 8'b11111111; // 2147 : 255 - 0xff
      12'h864: dout  = 8'b11111111; // 2148 : 255 - 0xff
      12'h865: dout  = 8'b10000000; // 2149 : 128 - 0x80
      12'h866: dout  = 8'b10000000; // 2150 : 128 - 0x80
      12'h867: dout  = 8'b11111111; // 2151 : 255 - 0xff
      12'h868: dout  = 8'b11111111; // 2152 : 255 - 0xff -- plane 1
      12'h869: dout  = 8'b10000000; // 2153 : 128 - 0x80
      12'h86A: dout  = 8'b10000000; // 2154 : 128 - 0x80
      12'h86B: dout  = 8'b10000000; // 2155 : 128 - 0x80
      12'h86C: dout  = 8'b10000000; // 2156 : 128 - 0x80
      12'h86D: dout  = 8'b11111111; // 2157 : 255 - 0xff
      12'h86E: dout  = 8'b11111111; // 2158 : 255 - 0xff
      12'h86F: dout  = 8'b10000000; // 2159 : 128 - 0x80
      12'h870: dout  = 8'b11111110; // 2160 : 254 - 0xfe -- Background 0x87
      12'h871: dout  = 8'b11111111; // 2161 : 255 - 0xff
      12'h872: dout  = 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout  = 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout  = 8'b11111111; // 2164 : 255 - 0xff
      12'h875: dout  = 8'b00000011; // 2165 :   3 - 0x3
      12'h876: dout  = 8'b00000011; // 2166 :   3 - 0x3
      12'h877: dout  = 8'b11111111; // 2167 : 255 - 0xff
      12'h878: dout  = 8'b11111110; // 2168 : 254 - 0xfe -- plane 1
      12'h879: dout  = 8'b00000011; // 2169 :   3 - 0x3
      12'h87A: dout  = 8'b00000011; // 2170 :   3 - 0x3
      12'h87B: dout  = 8'b00000011; // 2171 :   3 - 0x3
      12'h87C: dout  = 8'b00000011; // 2172 :   3 - 0x3
      12'h87D: dout  = 8'b11111111; // 2173 : 255 - 0xff
      12'h87E: dout  = 8'b11111111; // 2174 : 255 - 0xff
      12'h87F: dout  = 8'b00000011; // 2175 :   3 - 0x3
      12'h880: dout  = 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x88
      12'h881: dout  = 8'b11111111; // 2177 : 255 - 0xff
      12'h882: dout  = 8'b11111111; // 2178 : 255 - 0xff
      12'h883: dout  = 8'b11111111; // 2179 : 255 - 0xff
      12'h884: dout  = 8'b11111111; // 2180 : 255 - 0xff
      12'h885: dout  = 8'b11111111; // 2181 : 255 - 0xff
      12'h886: dout  = 8'b00000000; // 2182 :   0 - 0x0
      12'h887: dout  = 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout  = 8'b11111111; // 2185 : 255 - 0xff
      12'h88A: dout  = 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout  = 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout  = 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout  = 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout  = 8'b11111111; // 2190 : 255 - 0xff
      12'h88F: dout  = 8'b11111111; // 2191 : 255 - 0xff
      12'h890: dout  = 8'b00111100; // 2192 :  60 - 0x3c -- Background 0x89
      12'h891: dout  = 8'b11111100; // 2193 : 252 - 0xfc
      12'h892: dout  = 8'b11111100; // 2194 : 252 - 0xfc
      12'h893: dout  = 8'b11111100; // 2195 : 252 - 0xfc
      12'h894: dout  = 8'b11111100; // 2196 : 252 - 0xfc
      12'h895: dout  = 8'b11111100; // 2197 : 252 - 0xfc
      12'h896: dout  = 8'b00000100; // 2198 :   4 - 0x4
      12'h897: dout  = 8'b00000100; // 2199 :   4 - 0x4
      12'h898: dout  = 8'b00100011; // 2200 :  35 - 0x23 -- plane 1
      12'h899: dout  = 8'b11110011; // 2201 : 243 - 0xf3
      12'h89A: dout  = 8'b00001011; // 2202 :  11 - 0xb
      12'h89B: dout  = 8'b00001011; // 2203 :  11 - 0xb
      12'h89C: dout  = 8'b00001011; // 2204 :  11 - 0xb
      12'h89D: dout  = 8'b00000111; // 2205 :   7 - 0x7
      12'h89E: dout  = 8'b11111111; // 2206 : 255 - 0xff
      12'h89F: dout  = 8'b11111111; // 2207 : 255 - 0xff
      12'h8A0: dout  = 8'b11111111; // 2208 : 255 - 0xff -- Background 0x8a
      12'h8A1: dout  = 8'b11111111; // 2209 : 255 - 0xff
      12'h8A2: dout  = 8'b11111111; // 2210 : 255 - 0xff
      12'h8A3: dout  = 8'b11111111; // 2211 : 255 - 0xff
      12'h8A4: dout  = 8'b10000000; // 2212 : 128 - 0x80
      12'h8A5: dout  = 8'b11111111; // 2213 : 255 - 0xff
      12'h8A6: dout  = 8'b11111111; // 2214 : 255 - 0xff
      12'h8A7: dout  = 8'b11111111; // 2215 : 255 - 0xff
      12'h8A8: dout  = 8'b10000000; // 2216 : 128 - 0x80 -- plane 1
      12'h8A9: dout  = 8'b10000000; // 2217 : 128 - 0x80
      12'h8AA: dout  = 8'b10000000; // 2218 : 128 - 0x80
      12'h8AB: dout  = 8'b10000000; // 2219 : 128 - 0x80
      12'h8AC: dout  = 8'b11111111; // 2220 : 255 - 0xff
      12'h8AD: dout  = 8'b10000000; // 2221 : 128 - 0x80
      12'h8AE: dout  = 8'b10000000; // 2222 : 128 - 0x80
      12'h8AF: dout  = 8'b10000000; // 2223 : 128 - 0x80
      12'h8B0: dout  = 8'b11111111; // 2224 : 255 - 0xff -- Background 0x8b
      12'h8B1: dout  = 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout  = 8'b11111111; // 2226 : 255 - 0xff
      12'h8B3: dout  = 8'b11111111; // 2227 : 255 - 0xff
      12'h8B4: dout  = 8'b00000011; // 2228 :   3 - 0x3
      12'h8B5: dout  = 8'b11111111; // 2229 : 255 - 0xff
      12'h8B6: dout  = 8'b11111111; // 2230 : 255 - 0xff
      12'h8B7: dout  = 8'b11111111; // 2231 : 255 - 0xff
      12'h8B8: dout  = 8'b00000011; // 2232 :   3 - 0x3 -- plane 1
      12'h8B9: dout  = 8'b00000011; // 2233 :   3 - 0x3
      12'h8BA: dout  = 8'b00000011; // 2234 :   3 - 0x3
      12'h8BB: dout  = 8'b00000011; // 2235 :   3 - 0x3
      12'h8BC: dout  = 8'b11111111; // 2236 : 255 - 0xff
      12'h8BD: dout  = 8'b00000011; // 2237 :   3 - 0x3
      12'h8BE: dout  = 8'b00000011; // 2238 :   3 - 0x3
      12'h8BF: dout  = 8'b00000011; // 2239 :   3 - 0x3
      12'h8C0: dout  = 8'b11111111; // 2240 : 255 - 0xff -- Background 0x8c
      12'h8C1: dout  = 8'b11111111; // 2241 : 255 - 0xff
      12'h8C2: dout  = 8'b11111111; // 2242 : 255 - 0xff
      12'h8C3: dout  = 8'b11111111; // 2243 : 255 - 0xff
      12'h8C4: dout  = 8'b11111111; // 2244 : 255 - 0xff
      12'h8C5: dout  = 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout  = 8'b11111111; // 2246 : 255 - 0xff
      12'h8C7: dout  = 8'b11111111; // 2247 : 255 - 0xff
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout  = 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout  = 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout  = 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout  = 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout  = 8'b11111111; // 2253 : 255 - 0xff
      12'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b11111100; // 2256 : 252 - 0xfc -- Background 0x8d
      12'h8D1: dout  = 8'b11111100; // 2257 : 252 - 0xfc
      12'h8D2: dout  = 8'b11111110; // 2258 : 254 - 0xfe
      12'h8D3: dout  = 8'b11111110; // 2259 : 254 - 0xfe
      12'h8D4: dout  = 8'b11111110; // 2260 : 254 - 0xfe
      12'h8D5: dout  = 8'b00000010; // 2261 :   2 - 0x2
      12'h8D6: dout  = 8'b11111110; // 2262 : 254 - 0xfe
      12'h8D7: dout  = 8'b11111110; // 2263 : 254 - 0xfe
      12'h8D8: dout  = 8'b00000111; // 2264 :   7 - 0x7 -- plane 1
      12'h8D9: dout  = 8'b00000111; // 2265 :   7 - 0x7
      12'h8DA: dout  = 8'b00000011; // 2266 :   3 - 0x3
      12'h8DB: dout  = 8'b00000011; // 2267 :   3 - 0x3
      12'h8DC: dout  = 8'b00000011; // 2268 :   3 - 0x3
      12'h8DD: dout  = 8'b11111111; // 2269 : 255 - 0xff
      12'h8DE: dout  = 8'b00000011; // 2270 :   3 - 0x3
      12'h8DF: dout  = 8'b00000011; // 2271 :   3 - 0x3
      12'h8E0: dout  = 8'b11111111; // 2272 : 255 - 0xff -- Background 0x8e
      12'h8E1: dout  = 8'b10000000; // 2273 : 128 - 0x80
      12'h8E2: dout  = 8'b10000000; // 2274 : 128 - 0x80
      12'h8E3: dout  = 8'b10000000; // 2275 : 128 - 0x80
      12'h8E4: dout  = 8'b10000000; // 2276 : 128 - 0x80
      12'h8E5: dout  = 8'b10000000; // 2277 : 128 - 0x80
      12'h8E6: dout  = 8'b10000000; // 2278 : 128 - 0x80
      12'h8E7: dout  = 8'b10000000; // 2279 : 128 - 0x80
      12'h8E8: dout  = 8'b10000000; // 2280 : 128 - 0x80 -- plane 1
      12'h8E9: dout  = 8'b11111111; // 2281 : 255 - 0xff
      12'h8EA: dout  = 8'b11111111; // 2282 : 255 - 0xff
      12'h8EB: dout  = 8'b11111111; // 2283 : 255 - 0xff
      12'h8EC: dout  = 8'b11111111; // 2284 : 255 - 0xff
      12'h8ED: dout  = 8'b11111111; // 2285 : 255 - 0xff
      12'h8EE: dout  = 8'b11111111; // 2286 : 255 - 0xff
      12'h8EF: dout  = 8'b11111111; // 2287 : 255 - 0xff
      12'h8F0: dout  = 8'b11111111; // 2288 : 255 - 0xff -- Background 0x8f
      12'h8F1: dout  = 8'b00000011; // 2289 :   3 - 0x3
      12'h8F2: dout  = 8'b00000011; // 2290 :   3 - 0x3
      12'h8F3: dout  = 8'b00000011; // 2291 :   3 - 0x3
      12'h8F4: dout  = 8'b00000011; // 2292 :   3 - 0x3
      12'h8F5: dout  = 8'b00000011; // 2293 :   3 - 0x3
      12'h8F6: dout  = 8'b00000011; // 2294 :   3 - 0x3
      12'h8F7: dout  = 8'b00000011; // 2295 :   3 - 0x3
      12'h8F8: dout  = 8'b00000011; // 2296 :   3 - 0x3 -- plane 1
      12'h8F9: dout  = 8'b11111111; // 2297 : 255 - 0xff
      12'h8FA: dout  = 8'b11111111; // 2298 : 255 - 0xff
      12'h8FB: dout  = 8'b11111111; // 2299 : 255 - 0xff
      12'h8FC: dout  = 8'b11111111; // 2300 : 255 - 0xff
      12'h8FD: dout  = 8'b11111111; // 2301 : 255 - 0xff
      12'h8FE: dout  = 8'b11111111; // 2302 : 255 - 0xff
      12'h8FF: dout  = 8'b11111111; // 2303 : 255 - 0xff
      12'h900: dout  = 8'b00000010; // 2304 :   2 - 0x2 -- Background 0x90
      12'h901: dout  = 8'b00000010; // 2305 :   2 - 0x2
      12'h902: dout  = 8'b00000010; // 2306 :   2 - 0x2
      12'h903: dout  = 8'b00000010; // 2307 :   2 - 0x2
      12'h904: dout  = 8'b00000010; // 2308 :   2 - 0x2
      12'h905: dout  = 8'b00000010; // 2309 :   2 - 0x2
      12'h906: dout  = 8'b00000100; // 2310 :   4 - 0x4
      12'h907: dout  = 8'b00000100; // 2311 :   4 - 0x4
      12'h908: dout  = 8'b11111111; // 2312 : 255 - 0xff -- plane 1
      12'h909: dout  = 8'b11111111; // 2313 : 255 - 0xff
      12'h90A: dout  = 8'b11111111; // 2314 : 255 - 0xff
      12'h90B: dout  = 8'b11111111; // 2315 : 255 - 0xff
      12'h90C: dout  = 8'b11111111; // 2316 : 255 - 0xff
      12'h90D: dout  = 8'b11111111; // 2317 : 255 - 0xff
      12'h90E: dout  = 8'b11111111; // 2318 : 255 - 0xff
      12'h90F: dout  = 8'b11111111; // 2319 : 255 - 0xff
      12'h910: dout  = 8'b10000000; // 2320 : 128 - 0x80 -- Background 0x91
      12'h911: dout  = 8'b10000000; // 2321 : 128 - 0x80
      12'h912: dout  = 8'b10101010; // 2322 : 170 - 0xaa
      12'h913: dout  = 8'b11010101; // 2323 : 213 - 0xd5
      12'h914: dout  = 8'b10101010; // 2324 : 170 - 0xaa
      12'h915: dout  = 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout  = 8'b11111111; // 2326 : 255 - 0xff
      12'h917: dout  = 8'b11111111; // 2327 : 255 - 0xff
      12'h918: dout  = 8'b11111111; // 2328 : 255 - 0xff -- plane 1
      12'h919: dout  = 8'b11111111; // 2329 : 255 - 0xff
      12'h91A: dout  = 8'b11010101; // 2330 : 213 - 0xd5
      12'h91B: dout  = 8'b10101010; // 2331 : 170 - 0xaa
      12'h91C: dout  = 8'b11010101; // 2332 : 213 - 0xd5
      12'h91D: dout  = 8'b10000000; // 2333 : 128 - 0x80
      12'h91E: dout  = 8'b10000000; // 2334 : 128 - 0x80
      12'h91F: dout  = 8'b11111111; // 2335 : 255 - 0xff
      12'h920: dout  = 8'b00000011; // 2336 :   3 - 0x3 -- Background 0x92
      12'h921: dout  = 8'b00000011; // 2337 :   3 - 0x3
      12'h922: dout  = 8'b10101011; // 2338 : 171 - 0xab
      12'h923: dout  = 8'b01010111; // 2339 :  87 - 0x57
      12'h924: dout  = 8'b10101011; // 2340 : 171 - 0xab
      12'h925: dout  = 8'b11111111; // 2341 : 255 - 0xff
      12'h926: dout  = 8'b11111111; // 2342 : 255 - 0xff
      12'h927: dout  = 8'b11111110; // 2343 : 254 - 0xfe
      12'h928: dout  = 8'b11111111; // 2344 : 255 - 0xff -- plane 1
      12'h929: dout  = 8'b11111111; // 2345 : 255 - 0xff
      12'h92A: dout  = 8'b01010111; // 2346 :  87 - 0x57
      12'h92B: dout  = 8'b10101011; // 2347 : 171 - 0xab
      12'h92C: dout  = 8'b01010111; // 2348 :  87 - 0x57
      12'h92D: dout  = 8'b00000011; // 2349 :   3 - 0x3
      12'h92E: dout  = 8'b00000011; // 2350 :   3 - 0x3
      12'h92F: dout  = 8'b11111110; // 2351 : 254 - 0xfe
      12'h930: dout  = 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x93
      12'h931: dout  = 8'b01010101; // 2353 :  85 - 0x55
      12'h932: dout  = 8'b10101010; // 2354 : 170 - 0xaa
      12'h933: dout  = 8'b01010101; // 2355 :  85 - 0x55
      12'h934: dout  = 8'b11111111; // 2356 : 255 - 0xff
      12'h935: dout  = 8'b11111111; // 2357 : 255 - 0xff
      12'h936: dout  = 8'b11111111; // 2358 : 255 - 0xff
      12'h937: dout  = 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout  = 8'b11111111; // 2360 : 255 - 0xff -- plane 1
      12'h939: dout  = 8'b10101010; // 2361 : 170 - 0xaa
      12'h93A: dout  = 8'b01010101; // 2362 :  85 - 0x55
      12'h93B: dout  = 8'b10101010; // 2363 : 170 - 0xaa
      12'h93C: dout  = 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout  = 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout  = 8'b11111111; // 2366 : 255 - 0xff
      12'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout  = 8'b00000100; // 2368 :   4 - 0x4 -- Background 0x94
      12'h941: dout  = 8'b01010100; // 2369 :  84 - 0x54
      12'h942: dout  = 8'b10101100; // 2370 : 172 - 0xac
      12'h943: dout  = 8'b01011100; // 2371 :  92 - 0x5c
      12'h944: dout  = 8'b11111100; // 2372 : 252 - 0xfc
      12'h945: dout  = 8'b11111100; // 2373 : 252 - 0xfc
      12'h946: dout  = 8'b11111100; // 2374 : 252 - 0xfc
      12'h947: dout  = 8'b00111100; // 2375 :  60 - 0x3c
      12'h948: dout  = 8'b11111111; // 2376 : 255 - 0xff -- plane 1
      12'h949: dout  = 8'b10101111; // 2377 : 175 - 0xaf
      12'h94A: dout  = 8'b01010111; // 2378 :  87 - 0x57
      12'h94B: dout  = 8'b10101011; // 2379 : 171 - 0xab
      12'h94C: dout  = 8'b00001011; // 2380 :  11 - 0xb
      12'h94D: dout  = 8'b00001011; // 2381 :  11 - 0xb
      12'h94E: dout  = 8'b11110011; // 2382 : 243 - 0xf3
      12'h94F: dout  = 8'b00100011; // 2383 :  35 - 0x23
      12'h950: dout  = 8'b00111111; // 2384 :  63 - 0x3f -- Background 0x95
      12'h951: dout  = 8'b00111111; // 2385 :  63 - 0x3f
      12'h952: dout  = 8'b00111111; // 2386 :  63 - 0x3f
      12'h953: dout  = 8'b00111111; // 2387 :  63 - 0x3f
      12'h954: dout  = 8'b00000000; // 2388 :   0 - 0x0
      12'h955: dout  = 8'b00000000; // 2389 :   0 - 0x0
      12'h956: dout  = 8'b00000000; // 2390 :   0 - 0x0
      12'h957: dout  = 8'b11111111; // 2391 : 255 - 0xff
      12'h958: dout  = 8'b11111111; // 2392 : 255 - 0xff -- plane 1
      12'h959: dout  = 8'b11111111; // 2393 : 255 - 0xff
      12'h95A: dout  = 8'b11111111; // 2394 : 255 - 0xff
      12'h95B: dout  = 8'b11111111; // 2395 : 255 - 0xff
      12'h95C: dout  = 8'b11111111; // 2396 : 255 - 0xff
      12'h95D: dout  = 8'b11111111; // 2397 : 255 - 0xff
      12'h95E: dout  = 8'b11111111; // 2398 : 255 - 0xff
      12'h95F: dout  = 8'b11111111; // 2399 : 255 - 0xff
      12'h960: dout  = 8'b01111110; // 2400 : 126 - 0x7e -- Background 0x96
      12'h961: dout  = 8'b01111100; // 2401 : 124 - 0x7c
      12'h962: dout  = 8'b01111100; // 2402 : 124 - 0x7c
      12'h963: dout  = 8'b01111000; // 2403 : 120 - 0x78
      12'h964: dout  = 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout  = 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout  = 8'b11111111; // 2407 : 255 - 0xff
      12'h968: dout  = 8'b11111111; // 2408 : 255 - 0xff -- plane 1
      12'h969: dout  = 8'b11111111; // 2409 : 255 - 0xff
      12'h96A: dout  = 8'b11111111; // 2410 : 255 - 0xff
      12'h96B: dout  = 8'b11111111; // 2411 : 255 - 0xff
      12'h96C: dout  = 8'b11111111; // 2412 : 255 - 0xff
      12'h96D: dout  = 8'b11111111; // 2413 : 255 - 0xff
      12'h96E: dout  = 8'b11111111; // 2414 : 255 - 0xff
      12'h96F: dout  = 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout  = 8'b00011111; // 2416 :  31 - 0x1f -- Background 0x97
      12'h971: dout  = 8'b00001111; // 2417 :  15 - 0xf
      12'h972: dout  = 8'b00001111; // 2418 :  15 - 0xf
      12'h973: dout  = 8'b00000111; // 2419 :   7 - 0x7
      12'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout  = 8'b11111111; // 2423 : 255 - 0xff
      12'h978: dout  = 8'b11111111; // 2424 : 255 - 0xff -- plane 1
      12'h979: dout  = 8'b11111111; // 2425 : 255 - 0xff
      12'h97A: dout  = 8'b11111111; // 2426 : 255 - 0xff
      12'h97B: dout  = 8'b11111111; // 2427 : 255 - 0xff
      12'h97C: dout  = 8'b11111111; // 2428 : 255 - 0xff
      12'h97D: dout  = 8'b11111111; // 2429 : 255 - 0xff
      12'h97E: dout  = 8'b11111111; // 2430 : 255 - 0xff
      12'h97F: dout  = 8'b11111111; // 2431 : 255 - 0xff
      12'h980: dout  = 8'b11111110; // 2432 : 254 - 0xfe -- Background 0x98
      12'h981: dout  = 8'b11111100; // 2433 : 252 - 0xfc
      12'h982: dout  = 8'b11111100; // 2434 : 252 - 0xfc
      12'h983: dout  = 8'b11111000; // 2435 : 248 - 0xf8
      12'h984: dout  = 8'b00000000; // 2436 :   0 - 0x0
      12'h985: dout  = 8'b00000000; // 2437 :   0 - 0x0
      12'h986: dout  = 8'b00000000; // 2438 :   0 - 0x0
      12'h987: dout  = 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout  = 8'b11111111; // 2440 : 255 - 0xff -- plane 1
      12'h989: dout  = 8'b11111111; // 2441 : 255 - 0xff
      12'h98A: dout  = 8'b11111111; // 2442 : 255 - 0xff
      12'h98B: dout  = 8'b11111111; // 2443 : 255 - 0xff
      12'h98C: dout  = 8'b11111111; // 2444 : 255 - 0xff
      12'h98D: dout  = 8'b11111111; // 2445 : 255 - 0xff
      12'h98E: dout  = 8'b11111111; // 2446 : 255 - 0xff
      12'h98F: dout  = 8'b11111111; // 2447 : 255 - 0xff
      12'h990: dout  = 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x99
      12'h991: dout  = 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout  = 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout  = 8'b11111111; // 2452 : 255 - 0xff
      12'h995: dout  = 8'b11111111; // 2453 : 255 - 0xff
      12'h996: dout  = 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout  = 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout  = 8'b00000000; // 2456 :   0 - 0x0 -- plane 1
      12'h999: dout  = 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout  = 8'b00000000; // 2458 :   0 - 0x0
      12'h99B: dout  = 8'b00000000; // 2459 :   0 - 0x0
      12'h99C: dout  = 8'b00000000; // 2460 :   0 - 0x0
      12'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout  = 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout  = 8'b00011000; // 2464 :  24 - 0x18 -- Background 0x9a
      12'h9A1: dout  = 8'b00011000; // 2465 :  24 - 0x18
      12'h9A2: dout  = 8'b00011000; // 2466 :  24 - 0x18
      12'h9A3: dout  = 8'b00011000; // 2467 :  24 - 0x18
      12'h9A4: dout  = 8'b00011000; // 2468 :  24 - 0x18
      12'h9A5: dout  = 8'b00011000; // 2469 :  24 - 0x18
      12'h9A6: dout  = 8'b00011000; // 2470 :  24 - 0x18
      12'h9A7: dout  = 8'b00011000; // 2471 :  24 - 0x18
      12'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout  = 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout  = 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout  = 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout  = 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout  = 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout  = 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout  = 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout  = 8'b00000111; // 2480 :   7 - 0x7 -- Background 0x9b
      12'h9B1: dout  = 8'b00011111; // 2481 :  31 - 0x1f
      12'h9B2: dout  = 8'b00111111; // 2482 :  63 - 0x3f
      12'h9B3: dout  = 8'b11111111; // 2483 : 255 - 0xff
      12'h9B4: dout  = 8'b01111111; // 2484 : 127 - 0x7f
      12'h9B5: dout  = 8'b01111111; // 2485 : 127 - 0x7f
      12'h9B6: dout  = 8'b11111111; // 2486 : 255 - 0xff
      12'h9B7: dout  = 8'b11111111; // 2487 : 255 - 0xff
      12'h9B8: dout  = 8'b11111111; // 2488 : 255 - 0xff -- plane 1
      12'h9B9: dout  = 8'b11111111; // 2489 : 255 - 0xff
      12'h9BA: dout  = 8'b11111111; // 2490 : 255 - 0xff
      12'h9BB: dout  = 8'b11111111; // 2491 : 255 - 0xff
      12'h9BC: dout  = 8'b11111111; // 2492 : 255 - 0xff
      12'h9BD: dout  = 8'b11111111; // 2493 : 255 - 0xff
      12'h9BE: dout  = 8'b11111111; // 2494 : 255 - 0xff
      12'h9BF: dout  = 8'b11111111; // 2495 : 255 - 0xff
      12'h9C0: dout  = 8'b11100001; // 2496 : 225 - 0xe1 -- Background 0x9c
      12'h9C1: dout  = 8'b11111001; // 2497 : 249 - 0xf9
      12'h9C2: dout  = 8'b11111101; // 2498 : 253 - 0xfd
      12'h9C3: dout  = 8'b11111111; // 2499 : 255 - 0xff
      12'h9C4: dout  = 8'b11111110; // 2500 : 254 - 0xfe
      12'h9C5: dout  = 8'b11111110; // 2501 : 254 - 0xfe
      12'h9C6: dout  = 8'b11111111; // 2502 : 255 - 0xff
      12'h9C7: dout  = 8'b11111111; // 2503 : 255 - 0xff
      12'h9C8: dout  = 8'b11111111; // 2504 : 255 - 0xff -- plane 1
      12'h9C9: dout  = 8'b11111111; // 2505 : 255 - 0xff
      12'h9CA: dout  = 8'b11111111; // 2506 : 255 - 0xff
      12'h9CB: dout  = 8'b11111111; // 2507 : 255 - 0xff
      12'h9CC: dout  = 8'b11111111; // 2508 : 255 - 0xff
      12'h9CD: dout  = 8'b11111111; // 2509 : 255 - 0xff
      12'h9CE: dout  = 8'b11111111; // 2510 : 255 - 0xff
      12'h9CF: dout  = 8'b11111111; // 2511 : 255 - 0xff
      12'h9D0: dout  = 8'b11110000; // 2512 : 240 - 0xf0 -- Background 0x9d
      12'h9D1: dout  = 8'b00010000; // 2513 :  16 - 0x10
      12'h9D2: dout  = 8'b00010000; // 2514 :  16 - 0x10
      12'h9D3: dout  = 8'b00010000; // 2515 :  16 - 0x10
      12'h9D4: dout  = 8'b00010000; // 2516 :  16 - 0x10
      12'h9D5: dout  = 8'b00010000; // 2517 :  16 - 0x10
      12'h9D6: dout  = 8'b00010000; // 2518 :  16 - 0x10
      12'h9D7: dout  = 8'b11111111; // 2519 : 255 - 0xff
      12'h9D8: dout  = 8'b00000000; // 2520 :   0 - 0x0 -- plane 1
      12'h9D9: dout  = 8'b11100000; // 2521 : 224 - 0xe0
      12'h9DA: dout  = 8'b11100000; // 2522 : 224 - 0xe0
      12'h9DB: dout  = 8'b11100000; // 2523 : 224 - 0xe0
      12'h9DC: dout  = 8'b11100000; // 2524 : 224 - 0xe0
      12'h9DD: dout  = 8'b11100000; // 2525 : 224 - 0xe0
      12'h9DE: dout  = 8'b11100000; // 2526 : 224 - 0xe0
      12'h9DF: dout  = 8'b11100000; // 2527 : 224 - 0xe0
      12'h9E0: dout  = 8'b00011111; // 2528 :  31 - 0x1f -- Background 0x9e
      12'h9E1: dout  = 8'b00010000; // 2529 :  16 - 0x10
      12'h9E2: dout  = 8'b00010000; // 2530 :  16 - 0x10
      12'h9E3: dout  = 8'b00010000; // 2531 :  16 - 0x10
      12'h9E4: dout  = 8'b00010000; // 2532 :  16 - 0x10
      12'h9E5: dout  = 8'b00010000; // 2533 :  16 - 0x10
      12'h9E6: dout  = 8'b00010000; // 2534 :  16 - 0x10
      12'h9E7: dout  = 8'b11111111; // 2535 : 255 - 0xff
      12'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout  = 8'b00001111; // 2537 :  15 - 0xf
      12'h9EA: dout  = 8'b00001111; // 2538 :  15 - 0xf
      12'h9EB: dout  = 8'b00001111; // 2539 :  15 - 0xf
      12'h9EC: dout  = 8'b00001111; // 2540 :  15 - 0xf
      12'h9ED: dout  = 8'b00001111; // 2541 :  15 - 0xf
      12'h9EE: dout  = 8'b00001111; // 2542 :  15 - 0xf
      12'h9EF: dout  = 8'b00001111; // 2543 :  15 - 0xf
      12'h9F0: dout  = 8'b10010010; // 2544 : 146 - 0x92 -- Background 0x9f
      12'h9F1: dout  = 8'b10010010; // 2545 : 146 - 0x92
      12'h9F2: dout  = 8'b10010010; // 2546 : 146 - 0x92
      12'h9F3: dout  = 8'b11111110; // 2547 : 254 - 0xfe
      12'h9F4: dout  = 8'b11111110; // 2548 : 254 - 0xfe
      12'h9F5: dout  = 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout  = 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout  = 8'b01001000; // 2552 :  72 - 0x48 -- plane 1
      12'h9F9: dout  = 8'b01001000; // 2553 :  72 - 0x48
      12'h9FA: dout  = 8'b01101100; // 2554 : 108 - 0x6c
      12'h9FB: dout  = 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout  = 8'b11111110; // 2558 : 254 - 0xfe
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00001010; // 2560 :  10 - 0xa -- Background 0xa0
      12'hA01: dout  = 8'b00001010; // 2561 :  10 - 0xa
      12'hA02: dout  = 8'b00111010; // 2562 :  58 - 0x3a
      12'hA03: dout  = 8'b00001010; // 2563 :  10 - 0xa
      12'hA04: dout  = 8'b11111011; // 2564 : 251 - 0xfb
      12'hA05: dout  = 8'b00001011; // 2565 :  11 - 0xb
      12'hA06: dout  = 8'b00001011; // 2566 :  11 - 0xb
      12'hA07: dout  = 8'b00001011; // 2567 :  11 - 0xb
      12'hA08: dout  = 8'b00000101; // 2568 :   5 - 0x5 -- plane 1
      12'hA09: dout  = 8'b00000101; // 2569 :   5 - 0x5
      12'hA0A: dout  = 8'b11000101; // 2570 : 197 - 0xc5
      12'hA0B: dout  = 8'b11110101; // 2571 : 245 - 0xf5
      12'hA0C: dout  = 8'b11110100; // 2572 : 244 - 0xf4
      12'hA0D: dout  = 8'b00000100; // 2573 :   4 - 0x4
      12'hA0E: dout  = 8'b00000100; // 2574 :   4 - 0x4
      12'hA0F: dout  = 8'b00000100; // 2575 :   4 - 0x4
      12'hA10: dout  = 8'b10010000; // 2576 : 144 - 0x90 -- Background 0xa1
      12'hA11: dout  = 8'b10010000; // 2577 : 144 - 0x90
      12'hA12: dout  = 8'b10011111; // 2578 : 159 - 0x9f
      12'hA13: dout  = 8'b10010000; // 2579 : 144 - 0x90
      12'hA14: dout  = 8'b10011111; // 2580 : 159 - 0x9f
      12'hA15: dout  = 8'b10010000; // 2581 : 144 - 0x90
      12'hA16: dout  = 8'b10010000; // 2582 : 144 - 0x90
      12'hA17: dout  = 8'b10010000; // 2583 : 144 - 0x90
      12'hA18: dout  = 8'b01110000; // 2584 : 112 - 0x70 -- plane 1
      12'hA19: dout  = 8'b01110000; // 2585 : 112 - 0x70
      12'hA1A: dout  = 8'b01110000; // 2586 : 112 - 0x70
      12'hA1B: dout  = 8'b01111111; // 2587 : 127 - 0x7f
      12'hA1C: dout  = 8'b01111111; // 2588 : 127 - 0x7f
      12'hA1D: dout  = 8'b01110000; // 2589 : 112 - 0x70
      12'hA1E: dout  = 8'b01110000; // 2590 : 112 - 0x70
      12'hA1F: dout  = 8'b01110000; // 2591 : 112 - 0x70
      12'hA20: dout  = 8'b00000001; // 2592 :   1 - 0x1 -- Background 0xa2
      12'hA21: dout  = 8'b00000001; // 2593 :   1 - 0x1
      12'hA22: dout  = 8'b00000001; // 2594 :   1 - 0x1
      12'hA23: dout  = 8'b00000001; // 2595 :   1 - 0x1
      12'hA24: dout  = 8'b00000001; // 2596 :   1 - 0x1
      12'hA25: dout  = 8'b00000001; // 2597 :   1 - 0x1
      12'hA26: dout  = 8'b00000001; // 2598 :   1 - 0x1
      12'hA27: dout  = 8'b00000001; // 2599 :   1 - 0x1
      12'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout  = 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout  = 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout  = 8'b10000000; // 2608 : 128 - 0x80 -- Background 0xa3
      12'hA31: dout  = 8'b10000000; // 2609 : 128 - 0x80
      12'hA32: dout  = 8'b10000000; // 2610 : 128 - 0x80
      12'hA33: dout  = 8'b10000000; // 2611 : 128 - 0x80
      12'hA34: dout  = 8'b10000000; // 2612 : 128 - 0x80
      12'hA35: dout  = 8'b10000000; // 2613 : 128 - 0x80
      12'hA36: dout  = 8'b10000000; // 2614 : 128 - 0x80
      12'hA37: dout  = 8'b10000000; // 2615 : 128 - 0x80
      12'hA38: dout  = 8'b00000000; // 2616 :   0 - 0x0 -- plane 1
      12'hA39: dout  = 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout  = 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout  = 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout  = 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout  = 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout  = 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b00001000; // 2624 :   8 - 0x8 -- Background 0xa4
      12'hA41: dout  = 8'b10001000; // 2625 : 136 - 0x88
      12'hA42: dout  = 8'b10010001; // 2626 : 145 - 0x91
      12'hA43: dout  = 8'b11010001; // 2627 : 209 - 0xd1
      12'hA44: dout  = 8'b01010011; // 2628 :  83 - 0x53
      12'hA45: dout  = 8'b01010011; // 2629 :  83 - 0x53
      12'hA46: dout  = 8'b01110011; // 2630 : 115 - 0x73
      12'hA47: dout  = 8'b00111111; // 2631 :  63 - 0x3f
      12'hA48: dout  = 8'b11111111; // 2632 : 255 - 0xff -- plane 1
      12'hA49: dout  = 8'b11111111; // 2633 : 255 - 0xff
      12'hA4A: dout  = 8'b11111111; // 2634 : 255 - 0xff
      12'hA4B: dout  = 8'b11111111; // 2635 : 255 - 0xff
      12'hA4C: dout  = 8'b11111111; // 2636 : 255 - 0xff
      12'hA4D: dout  = 8'b11111110; // 2637 : 254 - 0xfe
      12'hA4E: dout  = 8'b10111110; // 2638 : 190 - 0xbe
      12'hA4F: dout  = 8'b11001110; // 2639 : 206 - 0xce
      12'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Background 0xa5
      12'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout  = 8'b00000111; // 2642 :   7 - 0x7
      12'hA53: dout  = 8'b00001111; // 2643 :  15 - 0xf
      12'hA54: dout  = 8'b00001100; // 2644 :  12 - 0xc
      12'hA55: dout  = 8'b00011011; // 2645 :  27 - 0x1b
      12'hA56: dout  = 8'b00011011; // 2646 :  27 - 0x1b
      12'hA57: dout  = 8'b00011011; // 2647 :  27 - 0x1b
      12'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout  = 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout  = 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout  = 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout  = 8'b00000011; // 2652 :   3 - 0x3
      12'hA5D: dout  = 8'b00000100; // 2653 :   4 - 0x4
      12'hA5E: dout  = 8'b00000100; // 2654 :   4 - 0x4
      12'hA5F: dout  = 8'b00000100; // 2655 :   4 - 0x4
      12'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Background 0xa6
      12'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout  = 8'b11100000; // 2658 : 224 - 0xe0
      12'hA63: dout  = 8'b11110000; // 2659 : 240 - 0xf0
      12'hA64: dout  = 8'b11110000; // 2660 : 240 - 0xf0
      12'hA65: dout  = 8'b11111000; // 2661 : 248 - 0xf8
      12'hA66: dout  = 8'b11111000; // 2662 : 248 - 0xf8
      12'hA67: dout  = 8'b11111000; // 2663 : 248 - 0xf8
      12'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b01100000; // 2666 :  96 - 0x60
      12'hA6B: dout  = 8'b00110000; // 2667 :  48 - 0x30
      12'hA6C: dout  = 8'b00110000; // 2668 :  48 - 0x30
      12'hA6D: dout  = 8'b10011000; // 2669 : 152 - 0x98
      12'hA6E: dout  = 8'b10011000; // 2670 : 152 - 0x98
      12'hA6F: dout  = 8'b10011000; // 2671 : 152 - 0x98
      12'hA70: dout  = 8'b00011011; // 2672 :  27 - 0x1b -- Background 0xa7
      12'hA71: dout  = 8'b00011011; // 2673 :  27 - 0x1b
      12'hA72: dout  = 8'b00011011; // 2674 :  27 - 0x1b
      12'hA73: dout  = 8'b00011011; // 2675 :  27 - 0x1b
      12'hA74: dout  = 8'b00011011; // 2676 :  27 - 0x1b
      12'hA75: dout  = 8'b00001111; // 2677 :  15 - 0xf
      12'hA76: dout  = 8'b00001111; // 2678 :  15 - 0xf
      12'hA77: dout  = 8'b00000111; // 2679 :   7 - 0x7
      12'hA78: dout  = 8'b00000100; // 2680 :   4 - 0x4 -- plane 1
      12'hA79: dout  = 8'b00000100; // 2681 :   4 - 0x4
      12'hA7A: dout  = 8'b00000100; // 2682 :   4 - 0x4
      12'hA7B: dout  = 8'b00000100; // 2683 :   4 - 0x4
      12'hA7C: dout  = 8'b00000100; // 2684 :   4 - 0x4
      12'hA7D: dout  = 8'b00000011; // 2685 :   3 - 0x3
      12'hA7E: dout  = 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout  = 8'b11111000; // 2688 : 248 - 0xf8 -- Background 0xa8
      12'hA81: dout  = 8'b11111000; // 2689 : 248 - 0xf8
      12'hA82: dout  = 8'b11111000; // 2690 : 248 - 0xf8
      12'hA83: dout  = 8'b11111000; // 2691 : 248 - 0xf8
      12'hA84: dout  = 8'b11111000; // 2692 : 248 - 0xf8
      12'hA85: dout  = 8'b11110000; // 2693 : 240 - 0xf0
      12'hA86: dout  = 8'b11110000; // 2694 : 240 - 0xf0
      12'hA87: dout  = 8'b11100000; // 2695 : 224 - 0xe0
      12'hA88: dout  = 8'b10011000; // 2696 : 152 - 0x98 -- plane 1
      12'hA89: dout  = 8'b10011000; // 2697 : 152 - 0x98
      12'hA8A: dout  = 8'b10011000; // 2698 : 152 - 0x98
      12'hA8B: dout  = 8'b10011000; // 2699 : 152 - 0x98
      12'hA8C: dout  = 8'b10011000; // 2700 : 152 - 0x98
      12'hA8D: dout  = 8'b00110000; // 2701 :  48 - 0x30
      12'hA8E: dout  = 8'b00110000; // 2702 :  48 - 0x30
      12'hA8F: dout  = 8'b01100000; // 2703 :  96 - 0x60
      12'hA90: dout  = 8'b11110001; // 2704 : 241 - 0xf1 -- Background 0xa9
      12'hA91: dout  = 8'b00010001; // 2705 :  17 - 0x11
      12'hA92: dout  = 8'b00010001; // 2706 :  17 - 0x11
      12'hA93: dout  = 8'b00011111; // 2707 :  31 - 0x1f
      12'hA94: dout  = 8'b00010000; // 2708 :  16 - 0x10
      12'hA95: dout  = 8'b00010000; // 2709 :  16 - 0x10
      12'hA96: dout  = 8'b00010000; // 2710 :  16 - 0x10
      12'hA97: dout  = 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout  = 8'b00001111; // 2712 :  15 - 0xf -- plane 1
      12'hA99: dout  = 8'b11101111; // 2713 : 239 - 0xef
      12'hA9A: dout  = 8'b11101111; // 2714 : 239 - 0xef
      12'hA9B: dout  = 8'b11101111; // 2715 : 239 - 0xef
      12'hA9C: dout  = 8'b11101111; // 2716 : 239 - 0xef
      12'hA9D: dout  = 8'b11101111; // 2717 : 239 - 0xef
      12'hA9E: dout  = 8'b11101111; // 2718 : 239 - 0xef
      12'hA9F: dout  = 8'b11100000; // 2719 : 224 - 0xe0
      12'hAA0: dout  = 8'b00011111; // 2720 :  31 - 0x1f -- Background 0xaa
      12'hAA1: dout  = 8'b00010000; // 2721 :  16 - 0x10
      12'hAA2: dout  = 8'b00010000; // 2722 :  16 - 0x10
      12'hAA3: dout  = 8'b11110000; // 2723 : 240 - 0xf0
      12'hAA4: dout  = 8'b00010000; // 2724 :  16 - 0x10
      12'hAA5: dout  = 8'b00010000; // 2725 :  16 - 0x10
      12'hAA6: dout  = 8'b00010000; // 2726 :  16 - 0x10
      12'hAA7: dout  = 8'b11111111; // 2727 : 255 - 0xff
      12'hAA8: dout  = 8'b11100000; // 2728 : 224 - 0xe0 -- plane 1
      12'hAA9: dout  = 8'b11101111; // 2729 : 239 - 0xef
      12'hAAA: dout  = 8'b11101111; // 2730 : 239 - 0xef
      12'hAAB: dout  = 8'b11101111; // 2731 : 239 - 0xef
      12'hAAC: dout  = 8'b11101111; // 2732 : 239 - 0xef
      12'hAAD: dout  = 8'b11101111; // 2733 : 239 - 0xef
      12'hAAE: dout  = 8'b11101111; // 2734 : 239 - 0xef
      12'hAAF: dout  = 8'b00001111; // 2735 :  15 - 0xf
      12'hAB0: dout  = 8'b01111111; // 2736 : 127 - 0x7f -- Background 0xab
      12'hAB1: dout  = 8'b10111111; // 2737 : 191 - 0xbf
      12'hAB2: dout  = 8'b11011111; // 2738 : 223 - 0xdf
      12'hAB3: dout  = 8'b11101111; // 2739 : 239 - 0xef
      12'hAB4: dout  = 8'b11110000; // 2740 : 240 - 0xf0
      12'hAB5: dout  = 8'b11110000; // 2741 : 240 - 0xf0
      12'hAB6: dout  = 8'b11110000; // 2742 : 240 - 0xf0
      12'hAB7: dout  = 8'b11110000; // 2743 : 240 - 0xf0
      12'hAB8: dout  = 8'b10000000; // 2744 : 128 - 0x80 -- plane 1
      12'hAB9: dout  = 8'b01000000; // 2745 :  64 - 0x40
      12'hABA: dout  = 8'b00100000; // 2746 :  32 - 0x20
      12'hABB: dout  = 8'b00010000; // 2747 :  16 - 0x10
      12'hABC: dout  = 8'b00001111; // 2748 :  15 - 0xf
      12'hABD: dout  = 8'b00001111; // 2749 :  15 - 0xf
      12'hABE: dout  = 8'b00001111; // 2750 :  15 - 0xf
      12'hABF: dout  = 8'b00001111; // 2751 :  15 - 0xf
      12'hAC0: dout  = 8'b11110000; // 2752 : 240 - 0xf0 -- Background 0xac
      12'hAC1: dout  = 8'b11110000; // 2753 : 240 - 0xf0
      12'hAC2: dout  = 8'b11110000; // 2754 : 240 - 0xf0
      12'hAC3: dout  = 8'b11110000; // 2755 : 240 - 0xf0
      12'hAC4: dout  = 8'b11111111; // 2756 : 255 - 0xff
      12'hAC5: dout  = 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout  = 8'b11111111; // 2758 : 255 - 0xff
      12'hAC7: dout  = 8'b11111111; // 2759 : 255 - 0xff
      12'hAC8: dout  = 8'b00001111; // 2760 :  15 - 0xf -- plane 1
      12'hAC9: dout  = 8'b00001111; // 2761 :  15 - 0xf
      12'hACA: dout  = 8'b00001111; // 2762 :  15 - 0xf
      12'hACB: dout  = 8'b00001111; // 2763 :  15 - 0xf
      12'hACC: dout  = 8'b00011111; // 2764 :  31 - 0x1f
      12'hACD: dout  = 8'b00111111; // 2765 :  63 - 0x3f
      12'hACE: dout  = 8'b01111111; // 2766 : 127 - 0x7f
      12'hACF: dout  = 8'b11111111; // 2767 : 255 - 0xff
      12'hAD0: dout  = 8'b11111111; // 2768 : 255 - 0xff -- Background 0xad
      12'hAD1: dout  = 8'b11111111; // 2769 : 255 - 0xff
      12'hAD2: dout  = 8'b11111111; // 2770 : 255 - 0xff
      12'hAD3: dout  = 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout  = 8'b00001111; // 2772 :  15 - 0xf
      12'hAD5: dout  = 8'b00001111; // 2773 :  15 - 0xf
      12'hAD6: dout  = 8'b00001111; // 2774 :  15 - 0xf
      12'hAD7: dout  = 8'b00001111; // 2775 :  15 - 0xf
      12'hAD8: dout  = 8'b00000001; // 2776 :   1 - 0x1 -- plane 1
      12'hAD9: dout  = 8'b00000011; // 2777 :   3 - 0x3
      12'hADA: dout  = 8'b00000111; // 2778 :   7 - 0x7
      12'hADB: dout  = 8'b00001111; // 2779 :  15 - 0xf
      12'hADC: dout  = 8'b11111111; // 2780 : 255 - 0xff
      12'hADD: dout  = 8'b11111111; // 2781 : 255 - 0xff
      12'hADE: dout  = 8'b11111111; // 2782 : 255 - 0xff
      12'hADF: dout  = 8'b11111111; // 2783 : 255 - 0xff
      12'hAE0: dout  = 8'b00001111; // 2784 :  15 - 0xf -- Background 0xae
      12'hAE1: dout  = 8'b00001111; // 2785 :  15 - 0xf
      12'hAE2: dout  = 8'b00001111; // 2786 :  15 - 0xf
      12'hAE3: dout  = 8'b00001111; // 2787 :  15 - 0xf
      12'hAE4: dout  = 8'b11110111; // 2788 : 247 - 0xf7
      12'hAE5: dout  = 8'b11111011; // 2789 : 251 - 0xfb
      12'hAE6: dout  = 8'b11111101; // 2790 : 253 - 0xfd
      12'hAE7: dout  = 8'b11111110; // 2791 : 254 - 0xfe
      12'hAE8: dout  = 8'b11111111; // 2792 : 255 - 0xff -- plane 1
      12'hAE9: dout  = 8'b11111111; // 2793 : 255 - 0xff
      12'hAEA: dout  = 8'b11111111; // 2794 : 255 - 0xff
      12'hAEB: dout  = 8'b11111111; // 2795 : 255 - 0xff
      12'hAEC: dout  = 8'b11111111; // 2796 : 255 - 0xff
      12'hAED: dout  = 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout  = 8'b11111111; // 2798 : 255 - 0xff
      12'hAEF: dout  = 8'b11111111; // 2799 : 255 - 0xff
      12'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Background 0xaf
      12'hAF1: dout  = 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout  = 8'b00000000; // 2802 :   0 - 0x0
      12'hAF3: dout  = 8'b00000000; // 2803 :   0 - 0x0
      12'hAF4: dout  = 8'b00000000; // 2804 :   0 - 0x0
      12'hAF5: dout  = 8'b00000000; // 2805 :   0 - 0x0
      12'hAF6: dout  = 8'b00011000; // 2806 :  24 - 0x18
      12'hAF7: dout  = 8'b00011000; // 2807 :  24 - 0x18
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout  = 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout  = 8'b00011111; // 2816 :  31 - 0x1f -- Background 0xb0
      12'hB01: dout  = 8'b00111111; // 2817 :  63 - 0x3f
      12'hB02: dout  = 8'b01111111; // 2818 : 127 - 0x7f
      12'hB03: dout  = 8'b01111111; // 2819 : 127 - 0x7f
      12'hB04: dout  = 8'b01111111; // 2820 : 127 - 0x7f
      12'hB05: dout  = 8'b11111111; // 2821 : 255 - 0xff
      12'hB06: dout  = 8'b11111111; // 2822 : 255 - 0xff
      12'hB07: dout  = 8'b11111111; // 2823 : 255 - 0xff
      12'hB08: dout  = 8'b00011111; // 2824 :  31 - 0x1f -- plane 1
      12'hB09: dout  = 8'b00100000; // 2825 :  32 - 0x20
      12'hB0A: dout  = 8'b01000000; // 2826 :  64 - 0x40
      12'hB0B: dout  = 8'b01000000; // 2827 :  64 - 0x40
      12'hB0C: dout  = 8'b01000000; // 2828 :  64 - 0x40
      12'hB0D: dout  = 8'b10000000; // 2829 : 128 - 0x80
      12'hB0E: dout  = 8'b10000010; // 2830 : 130 - 0x82
      12'hB0F: dout  = 8'b10000010; // 2831 : 130 - 0x82
      12'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Background 0xb1
      12'hB11: dout  = 8'b11111111; // 2833 : 255 - 0xff
      12'hB12: dout  = 8'b11111111; // 2834 : 255 - 0xff
      12'hB13: dout  = 8'b01111111; // 2835 : 127 - 0x7f
      12'hB14: dout  = 8'b01111111; // 2836 : 127 - 0x7f
      12'hB15: dout  = 8'b01111111; // 2837 : 127 - 0x7f
      12'hB16: dout  = 8'b00111111; // 2838 :  63 - 0x3f
      12'hB17: dout  = 8'b00011110; // 2839 :  30 - 0x1e
      12'hB18: dout  = 8'b10000010; // 2840 : 130 - 0x82 -- plane 1
      12'hB19: dout  = 8'b10000000; // 2841 : 128 - 0x80
      12'hB1A: dout  = 8'b10100000; // 2842 : 160 - 0xa0
      12'hB1B: dout  = 8'b01000100; // 2843 :  68 - 0x44
      12'hB1C: dout  = 8'b01000011; // 2844 :  67 - 0x43
      12'hB1D: dout  = 8'b01000000; // 2845 :  64 - 0x40
      12'hB1E: dout  = 8'b00100001; // 2846 :  33 - 0x21
      12'hB1F: dout  = 8'b00011110; // 2847 :  30 - 0x1e
      12'hB20: dout  = 8'b11111000; // 2848 : 248 - 0xf8 -- Background 0xb2
      12'hB21: dout  = 8'b11111100; // 2849 : 252 - 0xfc
      12'hB22: dout  = 8'b11111110; // 2850 : 254 - 0xfe
      12'hB23: dout  = 8'b11111110; // 2851 : 254 - 0xfe
      12'hB24: dout  = 8'b11111110; // 2852 : 254 - 0xfe
      12'hB25: dout  = 8'b11111111; // 2853 : 255 - 0xff
      12'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      12'hB27: dout  = 8'b11111111; // 2855 : 255 - 0xff
      12'hB28: dout  = 8'b11111000; // 2856 : 248 - 0xf8 -- plane 1
      12'hB29: dout  = 8'b00000100; // 2857 :   4 - 0x4
      12'hB2A: dout  = 8'b00000010; // 2858 :   2 - 0x2
      12'hB2B: dout  = 8'b00000010; // 2859 :   2 - 0x2
      12'hB2C: dout  = 8'b00000010; // 2860 :   2 - 0x2
      12'hB2D: dout  = 8'b00000001; // 2861 :   1 - 0x1
      12'hB2E: dout  = 8'b01000001; // 2862 :  65 - 0x41
      12'hB2F: dout  = 8'b01000001; // 2863 :  65 - 0x41
      12'hB30: dout  = 8'b11111111; // 2864 : 255 - 0xff -- Background 0xb3
      12'hB31: dout  = 8'b11111111; // 2865 : 255 - 0xff
      12'hB32: dout  = 8'b11111111; // 2866 : 255 - 0xff
      12'hB33: dout  = 8'b11111110; // 2867 : 254 - 0xfe
      12'hB34: dout  = 8'b11111110; // 2868 : 254 - 0xfe
      12'hB35: dout  = 8'b11111110; // 2869 : 254 - 0xfe
      12'hB36: dout  = 8'b11111100; // 2870 : 252 - 0xfc
      12'hB37: dout  = 8'b01111000; // 2871 : 120 - 0x78
      12'hB38: dout  = 8'b01000001; // 2872 :  65 - 0x41 -- plane 1
      12'hB39: dout  = 8'b00000001; // 2873 :   1 - 0x1
      12'hB3A: dout  = 8'b00000101; // 2874 :   5 - 0x5
      12'hB3B: dout  = 8'b00100010; // 2875 :  34 - 0x22
      12'hB3C: dout  = 8'b11000010; // 2876 : 194 - 0xc2
      12'hB3D: dout  = 8'b00000010; // 2877 :   2 - 0x2
      12'hB3E: dout  = 8'b10000100; // 2878 : 132 - 0x84
      12'hB3F: dout  = 8'b01111000; // 2879 : 120 - 0x78
      12'hB40: dout  = 8'b01111111; // 2880 : 127 - 0x7f -- Background 0xb4
      12'hB41: dout  = 8'b10000000; // 2881 : 128 - 0x80
      12'hB42: dout  = 8'b10000000; // 2882 : 128 - 0x80
      12'hB43: dout  = 8'b10000000; // 2883 : 128 - 0x80
      12'hB44: dout  = 8'b10000000; // 2884 : 128 - 0x80
      12'hB45: dout  = 8'b10000000; // 2885 : 128 - 0x80
      12'hB46: dout  = 8'b10000000; // 2886 : 128 - 0x80
      12'hB47: dout  = 8'b10000000; // 2887 : 128 - 0x80
      12'hB48: dout  = 8'b10000000; // 2888 : 128 - 0x80 -- plane 1
      12'hB49: dout  = 8'b01111111; // 2889 : 127 - 0x7f
      12'hB4A: dout  = 8'b01111111; // 2890 : 127 - 0x7f
      12'hB4B: dout  = 8'b01111111; // 2891 : 127 - 0x7f
      12'hB4C: dout  = 8'b01111111; // 2892 : 127 - 0x7f
      12'hB4D: dout  = 8'b01111111; // 2893 : 127 - 0x7f
      12'hB4E: dout  = 8'b01111111; // 2894 : 127 - 0x7f
      12'hB4F: dout  = 8'b01111111; // 2895 : 127 - 0x7f
      12'hB50: dout  = 8'b11011110; // 2896 : 222 - 0xde -- Background 0xb5
      12'hB51: dout  = 8'b01100001; // 2897 :  97 - 0x61
      12'hB52: dout  = 8'b01100001; // 2898 :  97 - 0x61
      12'hB53: dout  = 8'b01100001; // 2899 :  97 - 0x61
      12'hB54: dout  = 8'b01110001; // 2900 : 113 - 0x71
      12'hB55: dout  = 8'b01011110; // 2901 :  94 - 0x5e
      12'hB56: dout  = 8'b01111111; // 2902 : 127 - 0x7f
      12'hB57: dout  = 8'b01100001; // 2903 :  97 - 0x61
      12'hB58: dout  = 8'b01100001; // 2904 :  97 - 0x61 -- plane 1
      12'hB59: dout  = 8'b11011111; // 2905 : 223 - 0xdf
      12'hB5A: dout  = 8'b11011111; // 2906 : 223 - 0xdf
      12'hB5B: dout  = 8'b11011111; // 2907 : 223 - 0xdf
      12'hB5C: dout  = 8'b11011111; // 2908 : 223 - 0xdf
      12'hB5D: dout  = 8'b11111111; // 2909 : 255 - 0xff
      12'hB5E: dout  = 8'b11000001; // 2910 : 193 - 0xc1
      12'hB5F: dout  = 8'b11011111; // 2911 : 223 - 0xdf
      12'hB60: dout  = 8'b10000000; // 2912 : 128 - 0x80 -- Background 0xb6
      12'hB61: dout  = 8'b10000000; // 2913 : 128 - 0x80
      12'hB62: dout  = 8'b11000000; // 2914 : 192 - 0xc0
      12'hB63: dout  = 8'b11110000; // 2915 : 240 - 0xf0
      12'hB64: dout  = 8'b10111111; // 2916 : 191 - 0xbf
      12'hB65: dout  = 8'b10001111; // 2917 : 143 - 0x8f
      12'hB66: dout  = 8'b10000001; // 2918 : 129 - 0x81
      12'hB67: dout  = 8'b01111110; // 2919 : 126 - 0x7e
      12'hB68: dout  = 8'b01111111; // 2920 : 127 - 0x7f -- plane 1
      12'hB69: dout  = 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout  = 8'b11111111; // 2922 : 255 - 0xff
      12'hB6B: dout  = 8'b00111111; // 2923 :  63 - 0x3f
      12'hB6C: dout  = 8'b01001111; // 2924 :  79 - 0x4f
      12'hB6D: dout  = 8'b01110001; // 2925 : 113 - 0x71
      12'hB6E: dout  = 8'b01111111; // 2926 : 127 - 0x7f
      12'hB6F: dout  = 8'b11111111; // 2927 : 255 - 0xff
      12'hB70: dout  = 8'b01100001; // 2928 :  97 - 0x61 -- Background 0xb7
      12'hB71: dout  = 8'b01100001; // 2929 :  97 - 0x61
      12'hB72: dout  = 8'b11000001; // 2930 : 193 - 0xc1
      12'hB73: dout  = 8'b11000001; // 2931 : 193 - 0xc1
      12'hB74: dout  = 8'b10000001; // 2932 : 129 - 0x81
      12'hB75: dout  = 8'b10000001; // 2933 : 129 - 0x81
      12'hB76: dout  = 8'b10000011; // 2934 : 131 - 0x83
      12'hB77: dout  = 8'b11111110; // 2935 : 254 - 0xfe
      12'hB78: dout  = 8'b11011111; // 2936 : 223 - 0xdf -- plane 1
      12'hB79: dout  = 8'b11011111; // 2937 : 223 - 0xdf
      12'hB7A: dout  = 8'b10111111; // 2938 : 191 - 0xbf
      12'hB7B: dout  = 8'b10111111; // 2939 : 191 - 0xbf
      12'hB7C: dout  = 8'b01111111; // 2940 : 127 - 0x7f
      12'hB7D: dout  = 8'b01111111; // 2941 : 127 - 0x7f
      12'hB7E: dout  = 8'b01111111; // 2942 : 127 - 0x7f
      12'hB7F: dout  = 8'b01111111; // 2943 : 127 - 0x7f
      12'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Background 0xb8
      12'hB81: dout  = 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout  = 8'b00000011; // 2946 :   3 - 0x3
      12'hB83: dout  = 8'b00001111; // 2947 :  15 - 0xf
      12'hB84: dout  = 8'b00011111; // 2948 :  31 - 0x1f
      12'hB85: dout  = 8'b00111111; // 2949 :  63 - 0x3f
      12'hB86: dout  = 8'b01111111; // 2950 : 127 - 0x7f
      12'hB87: dout  = 8'b01111111; // 2951 : 127 - 0x7f
      12'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout  = 8'b00000011; // 2954 :   3 - 0x3
      12'hB8B: dout  = 8'b00001100; // 2955 :  12 - 0xc
      12'hB8C: dout  = 8'b00010000; // 2956 :  16 - 0x10
      12'hB8D: dout  = 8'b00100000; // 2957 :  32 - 0x20
      12'hB8E: dout  = 8'b01000000; // 2958 :  64 - 0x40
      12'hB8F: dout  = 8'b01000000; // 2959 :  64 - 0x40
      12'hB90: dout  = 8'b00000000; // 2960 :   0 - 0x0 -- Background 0xb9
      12'hB91: dout  = 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout  = 8'b11000000; // 2962 : 192 - 0xc0
      12'hB93: dout  = 8'b11110000; // 2963 : 240 - 0xf0
      12'hB94: dout  = 8'b11111000; // 2964 : 248 - 0xf8
      12'hB95: dout  = 8'b11111100; // 2965 : 252 - 0xfc
      12'hB96: dout  = 8'b11111110; // 2966 : 254 - 0xfe
      12'hB97: dout  = 8'b11111110; // 2967 : 254 - 0xfe
      12'hB98: dout  = 8'b00000000; // 2968 :   0 - 0x0 -- plane 1
      12'hB99: dout  = 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout  = 8'b11000000; // 2970 : 192 - 0xc0
      12'hB9B: dout  = 8'b00110000; // 2971 :  48 - 0x30
      12'hB9C: dout  = 8'b00001000; // 2972 :   8 - 0x8
      12'hB9D: dout  = 8'b00000100; // 2973 :   4 - 0x4
      12'hB9E: dout  = 8'b00000010; // 2974 :   2 - 0x2
      12'hB9F: dout  = 8'b00000010; // 2975 :   2 - 0x2
      12'hBA0: dout  = 8'b11111111; // 2976 : 255 - 0xff -- Background 0xba
      12'hBA1: dout  = 8'b11111111; // 2977 : 255 - 0xff
      12'hBA2: dout  = 8'b11111111; // 2978 : 255 - 0xff
      12'hBA3: dout  = 8'b11111111; // 2979 : 255 - 0xff
      12'hBA4: dout  = 8'b11111111; // 2980 : 255 - 0xff
      12'hBA5: dout  = 8'b11111111; // 2981 : 255 - 0xff
      12'hBA6: dout  = 8'b11111111; // 2982 : 255 - 0xff
      12'hBA7: dout  = 8'b11111111; // 2983 : 255 - 0xff
      12'hBA8: dout  = 8'b10000000; // 2984 : 128 - 0x80 -- plane 1
      12'hBA9: dout  = 8'b10000000; // 2985 : 128 - 0x80
      12'hBAA: dout  = 8'b10000000; // 2986 : 128 - 0x80
      12'hBAB: dout  = 8'b10000000; // 2987 : 128 - 0x80
      12'hBAC: dout  = 8'b10000000; // 2988 : 128 - 0x80
      12'hBAD: dout  = 8'b10000000; // 2989 : 128 - 0x80
      12'hBAE: dout  = 8'b10000000; // 2990 : 128 - 0x80
      12'hBAF: dout  = 8'b10000000; // 2991 : 128 - 0x80
      12'hBB0: dout  = 8'b11111111; // 2992 : 255 - 0xff -- Background 0xbb
      12'hBB1: dout  = 8'b11111111; // 2993 : 255 - 0xff
      12'hBB2: dout  = 8'b11111111; // 2994 : 255 - 0xff
      12'hBB3: dout  = 8'b11111111; // 2995 : 255 - 0xff
      12'hBB4: dout  = 8'b11111111; // 2996 : 255 - 0xff
      12'hBB5: dout  = 8'b11111111; // 2997 : 255 - 0xff
      12'hBB6: dout  = 8'b11111111; // 2998 : 255 - 0xff
      12'hBB7: dout  = 8'b11111111; // 2999 : 255 - 0xff
      12'hBB8: dout  = 8'b00000001; // 3000 :   1 - 0x1 -- plane 1
      12'hBB9: dout  = 8'b00000001; // 3001 :   1 - 0x1
      12'hBBA: dout  = 8'b00000001; // 3002 :   1 - 0x1
      12'hBBB: dout  = 8'b00000001; // 3003 :   1 - 0x1
      12'hBBC: dout  = 8'b00000001; // 3004 :   1 - 0x1
      12'hBBD: dout  = 8'b00000001; // 3005 :   1 - 0x1
      12'hBBE: dout  = 8'b00000001; // 3006 :   1 - 0x1
      12'hBBF: dout  = 8'b00000001; // 3007 :   1 - 0x1
      12'hBC0: dout  = 8'b01111111; // 3008 : 127 - 0x7f -- Background 0xbc
      12'hBC1: dout  = 8'b01111111; // 3009 : 127 - 0x7f
      12'hBC2: dout  = 8'b01111111; // 3010 : 127 - 0x7f
      12'hBC3: dout  = 8'b00111111; // 3011 :  63 - 0x3f
      12'hBC4: dout  = 8'b00111111; // 3012 :  63 - 0x3f
      12'hBC5: dout  = 8'b00011111; // 3013 :  31 - 0x1f
      12'hBC6: dout  = 8'b00001111; // 3014 :  15 - 0xf
      12'hBC7: dout  = 8'b00000111; // 3015 :   7 - 0x7
      12'hBC8: dout  = 8'b01000000; // 3016 :  64 - 0x40 -- plane 1
      12'hBC9: dout  = 8'b01000000; // 3017 :  64 - 0x40
      12'hBCA: dout  = 8'b01000000; // 3018 :  64 - 0x40
      12'hBCB: dout  = 8'b00100000; // 3019 :  32 - 0x20
      12'hBCC: dout  = 8'b00110000; // 3020 :  48 - 0x30
      12'hBCD: dout  = 8'b00011100; // 3021 :  28 - 0x1c
      12'hBCE: dout  = 8'b00001111; // 3022 :  15 - 0xf
      12'hBCF: dout  = 8'b00000111; // 3023 :   7 - 0x7
      12'hBD0: dout  = 8'b11111110; // 3024 : 254 - 0xfe -- Background 0xbd
      12'hBD1: dout  = 8'b11111110; // 3025 : 254 - 0xfe
      12'hBD2: dout  = 8'b11111110; // 3026 : 254 - 0xfe
      12'hBD3: dout  = 8'b11111100; // 3027 : 252 - 0xfc
      12'hBD4: dout  = 8'b11111100; // 3028 : 252 - 0xfc
      12'hBD5: dout  = 8'b11111000; // 3029 : 248 - 0xf8
      12'hBD6: dout  = 8'b11110000; // 3030 : 240 - 0xf0
      12'hBD7: dout  = 8'b11110000; // 3031 : 240 - 0xf0
      12'hBD8: dout  = 8'b00000010; // 3032 :   2 - 0x2 -- plane 1
      12'hBD9: dout  = 8'b00000010; // 3033 :   2 - 0x2
      12'hBDA: dout  = 8'b00000010; // 3034 :   2 - 0x2
      12'hBDB: dout  = 8'b00000100; // 3035 :   4 - 0x4
      12'hBDC: dout  = 8'b00001100; // 3036 :  12 - 0xc
      12'hBDD: dout  = 8'b00111000; // 3037 :  56 - 0x38
      12'hBDE: dout  = 8'b11110000; // 3038 : 240 - 0xf0
      12'hBDF: dout  = 8'b11110000; // 3039 : 240 - 0xf0
      12'hBE0: dout  = 8'b00001111; // 3040 :  15 - 0xf -- Background 0xbe
      12'hBE1: dout  = 8'b00001111; // 3041 :  15 - 0xf
      12'hBE2: dout  = 8'b00001111; // 3042 :  15 - 0xf
      12'hBE3: dout  = 8'b00001111; // 3043 :  15 - 0xf
      12'hBE4: dout  = 8'b00001111; // 3044 :  15 - 0xf
      12'hBE5: dout  = 8'b00001111; // 3045 :  15 - 0xf
      12'hBE6: dout  = 8'b00000111; // 3046 :   7 - 0x7
      12'hBE7: dout  = 8'b00001111; // 3047 :  15 - 0xf
      12'hBE8: dout  = 8'b00001000; // 3048 :   8 - 0x8 -- plane 1
      12'hBE9: dout  = 8'b00001000; // 3049 :   8 - 0x8
      12'hBEA: dout  = 8'b00001000; // 3050 :   8 - 0x8
      12'hBEB: dout  = 8'b00001000; // 3051 :   8 - 0x8
      12'hBEC: dout  = 8'b00001000; // 3052 :   8 - 0x8
      12'hBED: dout  = 8'b00001100; // 3053 :  12 - 0xc
      12'hBEE: dout  = 8'b00000101; // 3054 :   5 - 0x5
      12'hBEF: dout  = 8'b00001010; // 3055 :  10 - 0xa
      12'hBF0: dout  = 8'b11110000; // 3056 : 240 - 0xf0 -- Background 0xbf
      12'hBF1: dout  = 8'b11110000; // 3057 : 240 - 0xf0
      12'hBF2: dout  = 8'b11110000; // 3058 : 240 - 0xf0
      12'hBF3: dout  = 8'b11110000; // 3059 : 240 - 0xf0
      12'hBF4: dout  = 8'b11110000; // 3060 : 240 - 0xf0
      12'hBF5: dout  = 8'b11110000; // 3061 : 240 - 0xf0
      12'hBF6: dout  = 8'b11100000; // 3062 : 224 - 0xe0
      12'hBF7: dout  = 8'b11110000; // 3063 : 240 - 0xf0
      12'hBF8: dout  = 8'b00010000; // 3064 :  16 - 0x10 -- plane 1
      12'hBF9: dout  = 8'b01010000; // 3065 :  80 - 0x50
      12'hBFA: dout  = 8'b01010000; // 3066 :  80 - 0x50
      12'hBFB: dout  = 8'b01010000; // 3067 :  80 - 0x50
      12'hBFC: dout  = 8'b01010000; // 3068 :  80 - 0x50
      12'hBFD: dout  = 8'b00110000; // 3069 :  48 - 0x30
      12'hBFE: dout  = 8'b10100000; // 3070 : 160 - 0xa0
      12'hBFF: dout  = 8'b01010000; // 3071 :  80 - 0x50
      12'hC00: dout  = 8'b10000001; // 3072 : 129 - 0x81 -- Background 0xc0
      12'hC01: dout  = 8'b11000001; // 3073 : 193 - 0xc1
      12'hC02: dout  = 8'b10100011; // 3074 : 163 - 0xa3
      12'hC03: dout  = 8'b10100011; // 3075 : 163 - 0xa3
      12'hC04: dout  = 8'b10011101; // 3076 : 157 - 0x9d
      12'hC05: dout  = 8'b10000001; // 3077 : 129 - 0x81
      12'hC06: dout  = 8'b10000001; // 3078 : 129 - 0x81
      12'hC07: dout  = 8'b10000001; // 3079 : 129 - 0x81
      12'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout  = 8'b01000001; // 3081 :  65 - 0x41
      12'hC0A: dout  = 8'b00100010; // 3082 :  34 - 0x22
      12'hC0B: dout  = 8'b00100010; // 3083 :  34 - 0x22
      12'hC0C: dout  = 8'b00011100; // 3084 :  28 - 0x1c
      12'hC0D: dout  = 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout  = 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout  = 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout  = 8'b11100011; // 3088 : 227 - 0xe3 -- Background 0xc1
      12'hC11: dout  = 8'b11110111; // 3089 : 247 - 0xf7
      12'hC12: dout  = 8'b11000001; // 3090 : 193 - 0xc1
      12'hC13: dout  = 8'b11000001; // 3091 : 193 - 0xc1
      12'hC14: dout  = 8'b11000001; // 3092 : 193 - 0xc1
      12'hC15: dout  = 8'b11000001; // 3093 : 193 - 0xc1
      12'hC16: dout  = 8'b11110111; // 3094 : 247 - 0xf7
      12'hC17: dout  = 8'b11100011; // 3095 : 227 - 0xe3
      12'hC18: dout  = 8'b11100011; // 3096 : 227 - 0xe3 -- plane 1
      12'hC19: dout  = 8'b00010100; // 3097 :  20 - 0x14
      12'hC1A: dout  = 8'b00111110; // 3098 :  62 - 0x3e
      12'hC1B: dout  = 8'b00111110; // 3099 :  62 - 0x3e
      12'hC1C: dout  = 8'b00111110; // 3100 :  62 - 0x3e
      12'hC1D: dout  = 8'b00111110; // 3101 :  62 - 0x3e
      12'hC1E: dout  = 8'b00010100; // 3102 :  20 - 0x14
      12'hC1F: dout  = 8'b11100011; // 3103 : 227 - 0xe3
      12'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Background 0xc2
      12'hC21: dout  = 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout  = 8'b00000111; // 3106 :   7 - 0x7
      12'hC23: dout  = 8'b00001111; // 3107 :  15 - 0xf
      12'hC24: dout  = 8'b00001100; // 3108 :  12 - 0xc
      12'hC25: dout  = 8'b00011011; // 3109 :  27 - 0x1b
      12'hC26: dout  = 8'b00011011; // 3110 :  27 - 0x1b
      12'hC27: dout  = 8'b00011011; // 3111 :  27 - 0x1b
      12'hC28: dout  = 8'b11111111; // 3112 : 255 - 0xff -- plane 1
      12'hC29: dout  = 8'b11111111; // 3113 : 255 - 0xff
      12'hC2A: dout  = 8'b11111000; // 3114 : 248 - 0xf8
      12'hC2B: dout  = 8'b11110000; // 3115 : 240 - 0xf0
      12'hC2C: dout  = 8'b11110000; // 3116 : 240 - 0xf0
      12'hC2D: dout  = 8'b11100000; // 3117 : 224 - 0xe0
      12'hC2E: dout  = 8'b11100000; // 3118 : 224 - 0xe0
      12'hC2F: dout  = 8'b11100000; // 3119 : 224 - 0xe0
      12'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Background 0xc3
      12'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout  = 8'b11100000; // 3122 : 224 - 0xe0
      12'hC33: dout  = 8'b11110000; // 3123 : 240 - 0xf0
      12'hC34: dout  = 8'b11110000; // 3124 : 240 - 0xf0
      12'hC35: dout  = 8'b11111000; // 3125 : 248 - 0xf8
      12'hC36: dout  = 8'b11111000; // 3126 : 248 - 0xf8
      12'hC37: dout  = 8'b11111000; // 3127 : 248 - 0xf8
      12'hC38: dout  = 8'b11111111; // 3128 : 255 - 0xff -- plane 1
      12'hC39: dout  = 8'b11111111; // 3129 : 255 - 0xff
      12'hC3A: dout  = 8'b01111111; // 3130 : 127 - 0x7f
      12'hC3B: dout  = 8'b00111111; // 3131 :  63 - 0x3f
      12'hC3C: dout  = 8'b00111111; // 3132 :  63 - 0x3f
      12'hC3D: dout  = 8'b10011111; // 3133 : 159 - 0x9f
      12'hC3E: dout  = 8'b10011111; // 3134 : 159 - 0x9f
      12'hC3F: dout  = 8'b10011111; // 3135 : 159 - 0x9f
      12'hC40: dout  = 8'b00011011; // 3136 :  27 - 0x1b -- Background 0xc4
      12'hC41: dout  = 8'b00011011; // 3137 :  27 - 0x1b
      12'hC42: dout  = 8'b00011011; // 3138 :  27 - 0x1b
      12'hC43: dout  = 8'b00011011; // 3139 :  27 - 0x1b
      12'hC44: dout  = 8'b00011011; // 3140 :  27 - 0x1b
      12'hC45: dout  = 8'b00001111; // 3141 :  15 - 0xf
      12'hC46: dout  = 8'b00001111; // 3142 :  15 - 0xf
      12'hC47: dout  = 8'b00000111; // 3143 :   7 - 0x7
      12'hC48: dout  = 8'b11100000; // 3144 : 224 - 0xe0 -- plane 1
      12'hC49: dout  = 8'b11100000; // 3145 : 224 - 0xe0
      12'hC4A: dout  = 8'b11100000; // 3146 : 224 - 0xe0
      12'hC4B: dout  = 8'b11100000; // 3147 : 224 - 0xe0
      12'hC4C: dout  = 8'b11100000; // 3148 : 224 - 0xe0
      12'hC4D: dout  = 8'b11110011; // 3149 : 243 - 0xf3
      12'hC4E: dout  = 8'b11110000; // 3150 : 240 - 0xf0
      12'hC4F: dout  = 8'b11111000; // 3151 : 248 - 0xf8
      12'hC50: dout  = 8'b11111000; // 3152 : 248 - 0xf8 -- Background 0xc5
      12'hC51: dout  = 8'b11111000; // 3153 : 248 - 0xf8
      12'hC52: dout  = 8'b11111000; // 3154 : 248 - 0xf8
      12'hC53: dout  = 8'b11111000; // 3155 : 248 - 0xf8
      12'hC54: dout  = 8'b11111000; // 3156 : 248 - 0xf8
      12'hC55: dout  = 8'b11110000; // 3157 : 240 - 0xf0
      12'hC56: dout  = 8'b11110000; // 3158 : 240 - 0xf0
      12'hC57: dout  = 8'b11100000; // 3159 : 224 - 0xe0
      12'hC58: dout  = 8'b10011111; // 3160 : 159 - 0x9f -- plane 1
      12'hC59: dout  = 8'b10011111; // 3161 : 159 - 0x9f
      12'hC5A: dout  = 8'b10011111; // 3162 : 159 - 0x9f
      12'hC5B: dout  = 8'b10011111; // 3163 : 159 - 0x9f
      12'hC5C: dout  = 8'b10011111; // 3164 : 159 - 0x9f
      12'hC5D: dout  = 8'b00111111; // 3165 :  63 - 0x3f
      12'hC5E: dout  = 8'b00111111; // 3166 :  63 - 0x3f
      12'hC5F: dout  = 8'b01111111; // 3167 : 127 - 0x7f
      12'hC60: dout  = 8'b11100000; // 3168 : 224 - 0xe0 -- Background 0xc6
      12'hC61: dout  = 8'b11111111; // 3169 : 255 - 0xff
      12'hC62: dout  = 8'b11111111; // 3170 : 255 - 0xff
      12'hC63: dout  = 8'b11111111; // 3171 : 255 - 0xff
      12'hC64: dout  = 8'b11111111; // 3172 : 255 - 0xff
      12'hC65: dout  = 8'b11111111; // 3173 : 255 - 0xff
      12'hC66: dout  = 8'b11111111; // 3174 : 255 - 0xff
      12'hC67: dout  = 8'b11111111; // 3175 : 255 - 0xff
      12'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout  = 8'b01110000; // 3177 : 112 - 0x70
      12'hC6A: dout  = 8'b00011111; // 3178 :  31 - 0x1f
      12'hC6B: dout  = 8'b00010000; // 3179 :  16 - 0x10
      12'hC6C: dout  = 8'b01110000; // 3180 : 112 - 0x70
      12'hC6D: dout  = 8'b01111111; // 3181 : 127 - 0x7f
      12'hC6E: dout  = 8'b01111111; // 3182 : 127 - 0x7f
      12'hC6F: dout  = 8'b01111111; // 3183 : 127 - 0x7f
      12'hC70: dout  = 8'b00000111; // 3184 :   7 - 0x7 -- Background 0xc7
      12'hC71: dout  = 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout  = 8'b11111111; // 3186 : 255 - 0xff
      12'hC73: dout  = 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout  = 8'b11111111; // 3188 : 255 - 0xff
      12'hC75: dout  = 8'b11111111; // 3189 : 255 - 0xff
      12'hC76: dout  = 8'b11111111; // 3190 : 255 - 0xff
      12'hC77: dout  = 8'b11111111; // 3191 : 255 - 0xff
      12'hC78: dout  = 8'b00000000; // 3192 :   0 - 0x0 -- plane 1
      12'hC79: dout  = 8'b00000011; // 3193 :   3 - 0x3
      12'hC7A: dout  = 8'b11111000; // 3194 : 248 - 0xf8
      12'hC7B: dout  = 8'b00000000; // 3195 :   0 - 0x0
      12'hC7C: dout  = 8'b00000011; // 3196 :   3 - 0x3
      12'hC7D: dout  = 8'b11111011; // 3197 : 251 - 0xfb
      12'hC7E: dout  = 8'b11111011; // 3198 : 251 - 0xfb
      12'hC7F: dout  = 8'b11111011; // 3199 : 251 - 0xfb
      12'hC80: dout  = 8'b11111111; // 3200 : 255 - 0xff -- Background 0xc8
      12'hC81: dout  = 8'b11111111; // 3201 : 255 - 0xff
      12'hC82: dout  = 8'b11111111; // 3202 : 255 - 0xff
      12'hC83: dout  = 8'b11111111; // 3203 : 255 - 0xff
      12'hC84: dout  = 8'b11111111; // 3204 : 255 - 0xff
      12'hC85: dout  = 8'b11111110; // 3205 : 254 - 0xfe
      12'hC86: dout  = 8'b11111111; // 3206 : 255 - 0xff
      12'hC87: dout  = 8'b11101111; // 3207 : 239 - 0xef
      12'hC88: dout  = 8'b01111100; // 3208 : 124 - 0x7c -- plane 1
      12'hC89: dout  = 8'b01111011; // 3209 : 123 - 0x7b
      12'hC8A: dout  = 8'b01110110; // 3210 : 118 - 0x76
      12'hC8B: dout  = 8'b01110101; // 3211 : 117 - 0x75
      12'hC8C: dout  = 8'b01110101; // 3212 : 117 - 0x75
      12'hC8D: dout  = 8'b01110111; // 3213 : 119 - 0x77
      12'hC8E: dout  = 8'b00010111; // 3214 :  23 - 0x17
      12'hC8F: dout  = 8'b01100111; // 3215 : 103 - 0x67
      12'hC90: dout  = 8'b11111111; // 3216 : 255 - 0xff -- Background 0xc9
      12'hC91: dout  = 8'b11011111; // 3217 : 223 - 0xdf
      12'hC92: dout  = 8'b11101111; // 3218 : 239 - 0xef
      12'hC93: dout  = 8'b10101111; // 3219 : 175 - 0xaf
      12'hC94: dout  = 8'b10101111; // 3220 : 175 - 0xaf
      12'hC95: dout  = 8'b01101111; // 3221 : 111 - 0x6f
      12'hC96: dout  = 8'b11101111; // 3222 : 239 - 0xef
      12'hC97: dout  = 8'b11100111; // 3223 : 231 - 0xe7
      12'hC98: dout  = 8'b00111011; // 3224 :  59 - 0x3b -- plane 1
      12'hC99: dout  = 8'b11111011; // 3225 : 251 - 0xfb
      12'hC9A: dout  = 8'b01111011; // 3226 : 123 - 0x7b
      12'hC9B: dout  = 8'b11111011; // 3227 : 251 - 0xfb
      12'hC9C: dout  = 8'b11111011; // 3228 : 251 - 0xfb
      12'hC9D: dout  = 8'b11110011; // 3229 : 243 - 0xf3
      12'hC9E: dout  = 8'b11111000; // 3230 : 248 - 0xf8
      12'hC9F: dout  = 8'b11110011; // 3231 : 243 - 0xf3
      12'hCA0: dout  = 8'b00011111; // 3232 :  31 - 0x1f -- Background 0xca
      12'hCA1: dout  = 8'b00011111; // 3233 :  31 - 0x1f
      12'hCA2: dout  = 8'b00111111; // 3234 :  63 - 0x3f
      12'hCA3: dout  = 8'b00111111; // 3235 :  63 - 0x3f
      12'hCA4: dout  = 8'b01110000; // 3236 : 112 - 0x70
      12'hCA5: dout  = 8'b01100011; // 3237 :  99 - 0x63
      12'hCA6: dout  = 8'b11100111; // 3238 : 231 - 0xe7
      12'hCA7: dout  = 8'b11100101; // 3239 : 229 - 0xe5
      12'hCA8: dout  = 8'b00001111; // 3240 :  15 - 0xf -- plane 1
      12'hCA9: dout  = 8'b00001111; // 3241 :  15 - 0xf
      12'hCAA: dout  = 8'b00011111; // 3242 :  31 - 0x1f
      12'hCAB: dout  = 8'b00011111; // 3243 :  31 - 0x1f
      12'hCAC: dout  = 8'b00111111; // 3244 :  63 - 0x3f
      12'hCAD: dout  = 8'b00111100; // 3245 :  60 - 0x3c
      12'hCAE: dout  = 8'b01111000; // 3246 : 120 - 0x78
      12'hCAF: dout  = 8'b01111010; // 3247 : 122 - 0x7a
      12'hCB0: dout  = 8'b11110000; // 3248 : 240 - 0xf0 -- Background 0xcb
      12'hCB1: dout  = 8'b11110000; // 3249 : 240 - 0xf0
      12'hCB2: dout  = 8'b11111000; // 3250 : 248 - 0xf8
      12'hCB3: dout  = 8'b11111000; // 3251 : 248 - 0xf8
      12'hCB4: dout  = 8'b00001100; // 3252 :  12 - 0xc
      12'hCB5: dout  = 8'b11000100; // 3253 : 196 - 0xc4
      12'hCB6: dout  = 8'b11100100; // 3254 : 228 - 0xe4
      12'hCB7: dout  = 8'b10100110; // 3255 : 166 - 0xa6
      12'hCB8: dout  = 8'b11111000; // 3256 : 248 - 0xf8 -- plane 1
      12'hCB9: dout  = 8'b11111000; // 3257 : 248 - 0xf8
      12'hCBA: dout  = 8'b11111100; // 3258 : 252 - 0xfc
      12'hCBB: dout  = 8'b11111100; // 3259 : 252 - 0xfc
      12'hCBC: dout  = 8'b11111110; // 3260 : 254 - 0xfe
      12'hCBD: dout  = 8'b00111110; // 3261 :  62 - 0x3e
      12'hCBE: dout  = 8'b00011110; // 3262 :  30 - 0x1e
      12'hCBF: dout  = 8'b01011111; // 3263 :  95 - 0x5f
      12'hCC0: dout  = 8'b11101001; // 3264 : 233 - 0xe9 -- Background 0xcc
      12'hCC1: dout  = 8'b11101001; // 3265 : 233 - 0xe9
      12'hCC2: dout  = 8'b11101001; // 3266 : 233 - 0xe9
      12'hCC3: dout  = 8'b11101111; // 3267 : 239 - 0xef
      12'hCC4: dout  = 8'b11100010; // 3268 : 226 - 0xe2
      12'hCC5: dout  = 8'b11100011; // 3269 : 227 - 0xe3
      12'hCC6: dout  = 8'b11110000; // 3270 : 240 - 0xf0
      12'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout  = 8'b01110110; // 3272 : 118 - 0x76 -- plane 1
      12'hCC9: dout  = 8'b01110110; // 3273 : 118 - 0x76
      12'hCCA: dout  = 8'b01110110; // 3274 : 118 - 0x76
      12'hCCB: dout  = 8'b01110000; // 3275 : 112 - 0x70
      12'hCCC: dout  = 8'b01111101; // 3276 : 125 - 0x7d
      12'hCCD: dout  = 8'b01111100; // 3277 : 124 - 0x7c
      12'hCCE: dout  = 8'b01111111; // 3278 : 127 - 0x7f
      12'hCCF: dout  = 8'b01111111; // 3279 : 127 - 0x7f
      12'hCD0: dout  = 8'b10010110; // 3280 : 150 - 0x96 -- Background 0xcd
      12'hCD1: dout  = 8'b10010110; // 3281 : 150 - 0x96
      12'hCD2: dout  = 8'b10010110; // 3282 : 150 - 0x96
      12'hCD3: dout  = 8'b11110110; // 3283 : 246 - 0xf6
      12'hCD4: dout  = 8'b01000110; // 3284 :  70 - 0x46
      12'hCD5: dout  = 8'b11000110; // 3285 : 198 - 0xc6
      12'hCD6: dout  = 8'b00001110; // 3286 :  14 - 0xe
      12'hCD7: dout  = 8'b11111110; // 3287 : 254 - 0xfe
      12'hCD8: dout  = 8'b01101111; // 3288 : 111 - 0x6f -- plane 1
      12'hCD9: dout  = 8'b01101111; // 3289 : 111 - 0x6f
      12'hCDA: dout  = 8'b01101111; // 3290 : 111 - 0x6f
      12'hCDB: dout  = 8'b00001111; // 3291 :  15 - 0xf
      12'hCDC: dout  = 8'b10111111; // 3292 : 191 - 0xbf
      12'hCDD: dout  = 8'b00111111; // 3293 :  63 - 0x3f
      12'hCDE: dout  = 8'b11111111; // 3294 : 255 - 0xff
      12'hCDF: dout  = 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout  = 8'b00000000; // 3296 :   0 - 0x0 -- Background 0xce
      12'hCE1: dout  = 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout  = 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout  = 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout  = 8'b00000000; // 3300 :   0 - 0x0
      12'hCE5: dout  = 8'b00000000; // 3301 :   0 - 0x0
      12'hCE6: dout  = 8'b01111110; // 3302 : 126 - 0x7e
      12'hCE7: dout  = 8'b00111100; // 3303 :  60 - 0x3c
      12'hCE8: dout  = 8'b00111100; // 3304 :  60 - 0x3c -- plane 1
      12'hCE9: dout  = 8'b01111110; // 3305 : 126 - 0x7e
      12'hCEA: dout  = 8'b01111110; // 3306 : 126 - 0x7e
      12'hCEB: dout  = 8'b11111111; // 3307 : 255 - 0xff
      12'hCEC: dout  = 8'b11111111; // 3308 : 255 - 0xff
      12'hCED: dout  = 8'b11111111; // 3309 : 255 - 0xff
      12'hCEE: dout  = 8'b01000010; // 3310 :  66 - 0x42
      12'hCEF: dout  = 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout  = 8'b00111100; // 3312 :  60 - 0x3c -- Background 0xcf
      12'hCF1: dout  = 8'b01000010; // 3313 :  66 - 0x42
      12'hCF2: dout  = 8'b10011001; // 3314 : 153 - 0x99
      12'hCF3: dout  = 8'b10100001; // 3315 : 161 - 0xa1
      12'hCF4: dout  = 8'b10100001; // 3316 : 161 - 0xa1
      12'hCF5: dout  = 8'b10011001; // 3317 : 153 - 0x99
      12'hCF6: dout  = 8'b01000010; // 3318 :  66 - 0x42
      12'hCF7: dout  = 8'b00111100; // 3319 :  60 - 0x3c
      12'hCF8: dout  = 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout  = 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout  = 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout  = 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout  = 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00001111; // 3328 :  15 - 0xf -- Background 0xd0
      12'hD01: dout  = 8'b00011111; // 3329 :  31 - 0x1f
      12'hD02: dout  = 8'b00011111; // 3330 :  31 - 0x1f
      12'hD03: dout  = 8'b00111111; // 3331 :  63 - 0x3f
      12'hD04: dout  = 8'b00111111; // 3332 :  63 - 0x3f
      12'hD05: dout  = 8'b01111111; // 3333 : 127 - 0x7f
      12'hD06: dout  = 8'b01111111; // 3334 : 127 - 0x7f
      12'hD07: dout  = 8'b01111111; // 3335 : 127 - 0x7f
      12'hD08: dout  = 8'b11110000; // 3336 : 240 - 0xf0 -- plane 1
      12'hD09: dout  = 8'b11100000; // 3337 : 224 - 0xe0
      12'hD0A: dout  = 8'b11100000; // 3338 : 224 - 0xe0
      12'hD0B: dout  = 8'b11000000; // 3339 : 192 - 0xc0
      12'hD0C: dout  = 8'b11000000; // 3340 : 192 - 0xc0
      12'hD0D: dout  = 8'b10000000; // 3341 : 128 - 0x80
      12'hD0E: dout  = 8'b10000000; // 3342 : 128 - 0x80
      12'hD0F: dout  = 8'b10000000; // 3343 : 128 - 0x80
      12'hD10: dout  = 8'b11110000; // 3344 : 240 - 0xf0 -- Background 0xd1
      12'hD11: dout  = 8'b11111000; // 3345 : 248 - 0xf8
      12'hD12: dout  = 8'b11111000; // 3346 : 248 - 0xf8
      12'hD13: dout  = 8'b11111100; // 3347 : 252 - 0xfc
      12'hD14: dout  = 8'b11111100; // 3348 : 252 - 0xfc
      12'hD15: dout  = 8'b11111110; // 3349 : 254 - 0xfe
      12'hD16: dout  = 8'b11111110; // 3350 : 254 - 0xfe
      12'hD17: dout  = 8'b11111110; // 3351 : 254 - 0xfe
      12'hD18: dout  = 8'b00001111; // 3352 :  15 - 0xf -- plane 1
      12'hD19: dout  = 8'b00000111; // 3353 :   7 - 0x7
      12'hD1A: dout  = 8'b00000111; // 3354 :   7 - 0x7
      12'hD1B: dout  = 8'b00000011; // 3355 :   3 - 0x3
      12'hD1C: dout  = 8'b00000011; // 3356 :   3 - 0x3
      12'hD1D: dout  = 8'b00000001; // 3357 :   1 - 0x1
      12'hD1E: dout  = 8'b00000001; // 3358 :   1 - 0x1
      12'hD1F: dout  = 8'b00000001; // 3359 :   1 - 0x1
      12'hD20: dout  = 8'b01111111; // 3360 : 127 - 0x7f -- Background 0xd2
      12'hD21: dout  = 8'b01111111; // 3361 : 127 - 0x7f
      12'hD22: dout  = 8'b00111111; // 3362 :  63 - 0x3f
      12'hD23: dout  = 8'b00111111; // 3363 :  63 - 0x3f
      12'hD24: dout  = 8'b00111111; // 3364 :  63 - 0x3f
      12'hD25: dout  = 8'b00111111; // 3365 :  63 - 0x3f
      12'hD26: dout  = 8'b00011111; // 3366 :  31 - 0x1f
      12'hD27: dout  = 8'b00011111; // 3367 :  31 - 0x1f
      12'hD28: dout  = 8'b10000000; // 3368 : 128 - 0x80 -- plane 1
      12'hD29: dout  = 8'b10000000; // 3369 : 128 - 0x80
      12'hD2A: dout  = 8'b11000000; // 3370 : 192 - 0xc0
      12'hD2B: dout  = 8'b11000000; // 3371 : 192 - 0xc0
      12'hD2C: dout  = 8'b11100000; // 3372 : 224 - 0xe0
      12'hD2D: dout  = 8'b11111000; // 3373 : 248 - 0xf8
      12'hD2E: dout  = 8'b11111110; // 3374 : 254 - 0xfe
      12'hD2F: dout  = 8'b11111111; // 3375 : 255 - 0xff
      12'hD30: dout  = 8'b11111110; // 3376 : 254 - 0xfe -- Background 0xd3
      12'hD31: dout  = 8'b11111111; // 3377 : 255 - 0xff
      12'hD32: dout  = 8'b11111111; // 3378 : 255 - 0xff
      12'hD33: dout  = 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout  = 8'b11111100; // 3380 : 252 - 0xfc
      12'hD35: dout  = 8'b11111100; // 3381 : 252 - 0xfc
      12'hD36: dout  = 8'b11111110; // 3382 : 254 - 0xfe
      12'hD37: dout  = 8'b11111110; // 3383 : 254 - 0xfe
      12'hD38: dout  = 8'b11111111; // 3384 : 255 - 0xff -- plane 1
      12'hD39: dout  = 8'b01111111; // 3385 : 127 - 0x7f
      12'hD3A: dout  = 8'b00011111; // 3386 :  31 - 0x1f
      12'hD3B: dout  = 8'b00000111; // 3387 :   7 - 0x7
      12'hD3C: dout  = 8'b00000011; // 3388 :   3 - 0x3
      12'hD3D: dout  = 8'b00000011; // 3389 :   3 - 0x3
      12'hD3E: dout  = 8'b00000001; // 3390 :   1 - 0x1
      12'hD3F: dout  = 8'b10000001; // 3391 : 129 - 0x81
      12'hD40: dout  = 8'b01111111; // 3392 : 127 - 0x7f -- Background 0xd4
      12'hD41: dout  = 8'b01111111; // 3393 : 127 - 0x7f
      12'hD42: dout  = 8'b01111111; // 3394 : 127 - 0x7f
      12'hD43: dout  = 8'b00111111; // 3395 :  63 - 0x3f
      12'hD44: dout  = 8'b00111111; // 3396 :  63 - 0x3f
      12'hD45: dout  = 8'b00111111; // 3397 :  63 - 0x3f
      12'hD46: dout  = 8'b00111111; // 3398 :  63 - 0x3f
      12'hD47: dout  = 8'b00011111; // 3399 :  31 - 0x1f
      12'hD48: dout  = 8'b10000000; // 3400 : 128 - 0x80 -- plane 1
      12'hD49: dout  = 8'b10000000; // 3401 : 128 - 0x80
      12'hD4A: dout  = 8'b10000000; // 3402 : 128 - 0x80
      12'hD4B: dout  = 8'b11000000; // 3403 : 192 - 0xc0
      12'hD4C: dout  = 8'b11000000; // 3404 : 192 - 0xc0
      12'hD4D: dout  = 8'b11100000; // 3405 : 224 - 0xe0
      12'hD4E: dout  = 8'b11100000; // 3406 : 224 - 0xe0
      12'hD4F: dout  = 8'b11110000; // 3407 : 240 - 0xf0
      12'hD50: dout  = 8'b11111110; // 3408 : 254 - 0xfe -- Background 0xd5
      12'hD51: dout  = 8'b11111110; // 3409 : 254 - 0xfe
      12'hD52: dout  = 8'b11111111; // 3410 : 255 - 0xff
      12'hD53: dout  = 8'b11111111; // 3411 : 255 - 0xff
      12'hD54: dout  = 8'b11111111; // 3412 : 255 - 0xff
      12'hD55: dout  = 8'b11111111; // 3413 : 255 - 0xff
      12'hD56: dout  = 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout  = 8'b11111110; // 3415 : 254 - 0xfe
      12'hD58: dout  = 8'b00000001; // 3416 :   1 - 0x1 -- plane 1
      12'hD59: dout  = 8'b00000001; // 3417 :   1 - 0x1
      12'hD5A: dout  = 8'b00000001; // 3418 :   1 - 0x1
      12'hD5B: dout  = 8'b00000011; // 3419 :   3 - 0x3
      12'hD5C: dout  = 8'b00000011; // 3420 :   3 - 0x3
      12'hD5D: dout  = 8'b00000111; // 3421 :   7 - 0x7
      12'hD5E: dout  = 8'b00000111; // 3422 :   7 - 0x7
      12'hD5F: dout  = 8'b00001111; // 3423 :  15 - 0xf
      12'hD60: dout  = 8'b00011111; // 3424 :  31 - 0x1f -- Background 0xd6
      12'hD61: dout  = 8'b00001111; // 3425 :  15 - 0xf
      12'hD62: dout  = 8'b00001111; // 3426 :  15 - 0xf
      12'hD63: dout  = 8'b00000111; // 3427 :   7 - 0x7
      12'hD64: dout  = 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout  = 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout  = 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout  = 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout  = 8'b11111111; // 3432 : 255 - 0xff -- plane 1
      12'hD69: dout  = 8'b11111111; // 3433 : 255 - 0xff
      12'hD6A: dout  = 8'b11111111; // 3434 : 255 - 0xff
      12'hD6B: dout  = 8'b11111111; // 3435 : 255 - 0xff
      12'hD6C: dout  = 8'b11111111; // 3436 : 255 - 0xff
      12'hD6D: dout  = 8'b11111111; // 3437 : 255 - 0xff
      12'hD6E: dout  = 8'b11111111; // 3438 : 255 - 0xff
      12'hD6F: dout  = 8'b11111111; // 3439 : 255 - 0xff
      12'hD70: dout  = 8'b11111110; // 3440 : 254 - 0xfe -- Background 0xd7
      12'hD71: dout  = 8'b11111100; // 3441 : 252 - 0xfc
      12'hD72: dout  = 8'b11111100; // 3442 : 252 - 0xfc
      12'hD73: dout  = 8'b11111000; // 3443 : 248 - 0xf8
      12'hD74: dout  = 8'b00000000; // 3444 :   0 - 0x0
      12'hD75: dout  = 8'b00000000; // 3445 :   0 - 0x0
      12'hD76: dout  = 8'b00000000; // 3446 :   0 - 0x0
      12'hD77: dout  = 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout  = 8'b11111111; // 3448 : 255 - 0xff -- plane 1
      12'hD79: dout  = 8'b11111111; // 3449 : 255 - 0xff
      12'hD7A: dout  = 8'b11111111; // 3450 : 255 - 0xff
      12'hD7B: dout  = 8'b11111111; // 3451 : 255 - 0xff
      12'hD7C: dout  = 8'b11111111; // 3452 : 255 - 0xff
      12'hD7D: dout  = 8'b11111111; // 3453 : 255 - 0xff
      12'hD7E: dout  = 8'b11111111; // 3454 : 255 - 0xff
      12'hD7F: dout  = 8'b11111111; // 3455 : 255 - 0xff
      12'hD80: dout  = 8'b01111110; // 3456 : 126 - 0x7e -- Background 0xd8
      12'hD81: dout  = 8'b01111110; // 3457 : 126 - 0x7e
      12'hD82: dout  = 8'b01111110; // 3458 : 126 - 0x7e
      12'hD83: dout  = 8'b01111110; // 3459 : 126 - 0x7e
      12'hD84: dout  = 8'b01111111; // 3460 : 127 - 0x7f
      12'hD85: dout  = 8'b01111111; // 3461 : 127 - 0x7f
      12'hD86: dout  = 8'b01111111; // 3462 : 127 - 0x7f
      12'hD87: dout  = 8'b01111111; // 3463 : 127 - 0x7f
      12'hD88: dout  = 8'b10000001; // 3464 : 129 - 0x81 -- plane 1
      12'hD89: dout  = 8'b10000001; // 3465 : 129 - 0x81
      12'hD8A: dout  = 8'b10000001; // 3466 : 129 - 0x81
      12'hD8B: dout  = 8'b10000001; // 3467 : 129 - 0x81
      12'hD8C: dout  = 8'b10000001; // 3468 : 129 - 0x81
      12'hD8D: dout  = 8'b10000001; // 3469 : 129 - 0x81
      12'hD8E: dout  = 8'b10000001; // 3470 : 129 - 0x81
      12'hD8F: dout  = 8'b10000001; // 3471 : 129 - 0x81
      12'hD90: dout  = 8'b11111111; // 3472 : 255 - 0xff -- Background 0xd9
      12'hD91: dout  = 8'b11111111; // 3473 : 255 - 0xff
      12'hD92: dout  = 8'b11111111; // 3474 : 255 - 0xff
      12'hD93: dout  = 8'b11111111; // 3475 : 255 - 0xff
      12'hD94: dout  = 8'b11111111; // 3476 : 255 - 0xff
      12'hD95: dout  = 8'b11111111; // 3477 : 255 - 0xff
      12'hD96: dout  = 8'b11111111; // 3478 : 255 - 0xff
      12'hD97: dout  = 8'b11111110; // 3479 : 254 - 0xfe
      12'hD98: dout  = 8'b00000001; // 3480 :   1 - 0x1 -- plane 1
      12'hD99: dout  = 8'b00000001; // 3481 :   1 - 0x1
      12'hD9A: dout  = 8'b00000001; // 3482 :   1 - 0x1
      12'hD9B: dout  = 8'b00000011; // 3483 :   3 - 0x3
      12'hD9C: dout  = 8'b00000011; // 3484 :   3 - 0x3
      12'hD9D: dout  = 8'b00000111; // 3485 :   7 - 0x7
      12'hD9E: dout  = 8'b00000111; // 3486 :   7 - 0x7
      12'hD9F: dout  = 8'b00001111; // 3487 :  15 - 0xf
      12'hDA0: dout  = 8'b11111110; // 3488 : 254 - 0xfe -- Background 0xda
      12'hDA1: dout  = 8'b11111110; // 3489 : 254 - 0xfe
      12'hDA2: dout  = 8'b11111110; // 3490 : 254 - 0xfe
      12'hDA3: dout  = 8'b11111110; // 3491 : 254 - 0xfe
      12'hDA4: dout  = 8'b11111111; // 3492 : 255 - 0xff
      12'hDA5: dout  = 8'b11111111; // 3493 : 255 - 0xff
      12'hDA6: dout  = 8'b11111111; // 3494 : 255 - 0xff
      12'hDA7: dout  = 8'b11111111; // 3495 : 255 - 0xff
      12'hDA8: dout  = 8'b00000001; // 3496 :   1 - 0x1 -- plane 1
      12'hDA9: dout  = 8'b00000001; // 3497 :   1 - 0x1
      12'hDAA: dout  = 8'b00000001; // 3498 :   1 - 0x1
      12'hDAB: dout  = 8'b00000001; // 3499 :   1 - 0x1
      12'hDAC: dout  = 8'b00000001; // 3500 :   1 - 0x1
      12'hDAD: dout  = 8'b00000001; // 3501 :   1 - 0x1
      12'hDAE: dout  = 8'b00000001; // 3502 :   1 - 0x1
      12'hDAF: dout  = 8'b00000001; // 3503 :   1 - 0x1
      12'hDB0: dout  = 8'b01111111; // 3504 : 127 - 0x7f -- Background 0xdb
      12'hDB1: dout  = 8'b01111111; // 3505 : 127 - 0x7f
      12'hDB2: dout  = 8'b01111111; // 3506 : 127 - 0x7f
      12'hDB3: dout  = 8'b01111111; // 3507 : 127 - 0x7f
      12'hDB4: dout  = 8'b01111111; // 3508 : 127 - 0x7f
      12'hDB5: dout  = 8'b01111111; // 3509 : 127 - 0x7f
      12'hDB6: dout  = 8'b01111111; // 3510 : 127 - 0x7f
      12'hDB7: dout  = 8'b01111111; // 3511 : 127 - 0x7f
      12'hDB8: dout  = 8'b10000001; // 3512 : 129 - 0x81 -- plane 1
      12'hDB9: dout  = 8'b10000001; // 3513 : 129 - 0x81
      12'hDBA: dout  = 8'b10000001; // 3514 : 129 - 0x81
      12'hDBB: dout  = 8'b10000001; // 3515 : 129 - 0x81
      12'hDBC: dout  = 8'b10000001; // 3516 : 129 - 0x81
      12'hDBD: dout  = 8'b10000001; // 3517 : 129 - 0x81
      12'hDBE: dout  = 8'b10000001; // 3518 : 129 - 0x81
      12'hDBF: dout  = 8'b10000001; // 3519 : 129 - 0x81
      12'hDC0: dout  = 8'b11111111; // 3520 : 255 - 0xff -- Background 0xdc
      12'hDC1: dout  = 8'b11111111; // 3521 : 255 - 0xff
      12'hDC2: dout  = 8'b11111111; // 3522 : 255 - 0xff
      12'hDC3: dout  = 8'b11111111; // 3523 : 255 - 0xff
      12'hDC4: dout  = 8'b11111100; // 3524 : 252 - 0xfc
      12'hDC5: dout  = 8'b11111110; // 3525 : 254 - 0xfe
      12'hDC6: dout  = 8'b11111110; // 3526 : 254 - 0xfe
      12'hDC7: dout  = 8'b01111110; // 3527 : 126 - 0x7e
      12'hDC8: dout  = 8'b11111111; // 3528 : 255 - 0xff -- plane 1
      12'hDC9: dout  = 8'b00000011; // 3529 :   3 - 0x3
      12'hDCA: dout  = 8'b00000011; // 3530 :   3 - 0x3
      12'hDCB: dout  = 8'b00000011; // 3531 :   3 - 0x3
      12'hDCC: dout  = 8'b00000011; // 3532 :   3 - 0x3
      12'hDCD: dout  = 8'b00000011; // 3533 :   3 - 0x3
      12'hDCE: dout  = 8'b00000011; // 3534 :   3 - 0x3
      12'hDCF: dout  = 8'b11111111; // 3535 : 255 - 0xff
      12'hDD0: dout  = 8'b11111111; // 3536 : 255 - 0xff -- Background 0xdd
      12'hDD1: dout  = 8'b11111111; // 3537 : 255 - 0xff
      12'hDD2: dout  = 8'b11111111; // 3538 : 255 - 0xff
      12'hDD3: dout  = 8'b11111111; // 3539 : 255 - 0xff
      12'hDD4: dout  = 8'b00000000; // 3540 :   0 - 0x0
      12'hDD5: dout  = 8'b00000000; // 3541 :   0 - 0x0
      12'hDD6: dout  = 8'b00000000; // 3542 :   0 - 0x0
      12'hDD7: dout  = 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout  = 8'b11111111; // 3544 : 255 - 0xff -- plane 1
      12'hDD9: dout  = 8'b11111111; // 3545 : 255 - 0xff
      12'hDDA: dout  = 8'b11111111; // 3546 : 255 - 0xff
      12'hDDB: dout  = 8'b11111111; // 3547 : 255 - 0xff
      12'hDDC: dout  = 8'b11111111; // 3548 : 255 - 0xff
      12'hDDD: dout  = 8'b11111111; // 3549 : 255 - 0xff
      12'hDDE: dout  = 8'b11111111; // 3550 : 255 - 0xff
      12'hDDF: dout  = 8'b11111111; // 3551 : 255 - 0xff
      12'hDE0: dout  = 8'b01111111; // 3552 : 127 - 0x7f -- Background 0xde
      12'hDE1: dout  = 8'b01111111; // 3553 : 127 - 0x7f
      12'hDE2: dout  = 8'b01111111; // 3554 : 127 - 0x7f
      12'hDE3: dout  = 8'b01111111; // 3555 : 127 - 0x7f
      12'hDE4: dout  = 8'b01111111; // 3556 : 127 - 0x7f
      12'hDE5: dout  = 8'b01111111; // 3557 : 127 - 0x7f
      12'hDE6: dout  = 8'b01111111; // 3558 : 127 - 0x7f
      12'hDE7: dout  = 8'b01111111; // 3559 : 127 - 0x7f
      12'hDE8: dout  = 8'b10000000; // 3560 : 128 - 0x80 -- plane 1
      12'hDE9: dout  = 8'b10000000; // 3561 : 128 - 0x80
      12'hDEA: dout  = 8'b10000000; // 3562 : 128 - 0x80
      12'hDEB: dout  = 8'b10000000; // 3563 : 128 - 0x80
      12'hDEC: dout  = 8'b10000000; // 3564 : 128 - 0x80
      12'hDED: dout  = 8'b10000000; // 3565 : 128 - 0x80
      12'hDEE: dout  = 8'b10000000; // 3566 : 128 - 0x80
      12'hDEF: dout  = 8'b10000000; // 3567 : 128 - 0x80
      12'hDF0: dout  = 8'b11111111; // 3568 : 255 - 0xff -- Background 0xdf
      12'hDF1: dout  = 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout  = 8'b11111111; // 3570 : 255 - 0xff
      12'hDF3: dout  = 8'b11111111; // 3571 : 255 - 0xff
      12'hDF4: dout  = 8'b11111111; // 3572 : 255 - 0xff
      12'hDF5: dout  = 8'b11111111; // 3573 : 255 - 0xff
      12'hDF6: dout  = 8'b11111111; // 3574 : 255 - 0xff
      12'hDF7: dout  = 8'b11111110; // 3575 : 254 - 0xfe
      12'hDF8: dout  = 8'b00000001; // 3576 :   1 - 0x1 -- plane 1
      12'hDF9: dout  = 8'b00000001; // 3577 :   1 - 0x1
      12'hDFA: dout  = 8'b00000001; // 3578 :   1 - 0x1
      12'hDFB: dout  = 8'b00000011; // 3579 :   3 - 0x3
      12'hDFC: dout  = 8'b00000111; // 3580 :   7 - 0x7
      12'hDFD: dout  = 8'b00000011; // 3581 :   3 - 0x3
      12'hDFE: dout  = 8'b00000001; // 3582 :   1 - 0x1
      12'hDFF: dout  = 8'b00000001; // 3583 :   1 - 0x1
      12'hE00: dout  = 8'b01111110; // 3584 : 126 - 0x7e -- Background 0xe0
      12'hE01: dout  = 8'b01111110; // 3585 : 126 - 0x7e
      12'hE02: dout  = 8'b01111111; // 3586 : 127 - 0x7f
      12'hE03: dout  = 8'b01111111; // 3587 : 127 - 0x7f
      12'hE04: dout  = 8'b01111111; // 3588 : 127 - 0x7f
      12'hE05: dout  = 8'b01111111; // 3589 : 127 - 0x7f
      12'hE06: dout  = 8'b01111111; // 3590 : 127 - 0x7f
      12'hE07: dout  = 8'b01111111; // 3591 : 127 - 0x7f
      12'hE08: dout  = 8'b10000001; // 3592 : 129 - 0x81 -- plane 1
      12'hE09: dout  = 8'b10000001; // 3593 : 129 - 0x81
      12'hE0A: dout  = 8'b10000001; // 3594 : 129 - 0x81
      12'hE0B: dout  = 8'b10000001; // 3595 : 129 - 0x81
      12'hE0C: dout  = 8'b10000001; // 3596 : 129 - 0x81
      12'hE0D: dout  = 8'b10000001; // 3597 : 129 - 0x81
      12'hE0E: dout  = 8'b10000001; // 3598 : 129 - 0x81
      12'hE0F: dout  = 8'b10000001; // 3599 : 129 - 0x81
      12'hE10: dout  = 8'b00111111; // 3600 :  63 - 0x3f -- Background 0xe1
      12'hE11: dout  = 8'b00111111; // 3601 :  63 - 0x3f
      12'hE12: dout  = 8'b00111111; // 3602 :  63 - 0x3f
      12'hE13: dout  = 8'b00111111; // 3603 :  63 - 0x3f
      12'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout  = 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout  = 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout  = 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout  = 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout  = 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout  = 8'b11111111; // 3610 : 255 - 0xff
      12'hE1B: dout  = 8'b11111111; // 3611 : 255 - 0xff
      12'hE1C: dout  = 8'b11111111; // 3612 : 255 - 0xff
      12'hE1D: dout  = 8'b11111111; // 3613 : 255 - 0xff
      12'hE1E: dout  = 8'b11111111; // 3614 : 255 - 0xff
      12'hE1F: dout  = 8'b11111111; // 3615 : 255 - 0xff
      12'hE20: dout  = 8'b01111110; // 3616 : 126 - 0x7e -- Background 0xe2
      12'hE21: dout  = 8'b01111100; // 3617 : 124 - 0x7c
      12'hE22: dout  = 8'b01111100; // 3618 : 124 - 0x7c
      12'hE23: dout  = 8'b01111000; // 3619 : 120 - 0x78
      12'hE24: dout  = 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout  = 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout  = 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout  = 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout  = 8'b11111111; // 3624 : 255 - 0xff -- plane 1
      12'hE29: dout  = 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout  = 8'b11111111; // 3626 : 255 - 0xff
      12'hE2B: dout  = 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout  = 8'b11111111; // 3628 : 255 - 0xff
      12'hE2D: dout  = 8'b11111111; // 3629 : 255 - 0xff
      12'hE2E: dout  = 8'b11111111; // 3630 : 255 - 0xff
      12'hE2F: dout  = 8'b11111111; // 3631 : 255 - 0xff
      12'hE30: dout  = 8'b11111110; // 3632 : 254 - 0xfe -- Background 0xe3
      12'hE31: dout  = 8'b11111110; // 3633 : 254 - 0xfe
      12'hE32: dout  = 8'b11111111; // 3634 : 255 - 0xff
      12'hE33: dout  = 8'b11111111; // 3635 : 255 - 0xff
      12'hE34: dout  = 8'b01111111; // 3636 : 127 - 0x7f
      12'hE35: dout  = 8'b01111111; // 3637 : 127 - 0x7f
      12'hE36: dout  = 8'b01111111; // 3638 : 127 - 0x7f
      12'hE37: dout  = 8'b01111111; // 3639 : 127 - 0x7f
      12'hE38: dout  = 8'b10000001; // 3640 : 129 - 0x81 -- plane 1
      12'hE39: dout  = 8'b10000001; // 3641 : 129 - 0x81
      12'hE3A: dout  = 8'b10000001; // 3642 : 129 - 0x81
      12'hE3B: dout  = 8'b10000001; // 3643 : 129 - 0x81
      12'hE3C: dout  = 8'b10000001; // 3644 : 129 - 0x81
      12'hE3D: dout  = 8'b10000001; // 3645 : 129 - 0x81
      12'hE3E: dout  = 8'b10000001; // 3646 : 129 - 0x81
      12'hE3F: dout  = 8'b10000001; // 3647 : 129 - 0x81
      12'hE40: dout  = 8'b01111111; // 3648 : 127 - 0x7f -- Background 0xe4
      12'hE41: dout  = 8'b01111111; // 3649 : 127 - 0x7f
      12'hE42: dout  = 8'b00111111; // 3650 :  63 - 0x3f
      12'hE43: dout  = 8'b00111111; // 3651 :  63 - 0x3f
      12'hE44: dout  = 8'b00111111; // 3652 :  63 - 0x3f
      12'hE45: dout  = 8'b00111111; // 3653 :  63 - 0x3f
      12'hE46: dout  = 8'b00011111; // 3654 :  31 - 0x1f
      12'hE47: dout  = 8'b00011111; // 3655 :  31 - 0x1f
      12'hE48: dout  = 8'b10000000; // 3656 : 128 - 0x80 -- plane 1
      12'hE49: dout  = 8'b10000000; // 3657 : 128 - 0x80
      12'hE4A: dout  = 8'b11000000; // 3658 : 192 - 0xc0
      12'hE4B: dout  = 8'b11000000; // 3659 : 192 - 0xc0
      12'hE4C: dout  = 8'b11100000; // 3660 : 224 - 0xe0
      12'hE4D: dout  = 8'b11111000; // 3661 : 248 - 0xf8
      12'hE4E: dout  = 8'b11111110; // 3662 : 254 - 0xfe
      12'hE4F: dout  = 8'b11111111; // 3663 : 255 - 0xff
      12'hE50: dout  = 8'b00111111; // 3664 :  63 - 0x3f -- Background 0xe5
      12'hE51: dout  = 8'b10111111; // 3665 : 191 - 0xbf
      12'hE52: dout  = 8'b11111111; // 3666 : 255 - 0xff
      12'hE53: dout  = 8'b11111111; // 3667 : 255 - 0xff
      12'hE54: dout  = 8'b11111100; // 3668 : 252 - 0xfc
      12'hE55: dout  = 8'b11111100; // 3669 : 252 - 0xfc
      12'hE56: dout  = 8'b11111110; // 3670 : 254 - 0xfe
      12'hE57: dout  = 8'b11111110; // 3671 : 254 - 0xfe
      12'hE58: dout  = 8'b11111111; // 3672 : 255 - 0xff -- plane 1
      12'hE59: dout  = 8'b01111111; // 3673 : 127 - 0x7f
      12'hE5A: dout  = 8'b00011111; // 3674 :  31 - 0x1f
      12'hE5B: dout  = 8'b00000111; // 3675 :   7 - 0x7
      12'hE5C: dout  = 8'b00000011; // 3676 :   3 - 0x3
      12'hE5D: dout  = 8'b00000011; // 3677 :   3 - 0x3
      12'hE5E: dout  = 8'b00000001; // 3678 :   1 - 0x1
      12'hE5F: dout  = 8'b10000001; // 3679 : 129 - 0x81
      12'hE60: dout  = 8'b01111111; // 3680 : 127 - 0x7f -- Background 0xe6
      12'hE61: dout  = 8'b01111111; // 3681 : 127 - 0x7f
      12'hE62: dout  = 8'b01111110; // 3682 : 126 - 0x7e
      12'hE63: dout  = 8'b01111110; // 3683 : 126 - 0x7e
      12'hE64: dout  = 8'b01111111; // 3684 : 127 - 0x7f
      12'hE65: dout  = 8'b01111111; // 3685 : 127 - 0x7f
      12'hE66: dout  = 8'b01111111; // 3686 : 127 - 0x7f
      12'hE67: dout  = 8'b01111111; // 3687 : 127 - 0x7f
      12'hE68: dout  = 8'b10000001; // 3688 : 129 - 0x81 -- plane 1
      12'hE69: dout  = 8'b10000001; // 3689 : 129 - 0x81
      12'hE6A: dout  = 8'b10000001; // 3690 : 129 - 0x81
      12'hE6B: dout  = 8'b10000001; // 3691 : 129 - 0x81
      12'hE6C: dout  = 8'b10000001; // 3692 : 129 - 0x81
      12'hE6D: dout  = 8'b10000001; // 3693 : 129 - 0x81
      12'hE6E: dout  = 8'b10000001; // 3694 : 129 - 0x81
      12'hE6F: dout  = 8'b10000001; // 3695 : 129 - 0x81
      12'hE70: dout  = 8'b01111110; // 3696 : 126 - 0x7e -- Background 0xe7
      12'hE71: dout  = 8'b01111110; // 3697 : 126 - 0x7e
      12'hE72: dout  = 8'b01111110; // 3698 : 126 - 0x7e
      12'hE73: dout  = 8'b01111110; // 3699 : 126 - 0x7e
      12'hE74: dout  = 8'b01111111; // 3700 : 127 - 0x7f
      12'hE75: dout  = 8'b01111111; // 3701 : 127 - 0x7f
      12'hE76: dout  = 8'b01111111; // 3702 : 127 - 0x7f
      12'hE77: dout  = 8'b01111111; // 3703 : 127 - 0x7f
      12'hE78: dout  = 8'b10000001; // 3704 : 129 - 0x81 -- plane 1
      12'hE79: dout  = 8'b10000001; // 3705 : 129 - 0x81
      12'hE7A: dout  = 8'b10000001; // 3706 : 129 - 0x81
      12'hE7B: dout  = 8'b10000001; // 3707 : 129 - 0x81
      12'hE7C: dout  = 8'b10000001; // 3708 : 129 - 0x81
      12'hE7D: dout  = 8'b10000001; // 3709 : 129 - 0x81
      12'hE7E: dout  = 8'b10000001; // 3710 : 129 - 0x81
      12'hE7F: dout  = 8'b10000001; // 3711 : 129 - 0x81
      12'hE80: dout  = 8'b10000001; // 3712 : 129 - 0x81 -- Background 0xe8
      12'hE81: dout  = 8'b11000011; // 3713 : 195 - 0xc3
      12'hE82: dout  = 8'b11000011; // 3714 : 195 - 0xc3
      12'hE83: dout  = 8'b11100111; // 3715 : 231 - 0xe7
      12'hE84: dout  = 8'b11100111; // 3716 : 231 - 0xe7
      12'hE85: dout  = 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout  = 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout  = 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout  = 8'b01111110; // 3720 : 126 - 0x7e -- plane 1
      12'hE89: dout  = 8'b00111100; // 3721 :  60 - 0x3c
      12'hE8A: dout  = 8'b00111100; // 3722 :  60 - 0x3c
      12'hE8B: dout  = 8'b00011000; // 3723 :  24 - 0x18
      12'hE8C: dout  = 8'b00011000; // 3724 :  24 - 0x18
      12'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout  = 8'b00001111; // 3728 :  15 - 0xf -- Background 0xe9
      12'hE91: dout  = 8'b01000011; // 3729 :  67 - 0x43
      12'hE92: dout  = 8'b01011011; // 3730 :  91 - 0x5b
      12'hE93: dout  = 8'b01010011; // 3731 :  83 - 0x53
      12'hE94: dout  = 8'b00110001; // 3732 :  49 - 0x31
      12'hE95: dout  = 8'b00011001; // 3733 :  25 - 0x19
      12'hE96: dout  = 8'b00001111; // 3734 :  15 - 0xf
      12'hE97: dout  = 8'b00000111; // 3735 :   7 - 0x7
      12'hE98: dout  = 8'b11110010; // 3736 : 242 - 0xf2 -- plane 1
      12'hE99: dout  = 8'b11111110; // 3737 : 254 - 0xfe
      12'hE9A: dout  = 8'b11111110; // 3738 : 254 - 0xfe
      12'hE9B: dout  = 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout  = 8'b11111111; // 3740 : 255 - 0xff
      12'hE9D: dout  = 8'b11101111; // 3741 : 239 - 0xef
      12'hE9E: dout  = 8'b11110111; // 3742 : 247 - 0xf7
      12'hE9F: dout  = 8'b11111000; // 3743 : 248 - 0xf8
      12'hEA0: dout  = 8'b11000001; // 3744 : 193 - 0xc1 -- Background 0xea
      12'hEA1: dout  = 8'b11000011; // 3745 : 195 - 0xc3
      12'hEA2: dout  = 8'b11000110; // 3746 : 198 - 0xc6
      12'hEA3: dout  = 8'b10000100; // 3747 : 132 - 0x84
      12'hEA4: dout  = 8'b11111100; // 3748 : 252 - 0xfc
      12'hEA5: dout  = 8'b11111100; // 3749 : 252 - 0xfc
      12'hEA6: dout  = 8'b00001110; // 3750 :  14 - 0xe
      12'hEA7: dout  = 8'b00000010; // 3751 :   2 - 0x2
      12'hEA8: dout  = 8'b10111111; // 3752 : 191 - 0xbf -- plane 1
      12'hEA9: dout  = 8'b10111110; // 3753 : 190 - 0xbe
      12'hEAA: dout  = 8'b10111101; // 3754 : 189 - 0xbd
      12'hEAB: dout  = 8'b01111011; // 3755 : 123 - 0x7b
      12'hEAC: dout  = 8'b01111011; // 3756 : 123 - 0x7b
      12'hEAD: dout  = 8'b00000111; // 3757 :   7 - 0x7
      12'hEAE: dout  = 8'b11110011; // 3758 : 243 - 0xf3
      12'hEAF: dout  = 8'b11111101; // 3759 : 253 - 0xfd
      12'hEB0: dout  = 8'b00010000; // 3760 :  16 - 0x10 -- Background 0xeb
      12'hEB1: dout  = 8'b00100000; // 3761 :  32 - 0x20
      12'hEB2: dout  = 8'b00100010; // 3762 :  34 - 0x22
      12'hEB3: dout  = 8'b10111010; // 3763 : 186 - 0xba
      12'hEB4: dout  = 8'b11100110; // 3764 : 230 - 0xe6
      12'hEB5: dout  = 8'b11100001; // 3765 : 225 - 0xe1
      12'hEB6: dout  = 8'b11000000; // 3766 : 192 - 0xc0
      12'hEB7: dout  = 8'b11000000; // 3767 : 192 - 0xc0
      12'hEB8: dout  = 8'b11111111; // 3768 : 255 - 0xff -- plane 1
      12'hEB9: dout  = 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout  = 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout  = 8'b01100111; // 3771 : 103 - 0x67
      12'hEBC: dout  = 8'b01011001; // 3772 :  89 - 0x59
      12'hEBD: dout  = 8'b10011110; // 3773 : 158 - 0x9e
      12'hEBE: dout  = 8'b10111111; // 3774 : 191 - 0xbf
      12'hEBF: dout  = 8'b10111111; // 3775 : 191 - 0xbf
      12'hEC0: dout  = 8'b00100000; // 3776 :  32 - 0x20 -- Background 0xec
      12'hEC1: dout  = 8'b10100110; // 3777 : 166 - 0xa6
      12'hEC2: dout  = 8'b01010100; // 3778 :  84 - 0x54
      12'hEC3: dout  = 8'b00100110; // 3779 :  38 - 0x26
      12'hEC4: dout  = 8'b00100000; // 3780 :  32 - 0x20
      12'hEC5: dout  = 8'b11000110; // 3781 : 198 - 0xc6
      12'hEC6: dout  = 8'b01010100; // 3782 :  84 - 0x54
      12'hEC7: dout  = 8'b00100110; // 3783 :  38 - 0x26
      12'hEC8: dout  = 8'b00100000; // 3784 :  32 - 0x20 -- plane 1
      12'hEC9: dout  = 8'b11100110; // 3785 : 230 - 0xe6
      12'hECA: dout  = 8'b01010100; // 3786 :  84 - 0x54
      12'hECB: dout  = 8'b00100110; // 3787 :  38 - 0x26
      12'hECC: dout  = 8'b00100001; // 3788 :  33 - 0x21
      12'hECD: dout  = 8'b00000110; // 3789 :   6 - 0x6
      12'hECE: dout  = 8'b01010100; // 3790 :  84 - 0x54
      12'hECF: dout  = 8'b00100110; // 3791 :  38 - 0x26
      12'hED0: dout  = 8'b00100000; // 3792 :  32 - 0x20 -- Background 0xed
      12'hED1: dout  = 8'b10000101; // 3793 : 133 - 0x85
      12'hED2: dout  = 8'b00000001; // 3794 :   1 - 0x1
      12'hED3: dout  = 8'b01000100; // 3795 :  68 - 0x44
      12'hED4: dout  = 8'b00100000; // 3796 :  32 - 0x20
      12'hED5: dout  = 8'b10000110; // 3797 : 134 - 0x86
      12'hED6: dout  = 8'b01010100; // 3798 :  84 - 0x54
      12'hED7: dout  = 8'b01001000; // 3799 :  72 - 0x48
      12'hED8: dout  = 8'b00100000; // 3800 :  32 - 0x20 -- plane 1
      12'hED9: dout  = 8'b10011010; // 3801 : 154 - 0x9a
      12'hEDA: dout  = 8'b00000001; // 3802 :   1 - 0x1
      12'hEDB: dout  = 8'b01001001; // 3803 :  73 - 0x49
      12'hEDC: dout  = 8'b00100000; // 3804 :  32 - 0x20
      12'hEDD: dout  = 8'b10100101; // 3805 : 165 - 0xa5
      12'hEDE: dout  = 8'b11001001; // 3806 : 201 - 0xc9
      12'hEDF: dout  = 8'b01000110; // 3807 :  70 - 0x46
      12'hEE0: dout  = 8'b00100000; // 3808 :  32 - 0x20 -- Background 0xee
      12'hEE1: dout  = 8'b10111010; // 3809 : 186 - 0xba
      12'hEE2: dout  = 8'b11001001; // 3810 : 201 - 0xc9
      12'hEE3: dout  = 8'b01001010; // 3811 :  74 - 0x4a
      12'hEE4: dout  = 8'b00100000; // 3812 :  32 - 0x20
      12'hEE5: dout  = 8'b10100110; // 3813 : 166 - 0xa6
      12'hEE6: dout  = 8'b00001010; // 3814 :  10 - 0xa
      12'hEE7: dout  = 8'b11010000; // 3815 : 208 - 0xd0
      12'hEE8: dout  = 8'b11010001; // 3816 : 209 - 0xd1 -- plane 1
      12'hEE9: dout  = 8'b11011000; // 3817 : 216 - 0xd8
      12'hEEA: dout  = 8'b11011000; // 3818 : 216 - 0xd8
      12'hEEB: dout  = 8'b11011110; // 3819 : 222 - 0xde
      12'hEEC: dout  = 8'b11010001; // 3820 : 209 - 0xd1
      12'hEED: dout  = 8'b11010000; // 3821 : 208 - 0xd0
      12'hEEE: dout  = 8'b11011010; // 3822 : 218 - 0xda
      12'hEEF: dout  = 8'b11011110; // 3823 : 222 - 0xde
      12'hEF0: dout  = 8'b11010001; // 3824 : 209 - 0xd1 -- Background 0xef
      12'hEF1: dout  = 8'b00100000; // 3825 :  32 - 0x20
      12'hEF2: dout  = 8'b11000110; // 3826 : 198 - 0xc6
      12'hEF3: dout  = 8'b00001010; // 3827 :  10 - 0xa
      12'hEF4: dout  = 8'b11010010; // 3828 : 210 - 0xd2
      12'hEF5: dout  = 8'b11010011; // 3829 : 211 - 0xd3
      12'hEF6: dout  = 8'b11011011; // 3830 : 219 - 0xdb
      12'hEF7: dout  = 8'b11011011; // 3831 : 219 - 0xdb
      12'hEF8: dout  = 8'b11011011; // 3832 : 219 - 0xdb -- plane 1
      12'hEF9: dout  = 8'b11011001; // 3833 : 217 - 0xd9
      12'hEFA: dout  = 8'b11011011; // 3834 : 219 - 0xdb
      12'hEFB: dout  = 8'b11011100; // 3835 : 220 - 0xdc
      12'hEFC: dout  = 8'b11011011; // 3836 : 219 - 0xdb
      12'hEFD: dout  = 8'b11011111; // 3837 : 223 - 0xdf
      12'hEFE: dout  = 8'b00100000; // 3838 :  32 - 0x20
      12'hEFF: dout  = 8'b11100110; // 3839 : 230 - 0xe6
      12'hF00: dout  = 8'b00001010; // 3840 :  10 - 0xa -- Background 0xf0
      12'hF01: dout  = 8'b11010100; // 3841 : 212 - 0xd4
      12'hF02: dout  = 8'b11010101; // 3842 : 213 - 0xd5
      12'hF03: dout  = 8'b11010100; // 3843 : 212 - 0xd4
      12'hF04: dout  = 8'b11011001; // 3844 : 217 - 0xd9
      12'hF05: dout  = 8'b11011011; // 3845 : 219 - 0xdb
      12'hF06: dout  = 8'b11100010; // 3846 : 226 - 0xe2
      12'hF07: dout  = 8'b11010100; // 3847 : 212 - 0xd4
      12'hF08: dout  = 8'b11011010; // 3848 : 218 - 0xda -- plane 1
      12'hF09: dout  = 8'b11011011; // 3849 : 219 - 0xdb
      12'hF0A: dout  = 8'b11100000; // 3850 : 224 - 0xe0
      12'hF0B: dout  = 8'b00100001; // 3851 :  33 - 0x21
      12'hF0C: dout  = 8'b00000110; // 3852 :   6 - 0x6
      12'hF0D: dout  = 8'b00001010; // 3853 :  10 - 0xa
      12'hF0E: dout  = 8'b11010110; // 3854 : 214 - 0xd6
      12'hF0F: dout  = 8'b11010111; // 3855 : 215 - 0xd7
      12'hF10: dout  = 8'b11010110; // 3856 : 214 - 0xd6 -- Background 0xf1
      12'hF11: dout  = 8'b11010111; // 3857 : 215 - 0xd7
      12'hF12: dout  = 8'b11100001; // 3858 : 225 - 0xe1
      12'hF13: dout  = 8'b00100110; // 3859 :  38 - 0x26
      12'hF14: dout  = 8'b11010110; // 3860 : 214 - 0xd6
      12'hF15: dout  = 8'b11011101; // 3861 : 221 - 0xdd
      12'hF16: dout  = 8'b11100001; // 3862 : 225 - 0xe1
      12'hF17: dout  = 8'b11100001; // 3863 : 225 - 0xe1
      12'hF18: dout  = 8'b00100001; // 3864 :  33 - 0x21 -- plane 1
      12'hF19: dout  = 8'b00100110; // 3865 :  38 - 0x26
      12'hF1A: dout  = 8'b00010100; // 3866 :  20 - 0x14
      12'hF1B: dout  = 8'b11010000; // 3867 : 208 - 0xd0
      12'hF1C: dout  = 8'b11101000; // 3868 : 232 - 0xe8
      12'hF1D: dout  = 8'b11010001; // 3869 : 209 - 0xd1
      12'hF1E: dout  = 8'b11010000; // 3870 : 208 - 0xd0
      12'hF1F: dout  = 8'b11010001; // 3871 : 209 - 0xd1
      12'hF20: dout  = 8'b11011110; // 3872 : 222 - 0xde -- Background 0xf2
      12'hF21: dout  = 8'b11010001; // 3873 : 209 - 0xd1
      12'hF22: dout  = 8'b11011000; // 3874 : 216 - 0xd8
      12'hF23: dout  = 8'b11010000; // 3875 : 208 - 0xd0
      12'hF24: dout  = 8'b11010001; // 3876 : 209 - 0xd1
      12'hF25: dout  = 8'b00100110; // 3877 :  38 - 0x26
      12'hF26: dout  = 8'b11011110; // 3878 : 222 - 0xde
      12'hF27: dout  = 8'b11010001; // 3879 : 209 - 0xd1
      12'hF28: dout  = 8'b11011110; // 3880 : 222 - 0xde -- plane 1
      12'hF29: dout  = 8'b11010001; // 3881 : 209 - 0xd1
      12'hF2A: dout  = 8'b11010000; // 3882 : 208 - 0xd0
      12'hF2B: dout  = 8'b11010001; // 3883 : 209 - 0xd1
      12'hF2C: dout  = 8'b11010000; // 3884 : 208 - 0xd0
      12'hF2D: dout  = 8'b11010001; // 3885 : 209 - 0xd1
      12'hF2E: dout  = 8'b00100110; // 3886 :  38 - 0x26
      12'hF2F: dout  = 8'b00100001; // 3887 :  33 - 0x21
      12'hF30: dout  = 8'b01000110; // 3888 :  70 - 0x46 -- Background 0xf3
      12'hF31: dout  = 8'b00010100; // 3889 :  20 - 0x14
      12'hF32: dout  = 8'b11011011; // 3890 : 219 - 0xdb
      12'hF33: dout  = 8'b01000010; // 3891 :  66 - 0x42
      12'hF34: dout  = 8'b01000010; // 3892 :  66 - 0x42
      12'hF35: dout  = 8'b11011011; // 3893 : 219 - 0xdb
      12'hF36: dout  = 8'b01000010; // 3894 :  66 - 0x42
      12'hF37: dout  = 8'b11011011; // 3895 : 219 - 0xdb
      12'hF38: dout  = 8'b01000010; // 3896 :  66 - 0x42 -- plane 1
      12'hF39: dout  = 8'b11011011; // 3897 : 219 - 0xdb
      12'hF3A: dout  = 8'b11011011; // 3898 : 219 - 0xdb
      12'hF3B: dout  = 8'b01000010; // 3899 :  66 - 0x42
      12'hF3C: dout  = 8'b00100110; // 3900 :  38 - 0x26
      12'hF3D: dout  = 8'b11011011; // 3901 : 219 - 0xdb
      12'hF3E: dout  = 8'b01000010; // 3902 :  66 - 0x42
      12'hF3F: dout  = 8'b11011011; // 3903 : 219 - 0xdb
      12'hF40: dout  = 8'b01000010; // 3904 :  66 - 0x42 -- Background 0xf4
      12'hF41: dout  = 8'b11011011; // 3905 : 219 - 0xdb
      12'hF42: dout  = 8'b01000010; // 3906 :  66 - 0x42
      12'hF43: dout  = 8'b11011011; // 3907 : 219 - 0xdb
      12'hF44: dout  = 8'b01000010; // 3908 :  66 - 0x42
      12'hF45: dout  = 8'b00100110; // 3909 :  38 - 0x26
      12'hF46: dout  = 8'b00100001; // 3910 :  33 - 0x21
      12'hF47: dout  = 8'b01100110; // 3911 : 102 - 0x66
      12'hF48: dout  = 8'b01000110; // 3912 :  70 - 0x46 -- plane 1
      12'hF49: dout  = 8'b11011011; // 3913 : 219 - 0xdb
      12'hF4A: dout  = 8'b00100001; // 3914 :  33 - 0x21
      12'hF4B: dout  = 8'b01101100; // 3915 : 108 - 0x6c
      12'hF4C: dout  = 8'b00001110; // 3916 :  14 - 0xe
      12'hF4D: dout  = 8'b11011111; // 3917 : 223 - 0xdf
      12'hF4E: dout  = 8'b11011011; // 3918 : 219 - 0xdb
      12'hF4F: dout  = 8'b11011011; // 3919 : 219 - 0xdb
      12'hF50: dout  = 8'b11011011; // 3920 : 219 - 0xdb -- Background 0xf5
      12'hF51: dout  = 8'b00100110; // 3921 :  38 - 0x26
      12'hF52: dout  = 8'b11011011; // 3922 : 219 - 0xdb
      12'hF53: dout  = 8'b11011111; // 3923 : 223 - 0xdf
      12'hF54: dout  = 8'b11011011; // 3924 : 219 - 0xdb
      12'hF55: dout  = 8'b11011111; // 3925 : 223 - 0xdf
      12'hF56: dout  = 8'b11011011; // 3926 : 219 - 0xdb
      12'hF57: dout  = 8'b11011011; // 3927 : 219 - 0xdb
      12'hF58: dout  = 8'b11100100; // 3928 : 228 - 0xe4 -- plane 1
      12'hF59: dout  = 8'b11100101; // 3929 : 229 - 0xe5
      12'hF5A: dout  = 8'b00100110; // 3930 :  38 - 0x26
      12'hF5B: dout  = 8'b00100001; // 3931 :  33 - 0x21
      12'hF5C: dout  = 8'b10000110; // 3932 : 134 - 0x86
      12'hF5D: dout  = 8'b00010100; // 3933 :  20 - 0x14
      12'hF5E: dout  = 8'b11011011; // 3934 : 219 - 0xdb
      12'hF5F: dout  = 8'b11011011; // 3935 : 219 - 0xdb
      12'hF60: dout  = 8'b11011011; // 3936 : 219 - 0xdb -- Background 0xf6
      12'hF61: dout  = 8'b11011110; // 3937 : 222 - 0xde
      12'hF62: dout  = 8'b01000011; // 3938 :  67 - 0x43
      12'hF63: dout  = 8'b11011011; // 3939 : 219 - 0xdb
      12'hF64: dout  = 8'b11100000; // 3940 : 224 - 0xe0
      12'hF65: dout  = 8'b11011011; // 3941 : 219 - 0xdb
      12'hF66: dout  = 8'b11011011; // 3942 : 219 - 0xdb
      12'hF67: dout  = 8'b11011011; // 3943 : 219 - 0xdb
      12'hF68: dout  = 8'b00100110; // 3944 :  38 - 0x26 -- plane 1
      12'hF69: dout  = 8'b11011011; // 3945 : 219 - 0xdb
      12'hF6A: dout  = 8'b11100011; // 3946 : 227 - 0xe3
      12'hF6B: dout  = 8'b11011011; // 3947 : 219 - 0xdb
      12'hF6C: dout  = 8'b11100000; // 3948 : 224 - 0xe0
      12'hF6D: dout  = 8'b11011011; // 3949 : 219 - 0xdb
      12'hF6E: dout  = 8'b11011011; // 3950 : 219 - 0xdb
      12'hF6F: dout  = 8'b11100110; // 3951 : 230 - 0xe6
      12'hF70: dout  = 8'b11100011; // 3952 : 227 - 0xe3 -- Background 0xf7
      12'hF71: dout  = 8'b00100110; // 3953 :  38 - 0x26
      12'hF72: dout  = 8'b00100001; // 3954 :  33 - 0x21
      12'hF73: dout  = 8'b10100110; // 3955 : 166 - 0xa6
      12'hF74: dout  = 8'b00010100; // 3956 :  20 - 0x14
      12'hF75: dout  = 8'b11011011; // 3957 : 219 - 0xdb
      12'hF76: dout  = 8'b11011011; // 3958 : 219 - 0xdb
      12'hF77: dout  = 8'b11011011; // 3959 : 219 - 0xdb
      12'hF78: dout  = 8'b11011011; // 3960 : 219 - 0xdb -- plane 1
      12'hF79: dout  = 8'b01000010; // 3961 :  66 - 0x42
      12'hF7A: dout  = 8'b11011011; // 3962 : 219 - 0xdb
      12'hF7B: dout  = 8'b11011011; // 3963 : 219 - 0xdb
      12'hF7C: dout  = 8'b11011011; // 3964 : 219 - 0xdb
      12'hF7D: dout  = 8'b11010100; // 3965 : 212 - 0xd4
      12'hF7E: dout  = 8'b11011001; // 3966 : 217 - 0xd9
      12'hF7F: dout  = 8'b00100110; // 3967 :  38 - 0x26
      12'hF80: dout  = 8'b11011011; // 3968 : 219 - 0xdb -- Background 0xf8
      12'hF81: dout  = 8'b11011001; // 3969 : 217 - 0xd9
      12'hF82: dout  = 8'b11011011; // 3970 : 219 - 0xdb
      12'hF83: dout  = 8'b11011011; // 3971 : 219 - 0xdb
      12'hF84: dout  = 8'b11010100; // 3972 : 212 - 0xd4
      12'hF85: dout  = 8'b11011001; // 3973 : 217 - 0xd9
      12'hF86: dout  = 8'b11010100; // 3974 : 212 - 0xd4
      12'hF87: dout  = 8'b11011001; // 3975 : 217 - 0xd9
      12'hF88: dout  = 8'b11100111; // 3976 : 231 - 0xe7 -- plane 1
      12'hF89: dout  = 8'b00100001; // 3977 :  33 - 0x21
      12'hF8A: dout  = 8'b11000101; // 3978 : 197 - 0xc5
      12'hF8B: dout  = 8'b00010110; // 3979 :  22 - 0x16
      12'hF8C: dout  = 8'b01011111; // 3980 :  95 - 0x5f
      12'hF8D: dout  = 8'b10010101; // 3981 : 149 - 0x95
      12'hF8E: dout  = 8'b10010101; // 3982 : 149 - 0x95
      12'hF8F: dout  = 8'b10010101; // 3983 : 149 - 0x95
      12'hF90: dout  = 8'b10010101; // 3984 : 149 - 0x95 -- Background 0xf9
      12'hF91: dout  = 8'b10010101; // 3985 : 149 - 0x95
      12'hF92: dout  = 8'b10010101; // 3986 : 149 - 0x95
      12'hF93: dout  = 8'b10010101; // 3987 : 149 - 0x95
      12'hF94: dout  = 8'b10010101; // 3988 : 149 - 0x95
      12'hF95: dout  = 8'b10010111; // 3989 : 151 - 0x97
      12'hF96: dout  = 8'b10011000; // 3990 : 152 - 0x98
      12'hF97: dout  = 8'b01111000; // 3991 : 120 - 0x78
      12'hF98: dout  = 8'b10010101; // 3992 : 149 - 0x95 -- plane 1
      12'hF99: dout  = 8'b10010110; // 3993 : 150 - 0x96
      12'hF9A: dout  = 8'b10010101; // 3994 : 149 - 0x95
      12'hF9B: dout  = 8'b10010101; // 3995 : 149 - 0x95
      12'hF9C: dout  = 8'b10010111; // 3996 : 151 - 0x97
      12'hF9D: dout  = 8'b10011000; // 3997 : 152 - 0x98
      12'hF9E: dout  = 8'b10010111; // 3998 : 151 - 0x97
      12'hF9F: dout  = 8'b10011000; // 3999 : 152 - 0x98
      12'hFA0: dout  = 8'b10010101; // 4000 : 149 - 0x95 -- Background 0xfa
      12'hFA1: dout  = 8'b01111010; // 4001 : 122 - 0x7a
      12'hFA2: dout  = 8'b00100001; // 4002 :  33 - 0x21
      12'hFA3: dout  = 8'b11101101; // 4003 : 237 - 0xed
      12'hFA4: dout  = 8'b00001110; // 4004 :  14 - 0xe
      12'hFA5: dout  = 8'b11001111; // 4005 : 207 - 0xcf
      12'hFA6: dout  = 8'b00000001; // 4006 :   1 - 0x1
      12'hFA7: dout  = 8'b00001001; // 4007 :   9 - 0x9
      12'hFA8: dout  = 8'b00001000; // 4008 :   8 - 0x8 -- plane 1
      12'hFA9: dout  = 8'b00000101; // 4009 :   5 - 0x5
      12'hFAA: dout  = 8'b00100100; // 4010 :  36 - 0x24
      12'hFAB: dout  = 8'b00010111; // 4011 :  23 - 0x17
      12'hFAC: dout  = 8'b00010010; // 4012 :  18 - 0x12
      12'hFAD: dout  = 8'b00010111; // 4013 :  23 - 0x17
      12'hFAE: dout  = 8'b00011101; // 4014 :  29 - 0x1d
      12'hFAF: dout  = 8'b00001110; // 4015 :  14 - 0xe
      12'hFB0: dout  = 8'b00010111; // 4016 :  23 - 0x17 -- Background 0xfb
      12'hFB1: dout  = 8'b00001101; // 4017 :  13 - 0xd
      12'hFB2: dout  = 8'b00011000; // 4018 :  24 - 0x18
      12'hFB3: dout  = 8'b00100010; // 4019 :  34 - 0x22
      12'hFB4: dout  = 8'b01001011; // 4020 :  75 - 0x4b
      12'hFB5: dout  = 8'b00001101; // 4021 :  13 - 0xd
      12'hFB6: dout  = 8'b00000001; // 4022 :   1 - 0x1
      12'hFB7: dout  = 8'b00100100; // 4023 :  36 - 0x24
      12'hFB8: dout  = 8'b00011001; // 4024 :  25 - 0x19 -- plane 1
      12'hFB9: dout  = 8'b00010101; // 4025 :  21 - 0x15
      12'hFBA: dout  = 8'b00001010; // 4026 :  10 - 0xa
      12'hFBB: dout  = 8'b00100010; // 4027 :  34 - 0x22
      12'hFBC: dout  = 8'b00001110; // 4028 :  14 - 0xe
      12'hFBD: dout  = 8'b00011011; // 4029 :  27 - 0x1b
      12'hFBE: dout  = 8'b00100100; // 4030 :  36 - 0x24
      12'hFBF: dout  = 8'b00010000; // 4031 :  16 - 0x10
      12'hFC0: dout  = 8'b00001010; // 4032 :  10 - 0xa -- Background 0xfc
      12'hFC1: dout  = 8'b00010110; // 4033 :  22 - 0x16
      12'hFC2: dout  = 8'b00001110; // 4034 :  14 - 0xe
      12'hFC3: dout  = 8'b00100010; // 4035 :  34 - 0x22
      12'hFC4: dout  = 8'b10001011; // 4036 : 139 - 0x8b
      12'hFC5: dout  = 8'b00001101; // 4037 :  13 - 0xd
      12'hFC6: dout  = 8'b00000010; // 4038 :   2 - 0x2
      12'hFC7: dout  = 8'b00100100; // 4039 :  36 - 0x24
      12'hFC8: dout  = 8'b00011001; // 4040 :  25 - 0x19 -- plane 1
      12'hFC9: dout  = 8'b00010101; // 4041 :  21 - 0x15
      12'hFCA: dout  = 8'b00001010; // 4042 :  10 - 0xa
      12'hFCB: dout  = 8'b00100010; // 4043 :  34 - 0x22
      12'hFCC: dout  = 8'b00001110; // 4044 :  14 - 0xe
      12'hFCD: dout  = 8'b00011011; // 4045 :  27 - 0x1b
      12'hFCE: dout  = 8'b00100100; // 4046 :  36 - 0x24
      12'hFCF: dout  = 8'b00010000; // 4047 :  16 - 0x10
      12'hFD0: dout  = 8'b00001010; // 4048 :  10 - 0xa -- Background 0xfd
      12'hFD1: dout  = 8'b00010110; // 4049 :  22 - 0x16
      12'hFD2: dout  = 8'b00001110; // 4050 :  14 - 0xe
      12'hFD3: dout  = 8'b00100010; // 4051 :  34 - 0x22
      12'hFD4: dout  = 8'b11101100; // 4052 : 236 - 0xec
      12'hFD5: dout  = 8'b00000100; // 4053 :   4 - 0x4
      12'hFD6: dout  = 8'b00011101; // 4054 :  29 - 0x1d
      12'hFD7: dout  = 8'b00011000; // 4055 :  24 - 0x18
      12'hFD8: dout  = 8'b00011001; // 4056 :  25 - 0x19 -- plane 1
      12'hFD9: dout  = 8'b00101000; // 4057 :  40 - 0x28
      12'hFDA: dout  = 8'b00100010; // 4058 :  34 - 0x22
      12'hFDB: dout  = 8'b11110110; // 4059 : 246 - 0xf6
      12'hFDC: dout  = 8'b00000001; // 4060 :   1 - 0x1
      12'hFDD: dout  = 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout  = 8'b00100011; // 4062 :  35 - 0x23
      12'hFDF: dout  = 8'b11001001; // 4063 : 201 - 0xc9
      12'hFE0: dout  = 8'b01010110; // 4064 :  86 - 0x56 -- Background 0xfe
      12'hFE1: dout  = 8'b01010101; // 4065 :  85 - 0x55
      12'hFE2: dout  = 8'b00100011; // 4066 :  35 - 0x23
      12'hFE3: dout  = 8'b11100010; // 4067 : 226 - 0xe2
      12'hFE4: dout  = 8'b00000100; // 4068 :   4 - 0x4
      12'hFE5: dout  = 8'b10011001; // 4069 : 153 - 0x99
      12'hFE6: dout  = 8'b10101010; // 4070 : 170 - 0xaa
      12'hFE7: dout  = 8'b10101010; // 4071 : 170 - 0xaa
      12'hFE8: dout  = 8'b10101010; // 4072 : 170 - 0xaa -- plane 1
      12'hFE9: dout  = 8'b00100011; // 4073 :  35 - 0x23
      12'hFEA: dout  = 8'b11101010; // 4074 : 234 - 0xea
      12'hFEB: dout  = 8'b00000100; // 4075 :   4 - 0x4
      12'hFEC: dout  = 8'b10011001; // 4076 : 153 - 0x99
      12'hFED: dout  = 8'b10101010; // 4077 : 170 - 0xaa
      12'hFEE: dout  = 8'b10101010; // 4078 : 170 - 0xaa
      12'hFEF: dout  = 8'b10101010; // 4079 : 170 - 0xaa
      12'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Background 0xff
      12'hFF1: dout  = 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout  = 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout  = 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout  = 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout  = 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout  = 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout  = 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout  = 8'b11111111; // 4088 : 255 - 0xff -- plane 1
      12'hFF9: dout  = 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout  = 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout  = 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout  = 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout  = 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout  = 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout  = 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
