--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Pattern Table 0---------
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x1
    "00111000", --   17 - 0x11  :   56 - 0x38
    "01111100", --   18 - 0x12  :  124 - 0x7c
    "11111110", --   19 - 0x13  :  254 - 0xfe
    "11111110", --   20 - 0x14  :  254 - 0xfe
    "11111110", --   21 - 0x15  :  254 - 0xfe
    "01111100", --   22 - 0x16  :  124 - 0x7c
    "00111000", --   23 - 0x17  :   56 - 0x38
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00111000", --   25 - 0x19  :   56 - 0x38
    "01111100", --   26 - 0x1a  :  124 - 0x7c
    "11111110", --   27 - 0x1b  :  254 - 0xfe
    "11111110", --   28 - 0x1c  :  254 - 0xfe
    "11111110", --   29 - 0x1d  :  254 - 0xfe
    "01111100", --   30 - 0x1e  :  124 - 0x7c
    "00111000", --   31 - 0x1f  :   56 - 0x38
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00011000", --   51 - 0x33  :   24 - 0x18
    "00011000", --   52 - 0x34  :   24 - 0x18
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00011000", --   59 - 0x3b  :   24 - 0x18
    "00011000", --   60 - 0x3c  :   24 - 0x18
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00001111", --   88 - 0x58  :   15 - 0xf
    "00001111", --   89 - 0x59  :   15 - 0xf
    "00001111", --   90 - 0x5a  :   15 - 0xf
    "00001111", --   91 - 0x5b  :   15 - 0xf
    "00001111", --   92 - 0x5c  :   15 - 0xf
    "00001111", --   93 - 0x5d  :   15 - 0xf
    "00001111", --   94 - 0x5e  :   15 - 0xf
    "00001111", --   95 - 0x5f  :   15 - 0xf
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11110000", --  104 - 0x68  :  240 - 0xf0
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11110000", --  106 - 0x6a  :  240 - 0xf0
    "11110000", --  107 - 0x6b  :  240 - 0xf0
    "11110000", --  108 - 0x6c  :  240 - 0xf0
    "11110000", --  109 - 0x6d  :  240 - 0xf0
    "11110000", --  110 - 0x6e  :  240 - 0xf0
    "11110000", --  111 - 0x6f  :  240 - 0xf0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0x7
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x8
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x9
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00011000", --  147 - 0x93  :   24 - 0x18
    "00011000", --  148 - 0x94  :   24 - 0x18
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00011000", --  155 - 0x9b  :   24 - 0x18
    "00011000", --  156 - 0x9c  :   24 - 0x18
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0xa
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0xb
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0xd
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  257 - 0x101  :    0 - 0x0
    "11111111", --  258 - 0x102  :  255 - 0xff
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "11111111", --  261 - 0x105  :  255 - 0xff
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00100100", --  272 - 0x110  :   36 - 0x24 -- Sprite 0x11
    "00100100", --  273 - 0x111  :   36 - 0x24
    "00100100", --  274 - 0x112  :   36 - 0x24
    "00100100", --  275 - 0x113  :   36 - 0x24
    "00100100", --  276 - 0x114  :   36 - 0x24
    "00100100", --  277 - 0x115  :   36 - 0x24
    "00100100", --  278 - 0x116  :   36 - 0x24
    "00100100", --  279 - 0x117  :   36 - 0x24
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00100100", --  288 - 0x120  :   36 - 0x24 -- Sprite 0x12
    "00100100", --  289 - 0x121  :   36 - 0x24
    "11000011", --  290 - 0x122  :  195 - 0xc3
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "11111111", --  293 - 0x125  :  255 - 0xff
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  305 - 0x131  :    0 - 0x0
    "11111111", --  306 - 0x132  :  255 - 0xff
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "11000011", --  309 - 0x135  :  195 - 0xc3
    "00100100", --  310 - 0x136  :   36 - 0x24
    "00100100", --  311 - 0x137  :   36 - 0x24
    "00000000", --  312 - 0x138  :    0 - 0x0
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00100100", --  320 - 0x140  :   36 - 0x24 -- Sprite 0x14
    "00100100", --  321 - 0x141  :   36 - 0x24
    "11000100", --  322 - 0x142  :  196 - 0xc4
    "00000100", --  323 - 0x143  :    4 - 0x4
    "00000100", --  324 - 0x144  :    4 - 0x4
    "11000100", --  325 - 0x145  :  196 - 0xc4
    "00100100", --  326 - 0x146  :   36 - 0x24
    "00100100", --  327 - 0x147  :   36 - 0x24
    "00000000", --  328 - 0x148  :    0 - 0x0
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00100100", --  336 - 0x150  :   36 - 0x24 -- Sprite 0x15
    "00100100", --  337 - 0x151  :   36 - 0x24
    "00100011", --  338 - 0x152  :   35 - 0x23
    "00100000", --  339 - 0x153  :   32 - 0x20
    "00100000", --  340 - 0x154  :   32 - 0x20
    "00100011", --  341 - 0x155  :   35 - 0x23
    "00100100", --  342 - 0x156  :   36 - 0x24
    "00100100", --  343 - 0x157  :   36 - 0x24
    "00000000", --  344 - 0x158  :    0 - 0x0
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00001111", --  354 - 0x162  :   15 - 0xf
    "00010000", --  355 - 0x163  :   16 - 0x10
    "11110000", --  356 - 0x164  :  240 - 0xf0
    "00001111", --  357 - 0x165  :   15 - 0xf
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x17
    "00000000", --  369 - 0x171  :    0 - 0x0
    "11110000", --  370 - 0x172  :  240 - 0xf0
    "00001000", --  371 - 0x173  :    8 - 0x8
    "00001111", --  372 - 0x174  :   15 - 0xf
    "11110000", --  373 - 0x175  :  240 - 0xf0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  385 - 0x181  :    0 - 0x0
    "11110000", --  386 - 0x182  :  240 - 0xf0
    "00001000", --  387 - 0x183  :    8 - 0x8
    "00001000", --  388 - 0x184  :    8 - 0x8
    "11110000", --  389 - 0x185  :  240 - 0xf0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x19
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00001111", --  402 - 0x192  :   15 - 0xf
    "00010000", --  403 - 0x193  :   16 - 0x10
    "00010000", --  404 - 0x194  :   16 - 0x10
    "00001111", --  405 - 0x195  :   15 - 0xf
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00100100", --  416 - 0x1a0  :   36 - 0x24 -- Sprite 0x1a
    "00100100", --  417 - 0x1a1  :   36 - 0x24
    "00100100", --  418 - 0x1a2  :   36 - 0x24
    "00100100", --  419 - 0x1a3  :   36 - 0x24
    "00011000", --  420 - 0x1a4  :   24 - 0x18
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00011000", --  435 - 0x1b3  :   24 - 0x18
    "00100100", --  436 - 0x1b4  :   36 - 0x24
    "00100100", --  437 - 0x1b5  :   36 - 0x24
    "00100100", --  438 - 0x1b6  :   36 - 0x24
    "00100100", --  439 - 0x1b7  :   36 - 0x24
    "00000000", --  440 - 0x1b8  :    0 - 0x0
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00100100", --  448 - 0x1c0  :   36 - 0x24 -- Sprite 0x1c
    "00100100", --  449 - 0x1c1  :   36 - 0x24
    "11000100", --  450 - 0x1c2  :  196 - 0xc4
    "00000100", --  451 - 0x1c3  :    4 - 0x4
    "00001000", --  452 - 0x1c4  :    8 - 0x8
    "11110000", --  453 - 0x1c5  :  240 - 0xf0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x1d
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "11110000", --  466 - 0x1d2  :  240 - 0xf0
    "00001000", --  467 - 0x1d3  :    8 - 0x8
    "00000100", --  468 - 0x1d4  :    4 - 0x4
    "11000100", --  469 - 0x1d5  :  196 - 0xc4
    "00100100", --  470 - 0x1d6  :   36 - 0x24
    "00100100", --  471 - 0x1d7  :   36 - 0x24
    "00000000", --  472 - 0x1d8  :    0 - 0x0
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00100100", --  480 - 0x1e0  :   36 - 0x24 -- Sprite 0x1e
    "00100100", --  481 - 0x1e1  :   36 - 0x24
    "00100011", --  482 - 0x1e2  :   35 - 0x23
    "00100000", --  483 - 0x1e3  :   32 - 0x20
    "00010000", --  484 - 0x1e4  :   16 - 0x10
    "00001111", --  485 - 0x1e5  :   15 - 0xf
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00001111", --  498 - 0x1f2  :   15 - 0xf
    "00010000", --  499 - 0x1f3  :   16 - 0x10
    "00100000", --  500 - 0x1f4  :   32 - 0x20
    "00100011", --  501 - 0x1f5  :   35 - 0x23
    "00100100", --  502 - 0x1f6  :   36 - 0x24
    "00100100", --  503 - 0x1f7  :   36 - 0x24
    "00000000", --  504 - 0x1f8  :    0 - 0x0
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  529 - 0x211  :    0 - 0x0
    "11110000", --  530 - 0x212  :  240 - 0xf0
    "00001000", --  531 - 0x213  :    8 - 0x8
    "00001000", --  532 - 0x214  :    8 - 0x8
    "11110000", --  533 - 0x215  :  240 - 0xf0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00001111", --  536 - 0x218  :   15 - 0xf
    "00001111", --  537 - 0x219  :   15 - 0xf
    "00001111", --  538 - 0x21a  :   15 - 0xf
    "00000111", --  539 - 0x21b  :    7 - 0x7
    "00000111", --  540 - 0x21c  :    7 - 0x7
    "00001111", --  541 - 0x21d  :   15 - 0xf
    "00001111", --  542 - 0x21e  :   15 - 0xf
    "00001111", --  543 - 0x21f  :   15 - 0xf
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00001111", --  546 - 0x222  :   15 - 0xf
    "00010000", --  547 - 0x223  :   16 - 0x10
    "00010000", --  548 - 0x224  :   16 - 0x10
    "00001111", --  549 - 0x225  :   15 - 0xf
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "11110000", --  552 - 0x228  :  240 - 0xf0
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11110000", --  554 - 0x22a  :  240 - 0xf0
    "11100000", --  555 - 0x22b  :  224 - 0xe0
    "11100000", --  556 - 0x22c  :  224 - 0xe0
    "11110000", --  557 - 0x22d  :  240 - 0xf0
    "11110000", --  558 - 0x22e  :  240 - 0xf0
    "11110000", --  559 - 0x22f  :  240 - 0xf0
    "11111111", --  560 - 0x230  :  255 - 0xff -- Sprite 0x23
    "11111111", --  561 - 0x231  :  255 - 0xff
    "11100001", --  562 - 0x232  :  225 - 0xe1
    "11100001", --  563 - 0x233  :  225 - 0xe1
    "11100001", --  564 - 0x234  :  225 - 0xe1
    "11100001", --  565 - 0x235  :  225 - 0xe1
    "11100001", --  566 - 0x236  :  225 - 0xe1
    "11100001", --  567 - 0x237  :  225 - 0xe1
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11100001", --  570 - 0x23a  :  225 - 0xe1
    "11100001", --  571 - 0x23b  :  225 - 0xe1
    "11100001", --  572 - 0x23c  :  225 - 0xe1
    "11100001", --  573 - 0x23d  :  225 - 0xe1
    "11100001", --  574 - 0x23e  :  225 - 0xe1
    "11100001", --  575 - 0x23f  :  225 - 0xe1
    "10000111", --  576 - 0x240  :  135 - 0x87 -- Sprite 0x24
    "11000111", --  577 - 0x241  :  199 - 0xc7
    "11000000", --  578 - 0x242  :  192 - 0xc0
    "11000111", --  579 - 0x243  :  199 - 0xc7
    "11001111", --  580 - 0x244  :  207 - 0xcf
    "11001110", --  581 - 0x245  :  206 - 0xce
    "11001111", --  582 - 0x246  :  207 - 0xcf
    "11000111", --  583 - 0x247  :  199 - 0xc7
    "10000111", --  584 - 0x248  :  135 - 0x87
    "11000111", --  585 - 0x249  :  199 - 0xc7
    "11000000", --  586 - 0x24a  :  192 - 0xc0
    "11000111", --  587 - 0x24b  :  199 - 0xc7
    "11001111", --  588 - 0x24c  :  207 - 0xcf
    "11001110", --  589 - 0x24d  :  206 - 0xce
    "11001111", --  590 - 0x24e  :  207 - 0xcf
    "11000111", --  591 - 0x24f  :  199 - 0xc7
    "11111000", --  592 - 0x250  :  248 - 0xf8 -- Sprite 0x25
    "11111100", --  593 - 0x251  :  252 - 0xfc
    "00011100", --  594 - 0x252  :   28 - 0x1c
    "11111100", --  595 - 0x253  :  252 - 0xfc
    "11111100", --  596 - 0x254  :  252 - 0xfc
    "00011100", --  597 - 0x255  :   28 - 0x1c
    "11111100", --  598 - 0x256  :  252 - 0xfc
    "11111100", --  599 - 0x257  :  252 - 0xfc
    "11111000", --  600 - 0x258  :  248 - 0xf8
    "11111100", --  601 - 0x259  :  252 - 0xfc
    "00011100", --  602 - 0x25a  :   28 - 0x1c
    "11111100", --  603 - 0x25b  :  252 - 0xfc
    "11111100", --  604 - 0x25c  :  252 - 0xfc
    "00011100", --  605 - 0x25d  :   28 - 0x1c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x26
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11100111", --  610 - 0x262  :  231 - 0xe7
    "11100111", --  611 - 0x263  :  231 - 0xe7
    "11100111", --  612 - 0x264  :  231 - 0xe7
    "11100111", --  613 - 0x265  :  231 - 0xe7
    "11100111", --  614 - 0x266  :  231 - 0xe7
    "11100111", --  615 - 0x267  :  231 - 0xe7
    "11111111", --  616 - 0x268  :  255 - 0xff
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11100111", --  618 - 0x26a  :  231 - 0xe7
    "11100111", --  619 - 0x26b  :  231 - 0xe7
    "11100111", --  620 - 0x26c  :  231 - 0xe7
    "11100111", --  621 - 0x26d  :  231 - 0xe7
    "11100111", --  622 - 0x26e  :  231 - 0xe7
    "11100111", --  623 - 0x26f  :  231 - 0xe7
    "11110000", --  624 - 0x270  :  240 - 0xf0 -- Sprite 0x27
    "11111001", --  625 - 0x271  :  249 - 0xf9
    "00111001", --  626 - 0x272  :   57 - 0x39
    "00111001", --  627 - 0x273  :   57 - 0x39
    "00111001", --  628 - 0x274  :   57 - 0x39
    "00111001", --  629 - 0x275  :   57 - 0x39
    "00111001", --  630 - 0x276  :   57 - 0x39
    "00111000", --  631 - 0x277  :   56 - 0x38
    "11110000", --  632 - 0x278  :  240 - 0xf0
    "11111001", --  633 - 0x279  :  249 - 0xf9
    "00111001", --  634 - 0x27a  :   57 - 0x39
    "00111001", --  635 - 0x27b  :   57 - 0x39
    "00111001", --  636 - 0x27c  :   57 - 0x39
    "00111001", --  637 - 0x27d  :   57 - 0x39
    "00111001", --  638 - 0x27e  :   57 - 0x39
    "00111000", --  639 - 0x27f  :   56 - 0x38
    "11111111", --  640 - 0x280  :  255 - 0xff -- Sprite 0x28
    "11111111", --  641 - 0x281  :  255 - 0xff
    "11000000", --  642 - 0x282  :  192 - 0xc0
    "11000000", --  643 - 0x283  :  192 - 0xc0
    "11000000", --  644 - 0x284  :  192 - 0xc0
    "11000000", --  645 - 0x285  :  192 - 0xc0
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111111", --  648 - 0x288  :  255 - 0xff
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11000000", --  650 - 0x28a  :  192 - 0xc0
    "11000000", --  651 - 0x28b  :  192 - 0xc0
    "11000000", --  652 - 0x28c  :  192 - 0xc0
    "11000000", --  653 - 0x28d  :  192 - 0xc0
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "00011111", --  656 - 0x290  :   31 - 0x1f -- Sprite 0x29
    "00111111", --  657 - 0x291  :   63 - 0x3f
    "00110000", --  658 - 0x292  :   48 - 0x30
    "00110000", --  659 - 0x293  :   48 - 0x30
    "00110000", --  660 - 0x294  :   48 - 0x30
    "00110000", --  661 - 0x295  :   48 - 0x30
    "00111111", --  662 - 0x296  :   63 - 0x3f
    "00011111", --  663 - 0x297  :   31 - 0x1f
    "00011111", --  664 - 0x298  :   31 - 0x1f
    "00111111", --  665 - 0x299  :   63 - 0x3f
    "00110000", --  666 - 0x29a  :   48 - 0x30
    "00110000", --  667 - 0x29b  :   48 - 0x30
    "00110000", --  668 - 0x29c  :   48 - 0x30
    "00110000", --  669 - 0x29d  :   48 - 0x30
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "00011111", --  671 - 0x29f  :   31 - 0x1f
    "11100011", --  672 - 0x2a0  :  227 - 0xe3 -- Sprite 0x2a
    "11110011", --  673 - 0x2a1  :  243 - 0xf3
    "01110000", --  674 - 0x2a2  :  112 - 0x70
    "01110000", --  675 - 0x2a3  :  112 - 0x70
    "01110000", --  676 - 0x2a4  :  112 - 0x70
    "01110000", --  677 - 0x2a5  :  112 - 0x70
    "11110000", --  678 - 0x2a6  :  240 - 0xf0
    "11100000", --  679 - 0x2a7  :  224 - 0xe0
    "11100011", --  680 - 0x2a8  :  227 - 0xe3
    "11110011", --  681 - 0x2a9  :  243 - 0xf3
    "01110000", --  682 - 0x2aa  :  112 - 0x70
    "01110000", --  683 - 0x2ab  :  112 - 0x70
    "01110000", --  684 - 0x2ac  :  112 - 0x70
    "01110000", --  685 - 0x2ad  :  112 - 0x70
    "11110000", --  686 - 0x2ae  :  240 - 0xf0
    "11100000", --  687 - 0x2af  :  224 - 0xe0
    "11111110", --  688 - 0x2b0  :  254 - 0xfe -- Sprite 0x2b
    "11111110", --  689 - 0x2b1  :  254 - 0xfe
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "01110000", --  691 - 0x2b3  :  112 - 0x70
    "01110000", --  692 - 0x2b4  :  112 - 0x70
    "01110000", --  693 - 0x2b5  :  112 - 0x70
    "01110000", --  694 - 0x2b6  :  112 - 0x70
    "01110000", --  695 - 0x2b7  :  112 - 0x70
    "11111110", --  696 - 0x2b8  :  254 - 0xfe
    "11111110", --  697 - 0x2b9  :  254 - 0xfe
    "01110000", --  698 - 0x2ba  :  112 - 0x70
    "01110000", --  699 - 0x2bb  :  112 - 0x70
    "01110000", --  700 - 0x2bc  :  112 - 0x70
    "01110000", --  701 - 0x2bd  :  112 - 0x70
    "01110000", --  702 - 0x2be  :  112 - 0x70
    "01110000", --  703 - 0x2bf  :  112 - 0x70
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "11111111", --  728 - 0x2d8  :  255 - 0xff
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "11111111", --  735 - 0x2df  :  255 - 0xff
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00011000", --  739 - 0x2e3  :   24 - 0x18
    "00011000", --  740 - 0x2e4  :   24 - 0x18
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00011000", --  763 - 0x2fb  :   24 - 0x18
    "00011000", --  764 - 0x2fc  :   24 - 0x18
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00011100", --  768 - 0x300  :   28 - 0x1c -- Sprite 0x30
    "00100110", --  769 - 0x301  :   38 - 0x26
    "01100011", --  770 - 0x302  :   99 - 0x63
    "01100011", --  771 - 0x303  :   99 - 0x63
    "01100011", --  772 - 0x304  :   99 - 0x63
    "00110010", --  773 - 0x305  :   50 - 0x32
    "00011100", --  774 - 0x306  :   28 - 0x1c
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00001100", --  784 - 0x310  :   12 - 0xc -- Sprite 0x31
    "00011100", --  785 - 0x311  :   28 - 0x1c
    "00001100", --  786 - 0x312  :   12 - 0xc
    "00001100", --  787 - 0x313  :   12 - 0xc
    "00001100", --  788 - 0x314  :   12 - 0xc
    "00001100", --  789 - 0x315  :   12 - 0xc
    "00111111", --  790 - 0x316  :   63 - 0x3f
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00111110", --  800 - 0x320  :   62 - 0x3e -- Sprite 0x32
    "01100011", --  801 - 0x321  :   99 - 0x63
    "00000111", --  802 - 0x322  :    7 - 0x7
    "00011110", --  803 - 0x323  :   30 - 0x1e
    "00111100", --  804 - 0x324  :   60 - 0x3c
    "01110000", --  805 - 0x325  :  112 - 0x70
    "01111111", --  806 - 0x326  :  127 - 0x7f
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00111111", --  816 - 0x330  :   63 - 0x3f -- Sprite 0x33
    "00000110", --  817 - 0x331  :    6 - 0x6
    "00001100", --  818 - 0x332  :   12 - 0xc
    "00011110", --  819 - 0x333  :   30 - 0x1e
    "00000011", --  820 - 0x334  :    3 - 0x3
    "01100011", --  821 - 0x335  :   99 - 0x63
    "00111110", --  822 - 0x336  :   62 - 0x3e
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00001110", --  832 - 0x340  :   14 - 0xe -- Sprite 0x34
    "00011110", --  833 - 0x341  :   30 - 0x1e
    "00110110", --  834 - 0x342  :   54 - 0x36
    "01100110", --  835 - 0x343  :  102 - 0x66
    "01111111", --  836 - 0x344  :  127 - 0x7f
    "00000110", --  837 - 0x345  :    6 - 0x6
    "00000110", --  838 - 0x346  :    6 - 0x6
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "01111110", --  848 - 0x350  :  126 - 0x7e -- Sprite 0x35
    "01100000", --  849 - 0x351  :   96 - 0x60
    "01111110", --  850 - 0x352  :  126 - 0x7e
    "00000011", --  851 - 0x353  :    3 - 0x3
    "00000011", --  852 - 0x354  :    3 - 0x3
    "01100011", --  853 - 0x355  :   99 - 0x63
    "00111110", --  854 - 0x356  :   62 - 0x3e
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00011110", --  864 - 0x360  :   30 - 0x1e -- Sprite 0x36
    "00110000", --  865 - 0x361  :   48 - 0x30
    "01100000", --  866 - 0x362  :   96 - 0x60
    "01111110", --  867 - 0x363  :  126 - 0x7e
    "01100011", --  868 - 0x364  :   99 - 0x63
    "01100011", --  869 - 0x365  :   99 - 0x63
    "00111110", --  870 - 0x366  :   62 - 0x3e
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "01111111", --  880 - 0x370  :  127 - 0x7f -- Sprite 0x37
    "01100011", --  881 - 0x371  :   99 - 0x63
    "00000110", --  882 - 0x372  :    6 - 0x6
    "00001100", --  883 - 0x373  :   12 - 0xc
    "00011000", --  884 - 0x374  :   24 - 0x18
    "00011000", --  885 - 0x375  :   24 - 0x18
    "00011000", --  886 - 0x376  :   24 - 0x18
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00111100", --  896 - 0x380  :   60 - 0x3c -- Sprite 0x38
    "01100010", --  897 - 0x381  :   98 - 0x62
    "01110010", --  898 - 0x382  :  114 - 0x72
    "00111100", --  899 - 0x383  :   60 - 0x3c
    "01001111", --  900 - 0x384  :   79 - 0x4f
    "01000011", --  901 - 0x385  :   67 - 0x43
    "00111110", --  902 - 0x386  :   62 - 0x3e
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00111110", --  912 - 0x390  :   62 - 0x3e -- Sprite 0x39
    "01100011", --  913 - 0x391  :   99 - 0x63
    "01100011", --  914 - 0x392  :   99 - 0x63
    "00111111", --  915 - 0x393  :   63 - 0x3f
    "00000011", --  916 - 0x394  :    3 - 0x3
    "00000110", --  917 - 0x395  :    6 - 0x6
    "00111100", --  918 - 0x396  :   60 - 0x3c
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "01111110", --  931 - 0x3a3  :  126 - 0x7e
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x3b
    "00000010", --  945 - 0x3b1  :    2 - 0x2
    "00000100", --  946 - 0x3b2  :    4 - 0x4
    "00001000", --  947 - 0x3b3  :    8 - 0x8
    "00010000", --  948 - 0x3b4  :   16 - 0x10
    "00100000", --  949 - 0x3b5  :   32 - 0x20
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000111", --  961 - 0x3c1  :    7 - 0x7
    "00011111", --  962 - 0x3c2  :   31 - 0x1f
    "00111111", --  963 - 0x3c3  :   63 - 0x3f
    "00111111", --  964 - 0x3c4  :   63 - 0x3f
    "00001111", --  965 - 0x3c5  :   15 - 0xf
    "00000011", --  966 - 0x3c6  :    3 - 0x3
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000111", --  969 - 0x3c9  :    7 - 0x7
    "00011111", --  970 - 0x3ca  :   31 - 0x1f
    "00111111", --  971 - 0x3cb  :   63 - 0x3f
    "00111111", --  972 - 0x3cc  :   63 - 0x3f
    "00001111", --  973 - 0x3cd  :   15 - 0xf
    "00000011", --  974 - 0x3ce  :    3 - 0x3
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x3d
    "11000000", --  977 - 0x3d1  :  192 - 0xc0
    "11110000", --  978 - 0x3d2  :  240 - 0xf0
    "11111000", --  979 - 0x3d3  :  248 - 0xf8
    "11111000", --  980 - 0x3d4  :  248 - 0xf8
    "11111100", --  981 - 0x3d5  :  252 - 0xfc
    "11111100", --  982 - 0x3d6  :  252 - 0xfc
    "11111100", --  983 - 0x3d7  :  252 - 0xfc
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "11000000", --  985 - 0x3d9  :  192 - 0xc0
    "11110000", --  986 - 0x3da  :  240 - 0xf0
    "11111000", --  987 - 0x3db  :  248 - 0xf8
    "11111000", --  988 - 0x3dc  :  248 - 0xf8
    "11111100", --  989 - 0x3dd  :  252 - 0xfc
    "11111100", --  990 - 0x3de  :  252 - 0xfc
    "11111100", --  991 - 0x3df  :  252 - 0xfc
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000011", --  993 - 0x3e1  :    3 - 0x3
    "00001111", --  994 - 0x3e2  :   15 - 0xf
    "00111111", --  995 - 0x3e3  :   63 - 0x3f
    "00111111", --  996 - 0x3e4  :   63 - 0x3f
    "00011111", --  997 - 0x3e5  :   31 - 0x1f
    "00000111", --  998 - 0x3e6  :    7 - 0x7
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000011", -- 1001 - 0x3e9  :    3 - 0x3
    "00001111", -- 1002 - 0x3ea  :   15 - 0xf
    "00111111", -- 1003 - 0x3eb  :   63 - 0x3f
    "00111111", -- 1004 - 0x3ec  :   63 - 0x3f
    "00011111", -- 1005 - 0x3ed  :   31 - 0x1f
    "00000111", -- 1006 - 0x3ee  :    7 - 0x7
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "11111100", -- 1008 - 0x3f0  :  252 - 0xfc -- Sprite 0x3f
    "11111100", -- 1009 - 0x3f1  :  252 - 0xfc
    "11111100", -- 1010 - 0x3f2  :  252 - 0xfc
    "11111000", -- 1011 - 0x3f3  :  248 - 0xf8
    "11111000", -- 1012 - 0x3f4  :  248 - 0xf8
    "11110000", -- 1013 - 0x3f5  :  240 - 0xf0
    "11000000", -- 1014 - 0x3f6  :  192 - 0xc0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "11111100", -- 1016 - 0x3f8  :  252 - 0xfc
    "11111100", -- 1017 - 0x3f9  :  252 - 0xfc
    "11111100", -- 1018 - 0x3fa  :  252 - 0xfc
    "11111000", -- 1019 - 0x3fb  :  248 - 0xf8
    "11111000", -- 1020 - 0x3fc  :  248 - 0xf8
    "11110000", -- 1021 - 0x3fd  :  240 - 0xf0
    "11000000", -- 1022 - 0x3fe  :  192 - 0xc0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Sprite 0x40
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00011100", -- 1040 - 0x410  :   28 - 0x1c -- Sprite 0x41
    "00110110", -- 1041 - 0x411  :   54 - 0x36
    "01100011", -- 1042 - 0x412  :   99 - 0x63
    "01100011", -- 1043 - 0x413  :   99 - 0x63
    "01111111", -- 1044 - 0x414  :  127 - 0x7f
    "01100011", -- 1045 - 0x415  :   99 - 0x63
    "01100011", -- 1046 - 0x416  :   99 - 0x63
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "01111110", -- 1056 - 0x420  :  126 - 0x7e -- Sprite 0x42
    "01100011", -- 1057 - 0x421  :   99 - 0x63
    "01100011", -- 1058 - 0x422  :   99 - 0x63
    "01111110", -- 1059 - 0x423  :  126 - 0x7e
    "01100011", -- 1060 - 0x424  :   99 - 0x63
    "01100011", -- 1061 - 0x425  :   99 - 0x63
    "01111110", -- 1062 - 0x426  :  126 - 0x7e
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00011110", -- 1072 - 0x430  :   30 - 0x1e -- Sprite 0x43
    "00110011", -- 1073 - 0x431  :   51 - 0x33
    "01100000", -- 1074 - 0x432  :   96 - 0x60
    "01100000", -- 1075 - 0x433  :   96 - 0x60
    "01100000", -- 1076 - 0x434  :   96 - 0x60
    "00110011", -- 1077 - 0x435  :   51 - 0x33
    "00011110", -- 1078 - 0x436  :   30 - 0x1e
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "01111100", -- 1088 - 0x440  :  124 - 0x7c -- Sprite 0x44
    "01100110", -- 1089 - 0x441  :  102 - 0x66
    "01100011", -- 1090 - 0x442  :   99 - 0x63
    "01100011", -- 1091 - 0x443  :   99 - 0x63
    "01100011", -- 1092 - 0x444  :   99 - 0x63
    "01100110", -- 1093 - 0x445  :  102 - 0x66
    "01111100", -- 1094 - 0x446  :  124 - 0x7c
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "01111111", -- 1104 - 0x450  :  127 - 0x7f -- Sprite 0x45
    "01100000", -- 1105 - 0x451  :   96 - 0x60
    "01100000", -- 1106 - 0x452  :   96 - 0x60
    "01111110", -- 1107 - 0x453  :  126 - 0x7e
    "01100000", -- 1108 - 0x454  :   96 - 0x60
    "01100000", -- 1109 - 0x455  :   96 - 0x60
    "01111111", -- 1110 - 0x456  :  127 - 0x7f
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "01111111", -- 1120 - 0x460  :  127 - 0x7f -- Sprite 0x46
    "01100000", -- 1121 - 0x461  :   96 - 0x60
    "01100000", -- 1122 - 0x462  :   96 - 0x60
    "01111110", -- 1123 - 0x463  :  126 - 0x7e
    "01100000", -- 1124 - 0x464  :   96 - 0x60
    "01100000", -- 1125 - 0x465  :   96 - 0x60
    "01100000", -- 1126 - 0x466  :   96 - 0x60
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00011111", -- 1136 - 0x470  :   31 - 0x1f -- Sprite 0x47
    "00110000", -- 1137 - 0x471  :   48 - 0x30
    "01100000", -- 1138 - 0x472  :   96 - 0x60
    "01100111", -- 1139 - 0x473  :  103 - 0x67
    "01100011", -- 1140 - 0x474  :   99 - 0x63
    "00110011", -- 1141 - 0x475  :   51 - 0x33
    "00011111", -- 1142 - 0x476  :   31 - 0x1f
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "01100011", -- 1152 - 0x480  :   99 - 0x63 -- Sprite 0x48
    "01100011", -- 1153 - 0x481  :   99 - 0x63
    "01100011", -- 1154 - 0x482  :   99 - 0x63
    "01111111", -- 1155 - 0x483  :  127 - 0x7f
    "01100011", -- 1156 - 0x484  :   99 - 0x63
    "01100011", -- 1157 - 0x485  :   99 - 0x63
    "01100011", -- 1158 - 0x486  :   99 - 0x63
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00111111", -- 1168 - 0x490  :   63 - 0x3f -- Sprite 0x49
    "00001100", -- 1169 - 0x491  :   12 - 0xc
    "00001100", -- 1170 - 0x492  :   12 - 0xc
    "00001100", -- 1171 - 0x493  :   12 - 0xc
    "00001100", -- 1172 - 0x494  :   12 - 0xc
    "00001100", -- 1173 - 0x495  :   12 - 0xc
    "00111111", -- 1174 - 0x496  :   63 - 0x3f
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000011", -- 1184 - 0x4a0  :    3 - 0x3 -- Sprite 0x4a
    "00000011", -- 1185 - 0x4a1  :    3 - 0x3
    "00000011", -- 1186 - 0x4a2  :    3 - 0x3
    "00000011", -- 1187 - 0x4a3  :    3 - 0x3
    "00000011", -- 1188 - 0x4a4  :    3 - 0x3
    "01100011", -- 1189 - 0x4a5  :   99 - 0x63
    "00111110", -- 1190 - 0x4a6  :   62 - 0x3e
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "01100011", -- 1200 - 0x4b0  :   99 - 0x63 -- Sprite 0x4b
    "01100110", -- 1201 - 0x4b1  :  102 - 0x66
    "01101100", -- 1202 - 0x4b2  :  108 - 0x6c
    "01111000", -- 1203 - 0x4b3  :  120 - 0x78
    "01111100", -- 1204 - 0x4b4  :  124 - 0x7c
    "01100110", -- 1205 - 0x4b5  :  102 - 0x66
    "01100011", -- 1206 - 0x4b6  :   99 - 0x63
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "01100000", -- 1216 - 0x4c0  :   96 - 0x60 -- Sprite 0x4c
    "01100000", -- 1217 - 0x4c1  :   96 - 0x60
    "01100000", -- 1218 - 0x4c2  :   96 - 0x60
    "01100000", -- 1219 - 0x4c3  :   96 - 0x60
    "01100000", -- 1220 - 0x4c4  :   96 - 0x60
    "01100000", -- 1221 - 0x4c5  :   96 - 0x60
    "01111111", -- 1222 - 0x4c6  :  127 - 0x7f
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "01100011", -- 1232 - 0x4d0  :   99 - 0x63 -- Sprite 0x4d
    "01110111", -- 1233 - 0x4d1  :  119 - 0x77
    "01111111", -- 1234 - 0x4d2  :  127 - 0x7f
    "01111111", -- 1235 - 0x4d3  :  127 - 0x7f
    "01101011", -- 1236 - 0x4d4  :  107 - 0x6b
    "01100011", -- 1237 - 0x4d5  :   99 - 0x63
    "01100011", -- 1238 - 0x4d6  :   99 - 0x63
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "01100011", -- 1248 - 0x4e0  :   99 - 0x63 -- Sprite 0x4e
    "01110011", -- 1249 - 0x4e1  :  115 - 0x73
    "01111011", -- 1250 - 0x4e2  :  123 - 0x7b
    "01111111", -- 1251 - 0x4e3  :  127 - 0x7f
    "01101111", -- 1252 - 0x4e4  :  111 - 0x6f
    "01100111", -- 1253 - 0x4e5  :  103 - 0x67
    "01100011", -- 1254 - 0x4e6  :   99 - 0x63
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00111110", -- 1264 - 0x4f0  :   62 - 0x3e -- Sprite 0x4f
    "01100011", -- 1265 - 0x4f1  :   99 - 0x63
    "01100011", -- 1266 - 0x4f2  :   99 - 0x63
    "01100011", -- 1267 - 0x4f3  :   99 - 0x63
    "01100011", -- 1268 - 0x4f4  :   99 - 0x63
    "01100011", -- 1269 - 0x4f5  :   99 - 0x63
    "00111110", -- 1270 - 0x4f6  :   62 - 0x3e
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "01111110", -- 1280 - 0x500  :  126 - 0x7e -- Sprite 0x50
    "01100011", -- 1281 - 0x501  :   99 - 0x63
    "01100011", -- 1282 - 0x502  :   99 - 0x63
    "01100011", -- 1283 - 0x503  :   99 - 0x63
    "01111110", -- 1284 - 0x504  :  126 - 0x7e
    "01100000", -- 1285 - 0x505  :   96 - 0x60
    "01100000", -- 1286 - 0x506  :   96 - 0x60
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00111110", -- 1296 - 0x510  :   62 - 0x3e -- Sprite 0x51
    "01100011", -- 1297 - 0x511  :   99 - 0x63
    "01100011", -- 1298 - 0x512  :   99 - 0x63
    "01100011", -- 1299 - 0x513  :   99 - 0x63
    "01101111", -- 1300 - 0x514  :  111 - 0x6f
    "01100110", -- 1301 - 0x515  :  102 - 0x66
    "00111101", -- 1302 - 0x516  :   61 - 0x3d
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "01111110", -- 1312 - 0x520  :  126 - 0x7e -- Sprite 0x52
    "01100011", -- 1313 - 0x521  :   99 - 0x63
    "01100011", -- 1314 - 0x522  :   99 - 0x63
    "01100111", -- 1315 - 0x523  :  103 - 0x67
    "01111100", -- 1316 - 0x524  :  124 - 0x7c
    "01101110", -- 1317 - 0x525  :  110 - 0x6e
    "01100111", -- 1318 - 0x526  :  103 - 0x67
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00111100", -- 1328 - 0x530  :   60 - 0x3c -- Sprite 0x53
    "01100110", -- 1329 - 0x531  :  102 - 0x66
    "01100000", -- 1330 - 0x532  :   96 - 0x60
    "00111110", -- 1331 - 0x533  :   62 - 0x3e
    "00000011", -- 1332 - 0x534  :    3 - 0x3
    "01100011", -- 1333 - 0x535  :   99 - 0x63
    "00111110", -- 1334 - 0x536  :   62 - 0x3e
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00111111", -- 1344 - 0x540  :   63 - 0x3f -- Sprite 0x54
    "00001100", -- 1345 - 0x541  :   12 - 0xc
    "00001100", -- 1346 - 0x542  :   12 - 0xc
    "00001100", -- 1347 - 0x543  :   12 - 0xc
    "00001100", -- 1348 - 0x544  :   12 - 0xc
    "00001100", -- 1349 - 0x545  :   12 - 0xc
    "00001100", -- 1350 - 0x546  :   12 - 0xc
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "01100011", -- 1360 - 0x550  :   99 - 0x63 -- Sprite 0x55
    "01100011", -- 1361 - 0x551  :   99 - 0x63
    "01100011", -- 1362 - 0x552  :   99 - 0x63
    "01100011", -- 1363 - 0x553  :   99 - 0x63
    "01100011", -- 1364 - 0x554  :   99 - 0x63
    "01100011", -- 1365 - 0x555  :   99 - 0x63
    "00111110", -- 1366 - 0x556  :   62 - 0x3e
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "01100011", -- 1376 - 0x560  :   99 - 0x63 -- Sprite 0x56
    "01100011", -- 1377 - 0x561  :   99 - 0x63
    "01100011", -- 1378 - 0x562  :   99 - 0x63
    "01110111", -- 1379 - 0x563  :  119 - 0x77
    "00111110", -- 1380 - 0x564  :   62 - 0x3e
    "00011100", -- 1381 - 0x565  :   28 - 0x1c
    "00001000", -- 1382 - 0x566  :    8 - 0x8
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "01100011", -- 1392 - 0x570  :   99 - 0x63 -- Sprite 0x57
    "01100011", -- 1393 - 0x571  :   99 - 0x63
    "01101011", -- 1394 - 0x572  :  107 - 0x6b
    "01111111", -- 1395 - 0x573  :  127 - 0x7f
    "01111111", -- 1396 - 0x574  :  127 - 0x7f
    "01110111", -- 1397 - 0x575  :  119 - 0x77
    "01100011", -- 1398 - 0x576  :   99 - 0x63
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "01100011", -- 1408 - 0x580  :   99 - 0x63 -- Sprite 0x58
    "01110111", -- 1409 - 0x581  :  119 - 0x77
    "00111110", -- 1410 - 0x582  :   62 - 0x3e
    "00011100", -- 1411 - 0x583  :   28 - 0x1c
    "00111110", -- 1412 - 0x584  :   62 - 0x3e
    "01110111", -- 1413 - 0x585  :  119 - 0x77
    "01100011", -- 1414 - 0x586  :   99 - 0x63
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00110011", -- 1424 - 0x590  :   51 - 0x33 -- Sprite 0x59
    "00110011", -- 1425 - 0x591  :   51 - 0x33
    "00110011", -- 1426 - 0x592  :   51 - 0x33
    "00011110", -- 1427 - 0x593  :   30 - 0x1e
    "00001100", -- 1428 - 0x594  :   12 - 0xc
    "00001100", -- 1429 - 0x595  :   12 - 0xc
    "00001100", -- 1430 - 0x596  :   12 - 0xc
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01111111", -- 1440 - 0x5a0  :  127 - 0x7f -- Sprite 0x5a
    "00000111", -- 1441 - 0x5a1  :    7 - 0x7
    "00001110", -- 1442 - 0x5a2  :   14 - 0xe
    "00011100", -- 1443 - 0x5a3  :   28 - 0x1c
    "00111000", -- 1444 - 0x5a4  :   56 - 0x38
    "01110000", -- 1445 - 0x5a5  :  112 - 0x70
    "01111111", -- 1446 - 0x5a6  :  127 - 0x7f
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00110000", -- 1461 - 0x5b5  :   48 - 0x30
    "00110000", -- 1462 - 0x5b6  :   48 - 0x30
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0 -- Sprite 0x5c
    "11110000", -- 1473 - 0x5c1  :  240 - 0xf0
    "11111100", -- 1474 - 0x5c2  :  252 - 0xfc
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111100", -- 1476 - 0x5c4  :  252 - 0xfc
    "11110000", -- 1477 - 0x5c5  :  240 - 0xf0
    "11000000", -- 1478 - 0x5c6  :  192 - 0xc0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00111100", -- 1488 - 0x5d0  :   60 - 0x3c -- Sprite 0x5d
    "01000010", -- 1489 - 0x5d1  :   66 - 0x42
    "10011001", -- 1490 - 0x5d2  :  153 - 0x99
    "10100001", -- 1491 - 0x5d3  :  161 - 0xa1
    "10100001", -- 1492 - 0x5d4  :  161 - 0xa1
    "10011001", -- 1493 - 0x5d5  :  153 - 0x99
    "01000010", -- 1494 - 0x5d6  :   66 - 0x42
    "00111100", -- 1495 - 0x5d7  :   60 - 0x3c
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00010000", -- 1506 - 0x5e2  :   16 - 0x10
    "00010000", -- 1507 - 0x5e3  :   16 - 0x10
    "00010000", -- 1508 - 0x5e4  :   16 - 0x10
    "00010000", -- 1509 - 0x5e5  :   16 - 0x10
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00010000", -- 1514 - 0x5ea  :   16 - 0x10
    "00010000", -- 1515 - 0x5eb  :   16 - 0x10
    "00010000", -- 1516 - 0x5ec  :   16 - 0x10
    "00010000", -- 1517 - 0x5ed  :   16 - 0x10
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00110110", -- 1520 - 0x5f0  :   54 - 0x36 -- Sprite 0x5f
    "00110110", -- 1521 - 0x5f1  :   54 - 0x36
    "00010010", -- 1522 - 0x5f2  :   18 - 0x12
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000001", -- 1541 - 0x605  :    1 - 0x1
    "00011110", -- 1542 - 0x606  :   30 - 0x1e
    "00111011", -- 1543 - 0x607  :   59 - 0x3b
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0x61
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00001100", -- 1554 - 0x612  :   12 - 0xc
    "00111100", -- 1555 - 0x613  :   60 - 0x3c
    "11010000", -- 1556 - 0x614  :  208 - 0xd0
    "00010000", -- 1557 - 0x615  :   16 - 0x10
    "00100000", -- 1558 - 0x616  :   32 - 0x20
    "01000000", -- 1559 - 0x617  :   64 - 0x40
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00111110", -- 1568 - 0x620  :   62 - 0x3e -- Sprite 0x62
    "00101101", -- 1569 - 0x621  :   45 - 0x2d
    "00110101", -- 1570 - 0x622  :   53 - 0x35
    "00011101", -- 1571 - 0x623  :   29 - 0x1d
    "00000001", -- 1572 - 0x624  :    1 - 0x1
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "10110000", -- 1584 - 0x630  :  176 - 0xb0 -- Sprite 0x63
    "10111000", -- 1585 - 0x631  :  184 - 0xb8
    "11111000", -- 1586 - 0x632  :  248 - 0xf8
    "01111000", -- 1587 - 0x633  :  120 - 0x78
    "10011000", -- 1588 - 0x634  :  152 - 0x98
    "11110000", -- 1589 - 0x635  :  240 - 0xf0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000111", -- 1602 - 0x642  :    7 - 0x7
    "00000011", -- 1603 - 0x643  :    3 - 0x3
    "00001101", -- 1604 - 0x644  :   13 - 0xd
    "00011110", -- 1605 - 0x645  :   30 - 0x1e
    "00010111", -- 1606 - 0x646  :   23 - 0x17
    "00011101", -- 1607 - 0x647  :   29 - 0x1d
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "10000000", -- 1617 - 0x651  :  128 - 0x80
    "01110000", -- 1618 - 0x652  :  112 - 0x70
    "11100000", -- 1619 - 0x653  :  224 - 0xe0
    "11011000", -- 1620 - 0x654  :  216 - 0xd8
    "10111100", -- 1621 - 0x655  :  188 - 0xbc
    "01110100", -- 1622 - 0x656  :  116 - 0x74
    "11011100", -- 1623 - 0x657  :  220 - 0xdc
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00011111", -- 1632 - 0x660  :   31 - 0x1f -- Sprite 0x66
    "00001011", -- 1633 - 0x661  :   11 - 0xb
    "00001111", -- 1634 - 0x662  :   15 - 0xf
    "00000101", -- 1635 - 0x663  :    5 - 0x5
    "00000011", -- 1636 - 0x664  :    3 - 0x3
    "00000001", -- 1637 - 0x665  :    1 - 0x1
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11111100", -- 1648 - 0x670  :  252 - 0xfc -- Sprite 0x67
    "01101000", -- 1649 - 0x671  :  104 - 0x68
    "11111000", -- 1650 - 0x672  :  248 - 0xf8
    "10110000", -- 1651 - 0x673  :  176 - 0xb0
    "11100000", -- 1652 - 0x674  :  224 - 0xe0
    "10000000", -- 1653 - 0x675  :  128 - 0x80
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000001", -- 1675 - 0x68b  :    1 - 0x1
    "00000001", -- 1676 - 0x68c  :    1 - 0x1
    "00001011", -- 1677 - 0x68d  :   11 - 0xb
    "00011100", -- 1678 - 0x68e  :   28 - 0x1c
    "00111111", -- 1679 - 0x68f  :   63 - 0x3f
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00110000", -- 1690 - 0x69a  :   48 - 0x30
    "01111000", -- 1691 - 0x69b  :  120 - 0x78
    "10000000", -- 1692 - 0x69c  :  128 - 0x80
    "11110000", -- 1693 - 0x69d  :  240 - 0xf0
    "11111000", -- 1694 - 0x69e  :  248 - 0xf8
    "11111100", -- 1695 - 0x69f  :  252 - 0xfc
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00111111", -- 1704 - 0x6a8  :   63 - 0x3f
    "00111111", -- 1705 - 0x6a9  :   63 - 0x3f
    "00111111", -- 1706 - 0x6aa  :   63 - 0x3f
    "00011111", -- 1707 - 0x6ab  :   31 - 0x1f
    "00011111", -- 1708 - 0x6ac  :   31 - 0x1f
    "00000111", -- 1709 - 0x6ad  :    7 - 0x7
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0x6b
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "11111100", -- 1720 - 0x6b8  :  252 - 0xfc
    "11101100", -- 1721 - 0x6b9  :  236 - 0xec
    "11101100", -- 1722 - 0x6ba  :  236 - 0xec
    "11011000", -- 1723 - 0x6bb  :  216 - 0xd8
    "11111000", -- 1724 - 0x6bc  :  248 - 0xf8
    "11100000", -- 1725 - 0x6bd  :  224 - 0xe0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0x6c
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000001", -- 1730 - 0x6c2  :    1 - 0x1
    "00011101", -- 1731 - 0x6c3  :   29 - 0x1d
    "00111110", -- 1732 - 0x6c4  :   62 - 0x3e
    "00111111", -- 1733 - 0x6c5  :   63 - 0x3f
    "00111111", -- 1734 - 0x6c6  :   63 - 0x3f
    "00111111", -- 1735 - 0x6c7  :   63 - 0x3f
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000001", -- 1738 - 0x6ca  :    1 - 0x1
    "00011101", -- 1739 - 0x6cb  :   29 - 0x1d
    "00111110", -- 1740 - 0x6cc  :   62 - 0x3e
    "00111111", -- 1741 - 0x6cd  :   63 - 0x3f
    "00111111", -- 1742 - 0x6ce  :   63 - 0x3f
    "00111111", -- 1743 - 0x6cf  :   63 - 0x3f
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0x6d
    "10000000", -- 1745 - 0x6d1  :  128 - 0x80
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "01110000", -- 1747 - 0x6d3  :  112 - 0x70
    "11111000", -- 1748 - 0x6d4  :  248 - 0xf8
    "11111100", -- 1749 - 0x6d5  :  252 - 0xfc
    "11111100", -- 1750 - 0x6d6  :  252 - 0xfc
    "11111100", -- 1751 - 0x6d7  :  252 - 0xfc
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "01110000", -- 1755 - 0x6db  :  112 - 0x70
    "11111000", -- 1756 - 0x6dc  :  248 - 0xf8
    "11111100", -- 1757 - 0x6dd  :  252 - 0xfc
    "11111100", -- 1758 - 0x6de  :  252 - 0xfc
    "11111100", -- 1759 - 0x6df  :  252 - 0xfc
    "00111111", -- 1760 - 0x6e0  :   63 - 0x3f -- Sprite 0x6e
    "00111111", -- 1761 - 0x6e1  :   63 - 0x3f
    "00011111", -- 1762 - 0x6e2  :   31 - 0x1f
    "00011111", -- 1763 - 0x6e3  :   31 - 0x1f
    "00001111", -- 1764 - 0x6e4  :   15 - 0xf
    "00000110", -- 1765 - 0x6e5  :    6 - 0x6
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00111111", -- 1768 - 0x6e8  :   63 - 0x3f
    "00111111", -- 1769 - 0x6e9  :   63 - 0x3f
    "00011111", -- 1770 - 0x6ea  :   31 - 0x1f
    "00011111", -- 1771 - 0x6eb  :   31 - 0x1f
    "00001111", -- 1772 - 0x6ec  :   15 - 0xf
    "00000110", -- 1773 - 0x6ed  :    6 - 0x6
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11101100", -- 1776 - 0x6f0  :  236 - 0xec -- Sprite 0x6f
    "11101100", -- 1777 - 0x6f1  :  236 - 0xec
    "11011000", -- 1778 - 0x6f2  :  216 - 0xd8
    "11111000", -- 1779 - 0x6f3  :  248 - 0xf8
    "11110000", -- 1780 - 0x6f4  :  240 - 0xf0
    "11100000", -- 1781 - 0x6f5  :  224 - 0xe0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "11101100", -- 1784 - 0x6f8  :  236 - 0xec
    "11101100", -- 1785 - 0x6f9  :  236 - 0xec
    "11011000", -- 1786 - 0x6fa  :  216 - 0xd8
    "11111000", -- 1787 - 0x6fb  :  248 - 0xf8
    "11110000", -- 1788 - 0x6fc  :  240 - 0xf0
    "11100000", -- 1789 - 0x6fd  :  224 - 0xe0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0x70
    "00000100", -- 1793 - 0x701  :    4 - 0x4
    "00000011", -- 1794 - 0x702  :    3 - 0x3
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000001", -- 1796 - 0x704  :    1 - 0x1
    "00000111", -- 1797 - 0x705  :    7 - 0x7
    "00001111", -- 1798 - 0x706  :   15 - 0xf
    "00001100", -- 1799 - 0x707  :   12 - 0xc
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0x71
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "11100000", -- 1810 - 0x712  :  224 - 0xe0
    "10000000", -- 1811 - 0x713  :  128 - 0x80
    "01000000", -- 1812 - 0x714  :   64 - 0x40
    "11110000", -- 1813 - 0x715  :  240 - 0xf0
    "10011000", -- 1814 - 0x716  :  152 - 0x98
    "11111000", -- 1815 - 0x717  :  248 - 0xf8
    "00000000", -- 1816 - 0x718  :    0 - 0x0
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00011111", -- 1824 - 0x720  :   31 - 0x1f -- Sprite 0x72
    "00010011", -- 1825 - 0x721  :   19 - 0x13
    "00011111", -- 1826 - 0x722  :   31 - 0x1f
    "00001111", -- 1827 - 0x723  :   15 - 0xf
    "00001001", -- 1828 - 0x724  :    9 - 0x9
    "00000111", -- 1829 - 0x725  :    7 - 0x7
    "00000001", -- 1830 - 0x726  :    1 - 0x1
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "11100100", -- 1840 - 0x730  :  228 - 0xe4 -- Sprite 0x73
    "00111100", -- 1841 - 0x731  :   60 - 0x3c
    "11100100", -- 1842 - 0x732  :  228 - 0xe4
    "00111000", -- 1843 - 0x733  :   56 - 0x38
    "11111000", -- 1844 - 0x734  :  248 - 0xf8
    "11110000", -- 1845 - 0x735  :  240 - 0xf0
    "11000000", -- 1846 - 0x736  :  192 - 0xc0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0x74
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00010001", -- 1868 - 0x74c  :   17 - 0x11
    "00010011", -- 1869 - 0x74d  :   19 - 0x13
    "00011111", -- 1870 - 0x74e  :   31 - 0x1f
    "00011111", -- 1871 - 0x74f  :   31 - 0x1f
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0x75
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "10000000", -- 1883 - 0x75b  :  128 - 0x80
    "11000100", -- 1884 - 0x75c  :  196 - 0xc4
    "11100100", -- 1885 - 0x75d  :  228 - 0xe4
    "11111100", -- 1886 - 0x75e  :  252 - 0xfc
    "11111100", -- 1887 - 0x75f  :  252 - 0xfc
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0x76
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00011111", -- 1896 - 0x768  :   31 - 0x1f
    "00001110", -- 1897 - 0x769  :   14 - 0xe
    "00000110", -- 1898 - 0x76a  :    6 - 0x6
    "00000010", -- 1899 - 0x76b  :    2 - 0x2
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0x77
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "11111100", -- 1912 - 0x778  :  252 - 0xfc
    "10111000", -- 1913 - 0x779  :  184 - 0xb8
    "10110000", -- 1914 - 0x77a  :  176 - 0xb0
    "10100000", -- 1915 - 0x77b  :  160 - 0xa0
    "10000000", -- 1916 - 0x77c  :  128 - 0x80
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000001", -- 1931 - 0x78b  :    1 - 0x1
    "00000011", -- 1932 - 0x78c  :    3 - 0x3
    "00000110", -- 1933 - 0x78d  :    6 - 0x6
    "00000110", -- 1934 - 0x78e  :    6 - 0x6
    "00001111", -- 1935 - 0x78f  :   15 - 0xf
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0x79
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0
    "00011000", -- 1945 - 0x799  :   24 - 0x18
    "11110100", -- 1946 - 0x79a  :  244 - 0xf4
    "11111000", -- 1947 - 0x79b  :  248 - 0xf8
    "00111000", -- 1948 - 0x79c  :   56 - 0x38
    "01111100", -- 1949 - 0x79d  :  124 - 0x7c
    "11111100", -- 1950 - 0x79e  :  252 - 0xfc
    "11111100", -- 1951 - 0x79f  :  252 - 0xfc
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00001111", -- 1960 - 0x7a8  :   15 - 0xf
    "00011111", -- 1961 - 0x7a9  :   31 - 0x1f
    "00110000", -- 1962 - 0x7aa  :   48 - 0x30
    "00111000", -- 1963 - 0x7ab  :   56 - 0x38
    "00011101", -- 1964 - 0x7ac  :   29 - 0x1d
    "00000011", -- 1965 - 0x7ad  :    3 - 0x3
    "00000011", -- 1966 - 0x7ae  :    3 - 0x3
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0x7b
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "11111100", -- 1976 - 0x7b8  :  252 - 0xfc
    "11111100", -- 1977 - 0x7b9  :  252 - 0xfc
    "01111100", -- 1978 - 0x7ba  :  124 - 0x7c
    "10001110", -- 1979 - 0x7bb  :  142 - 0x8e
    "10000110", -- 1980 - 0x7bc  :  134 - 0x86
    "10011100", -- 1981 - 0x7bd  :  156 - 0x9c
    "01111000", -- 1982 - 0x7be  :  120 - 0x78
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0x7c
    "00000001", -- 1985 - 0x7c1  :    1 - 0x1
    "00000110", -- 1986 - 0x7c2  :    6 - 0x6
    "00000111", -- 1987 - 0x7c3  :    7 - 0x7
    "00000111", -- 1988 - 0x7c4  :    7 - 0x7
    "00000111", -- 1989 - 0x7c5  :    7 - 0x7
    "00000001", -- 1990 - 0x7c6  :    1 - 0x1
    "00000011", -- 1991 - 0x7c7  :    3 - 0x3
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000001", -- 1993 - 0x7c9  :    1 - 0x1
    "00000110", -- 1994 - 0x7ca  :    6 - 0x6
    "00000111", -- 1995 - 0x7cb  :    7 - 0x7
    "00000111", -- 1996 - 0x7cc  :    7 - 0x7
    "00000111", -- 1997 - 0x7cd  :    7 - 0x7
    "00000001", -- 1998 - 0x7ce  :    1 - 0x1
    "00000011", -- 1999 - 0x7cf  :    3 - 0x3
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0x7d
    "11000000", -- 2001 - 0x7d1  :  192 - 0xc0
    "00110000", -- 2002 - 0x7d2  :   48 - 0x30
    "11110000", -- 2003 - 0x7d3  :  240 - 0xf0
    "11110000", -- 2004 - 0x7d4  :  240 - 0xf0
    "11110000", -- 2005 - 0x7d5  :  240 - 0xf0
    "01000000", -- 2006 - 0x7d6  :   64 - 0x40
    "01000000", -- 2007 - 0x7d7  :   64 - 0x40
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "11000000", -- 2009 - 0x7d9  :  192 - 0xc0
    "00110000", -- 2010 - 0x7da  :   48 - 0x30
    "11110000", -- 2011 - 0x7db  :  240 - 0xf0
    "11110000", -- 2012 - 0x7dc  :  240 - 0xf0
    "11110000", -- 2013 - 0x7dd  :  240 - 0xf0
    "01000000", -- 2014 - 0x7de  :   64 - 0x40
    "01000000", -- 2015 - 0x7df  :   64 - 0x40
    "00000001", -- 2016 - 0x7e0  :    1 - 0x1 -- Sprite 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000001", -- 2018 - 0x7e2  :    1 - 0x1
    "00000011", -- 2019 - 0x7e3  :    3 - 0x3
    "00000001", -- 2020 - 0x7e4  :    1 - 0x1
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000001", -- 2024 - 0x7e8  :    1 - 0x1
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000001", -- 2026 - 0x7ea  :    1 - 0x1
    "00000011", -- 2027 - 0x7eb  :    3 - 0x3
    "00000001", -- 2028 - 0x7ec  :    1 - 0x1
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "01000000", -- 2032 - 0x7f0  :   64 - 0x40 -- Sprite 0x7f
    "01000000", -- 2033 - 0x7f1  :   64 - 0x40
    "01000000", -- 2034 - 0x7f2  :   64 - 0x40
    "01000000", -- 2035 - 0x7f3  :   64 - 0x40
    "01000000", -- 2036 - 0x7f4  :   64 - 0x40
    "10000000", -- 2037 - 0x7f5  :  128 - 0x80
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "01000000", -- 2040 - 0x7f8  :   64 - 0x40
    "01000000", -- 2041 - 0x7f9  :   64 - 0x40
    "01000000", -- 2042 - 0x7fa  :   64 - 0x40
    "01000000", -- 2043 - 0x7fb  :   64 - 0x40
    "01000000", -- 2044 - 0x7fc  :   64 - 0x40
    "10000000", -- 2045 - 0x7fd  :  128 - 0x80
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000", -- 2047 - 0x7ff  :    0 - 0x0
    "11111111", -- 2048 - 0x800  :  255 - 0xff -- Sprite 0x80
    "11111111", -- 2049 - 0x801  :  255 - 0xff
    "11111111", -- 2050 - 0x802  :  255 - 0xff
    "11111111", -- 2051 - 0x803  :  255 - 0xff
    "11000000", -- 2052 - 0x804  :  192 - 0xc0
    "11000000", -- 2053 - 0x805  :  192 - 0xc0
    "11000000", -- 2054 - 0x806  :  192 - 0xc0
    "11000111", -- 2055 - 0x807  :  199 - 0xc7
    "00000000", -- 2056 - 0x808  :    0 - 0x0
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000000", -- 2059 - 0x80b  :    0 - 0x0
    "00000000", -- 2060 - 0x80c  :    0 - 0x0
    "00011111", -- 2061 - 0x80d  :   31 - 0x1f
    "00010000", -- 2062 - 0x80e  :   16 - 0x10
    "00010111", -- 2063 - 0x80f  :   23 - 0x17
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Sprite 0x81
    "11111111", -- 2065 - 0x811  :  255 - 0xff
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "11111111", -- 2067 - 0x813  :  255 - 0xff
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "11111111", -- 2071 - 0x817  :  255 - 0xff
    "00000000", -- 2072 - 0x818  :    0 - 0x0
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00000000", -- 2075 - 0x81b  :    0 - 0x0
    "00000000", -- 2076 - 0x81c  :    0 - 0x0
    "11111111", -- 2077 - 0x81d  :  255 - 0xff
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "11111111", -- 2079 - 0x81f  :  255 - 0xff
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Sprite 0x82
    "11111111", -- 2081 - 0x821  :  255 - 0xff
    "11111111", -- 2082 - 0x822  :  255 - 0xff
    "11111111", -- 2083 - 0x823  :  255 - 0xff
    "01111111", -- 2084 - 0x824  :  127 - 0x7f
    "00111111", -- 2085 - 0x825  :   63 - 0x3f
    "00011111", -- 2086 - 0x826  :   31 - 0x1f
    "11001111", -- 2087 - 0x827  :  207 - 0xcf
    "00000000", -- 2088 - 0x828  :    0 - 0x0
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "00000000", -- 2091 - 0x82b  :    0 - 0x0
    "00000000", -- 2092 - 0x82c  :    0 - 0x0
    "10000000", -- 2093 - 0x82d  :  128 - 0x80
    "00000000", -- 2094 - 0x82e  :    0 - 0x0
    "11000000", -- 2095 - 0x82f  :  192 - 0xc0
    "11111111", -- 2096 - 0x830  :  255 - 0xff -- Sprite 0x83
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "11111111", -- 2098 - 0x832  :  255 - 0xff
    "11110111", -- 2099 - 0x833  :  247 - 0xf7
    "11110111", -- 2100 - 0x834  :  247 - 0xf7
    "11100010", -- 2101 - 0x835  :  226 - 0xe2
    "11100000", -- 2102 - 0x836  :  224 - 0xe0
    "11000110", -- 2103 - 0x837  :  198 - 0xc6
    "00000000", -- 2104 - 0x838  :    0 - 0x0
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00001000", -- 2109 - 0x83d  :    8 - 0x8
    "00001000", -- 2110 - 0x83e  :    8 - 0x8
    "00010110", -- 2111 - 0x83f  :   22 - 0x16
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Sprite 0x84
    "11111111", -- 2113 - 0x841  :  255 - 0xff
    "11111111", -- 2114 - 0x842  :  255 - 0xff
    "11111111", -- 2115 - 0x843  :  255 - 0xff
    "10111111", -- 2116 - 0x844  :  191 - 0xbf
    "10111111", -- 2117 - 0x845  :  191 - 0xbf
    "00011111", -- 2118 - 0x846  :   31 - 0x1f
    "00011111", -- 2119 - 0x847  :   31 - 0x1f
    "00000000", -- 2120 - 0x848  :    0 - 0x0
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "00000000", -- 2124 - 0x84c  :    0 - 0x0
    "00000000", -- 2125 - 0x84d  :    0 - 0x0
    "01000000", -- 2126 - 0x84e  :   64 - 0x40
    "11000000", -- 2127 - 0x84f  :  192 - 0xc0
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Sprite 0x85
    "11111111", -- 2129 - 0x851  :  255 - 0xff
    "11111111", -- 2130 - 0x852  :  255 - 0xff
    "11111111", -- 2131 - 0x853  :  255 - 0xff
    "11111110", -- 2132 - 0x854  :  254 - 0xfe
    "11111000", -- 2133 - 0x855  :  248 - 0xf8
    "11100000", -- 2134 - 0x856  :  224 - 0xe0
    "11000000", -- 2135 - 0x857  :  192 - 0xc0
    "00000000", -- 2136 - 0x858  :    0 - 0x0
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000001", -- 2141 - 0x85d  :    1 - 0x1
    "00000111", -- 2142 - 0x85e  :    7 - 0x7
    "00001100", -- 2143 - 0x85f  :   12 - 0xc
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11111111", -- 2147 - 0x863  :  255 - 0xff
    "00000111", -- 2148 - 0x864  :    7 - 0x7
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00111111", -- 2150 - 0x866  :   63 - 0x3f
    "11111111", -- 2151 - 0x867  :  255 - 0xff
    "00000000", -- 2152 - 0x868  :    0 - 0x0
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "11000000", -- 2157 - 0x86d  :  192 - 0xc0
    "00111111", -- 2158 - 0x86e  :   63 - 0x3f
    "11111111", -- 2159 - 0x86f  :  255 - 0xff
    "11111111", -- 2160 - 0x870  :  255 - 0xff -- Sprite 0x87
    "11111111", -- 2161 - 0x871  :  255 - 0xff
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "11111111", -- 2164 - 0x874  :  255 - 0xff
    "11111111", -- 2165 - 0x875  :  255 - 0xff
    "00111111", -- 2166 - 0x876  :   63 - 0x3f
    "11001111", -- 2167 - 0x877  :  207 - 0xcf
    "00000000", -- 2168 - 0x878  :    0 - 0x0
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "11000000", -- 2175 - 0x87f  :  192 - 0xc0
    "11111111", -- 2176 - 0x880  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "11111111", -- 2178 - 0x882  :  255 - 0xff
    "11111111", -- 2179 - 0x883  :  255 - 0xff
    "11111111", -- 2180 - 0x884  :  255 - 0xff
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "11111111", -- 2182 - 0x886  :  255 - 0xff
    "11111111", -- 2183 - 0x887  :  255 - 0xff
    "00000000", -- 2184 - 0x888  :    0 - 0x0
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "00000000", -- 2190 - 0x88e  :    0 - 0x0
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "11111111", -- 2192 - 0x890  :  255 - 0xff -- Sprite 0x89
    "11111111", -- 2193 - 0x891  :  255 - 0xff
    "11111111", -- 2194 - 0x892  :  255 - 0xff
    "01110111", -- 2195 - 0x893  :  119 - 0x77
    "00010011", -- 2196 - 0x894  :   19 - 0x13
    "00000001", -- 2197 - 0x895  :    1 - 0x1
    "00010000", -- 2198 - 0x896  :   16 - 0x10
    "00011000", -- 2199 - 0x897  :   24 - 0x18
    "00000000", -- 2200 - 0x898  :    0 - 0x0
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000000", -- 2203 - 0x89b  :    0 - 0x0
    "00000000", -- 2204 - 0x89c  :    0 - 0x0
    "01000100", -- 2205 - 0x89d  :   68 - 0x44
    "01010110", -- 2206 - 0x89e  :   86 - 0x56
    "01011011", -- 2207 - 0x89f  :   91 - 0x5b
    "11111111", -- 2208 - 0x8a0  :  255 - 0xff -- Sprite 0x8a
    "11111111", -- 2209 - 0x8a1  :  255 - 0xff
    "11111111", -- 2210 - 0x8a2  :  255 - 0xff
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "11111111", -- 2212 - 0x8a4  :  255 - 0xff
    "11111111", -- 2213 - 0x8a5  :  255 - 0xff
    "11111111", -- 2214 - 0x8a6  :  255 - 0xff
    "01111111", -- 2215 - 0x8a7  :  127 - 0x7f
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00000000", -- 2222 - 0x8ae  :    0 - 0x0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "11111111", -- 2224 - 0x8b0  :  255 - 0xff -- Sprite 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11111111", -- 2226 - 0x8b2  :  255 - 0xff
    "11110111", -- 2227 - 0x8b3  :  247 - 0xf7
    "11100101", -- 2228 - 0x8b4  :  229 - 0xe5
    "11000001", -- 2229 - 0x8b5  :  193 - 0xc1
    "10000100", -- 2230 - 0x8b6  :  132 - 0x84
    "00001100", -- 2231 - 0x8b7  :   12 - 0xc
    "00000000", -- 2232 - 0x8b8  :    0 - 0x0
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00000000", -- 2234 - 0x8ba  :    0 - 0x0
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00000000", -- 2236 - 0x8bc  :    0 - 0x0
    "00010000", -- 2237 - 0x8bd  :   16 - 0x10
    "00110100", -- 2238 - 0x8be  :   52 - 0x34
    "01101101", -- 2239 - 0x8bf  :  109 - 0x6d
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Sprite 0x8c
    "11111111", -- 2241 - 0x8c1  :  255 - 0xff
    "11111111", -- 2242 - 0x8c2  :  255 - 0xff
    "11111111", -- 2243 - 0x8c3  :  255 - 0xff
    "11111111", -- 2244 - 0x8c4  :  255 - 0xff
    "01111111", -- 2245 - 0x8c5  :  127 - 0x7f
    "01111110", -- 2246 - 0x8c6  :  126 - 0x7e
    "01111110", -- 2247 - 0x8c7  :  126 - 0x7e
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "11111111", -- 2256 - 0x8d0  :  255 - 0xff -- Sprite 0x8d
    "11111111", -- 2257 - 0x8d1  :  255 - 0xff
    "10111111", -- 2258 - 0x8d2  :  191 - 0xbf
    "10110111", -- 2259 - 0x8d3  :  183 - 0xb7
    "00010111", -- 2260 - 0x8d4  :   23 - 0x17
    "00000011", -- 2261 - 0x8d5  :    3 - 0x3
    "00100011", -- 2262 - 0x8d6  :   35 - 0x23
    "00100001", -- 2263 - 0x8d7  :   33 - 0x21
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "00000000", -- 2267 - 0x8db  :    0 - 0x0
    "01000000", -- 2268 - 0x8dc  :   64 - 0x40
    "01001000", -- 2269 - 0x8dd  :   72 - 0x48
    "10101000", -- 2270 - 0x8de  :  168 - 0xa8
    "10101100", -- 2271 - 0x8df  :  172 - 0xac
    "11111111", -- 2272 - 0x8e0  :  255 - 0xff -- Sprite 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11111011", -- 2274 - 0x8e2  :  251 - 0xfb
    "11111001", -- 2275 - 0x8e3  :  249 - 0xf9
    "11111000", -- 2276 - 0x8e4  :  248 - 0xf8
    "11111000", -- 2277 - 0x8e5  :  248 - 0xf8
    "11111000", -- 2278 - 0x8e6  :  248 - 0xf8
    "11111000", -- 2279 - 0x8e7  :  248 - 0xf8
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "00000000", -- 2283 - 0x8eb  :    0 - 0x0
    "00000010", -- 2284 - 0x8ec  :    2 - 0x2
    "00000010", -- 2285 - 0x8ed  :    2 - 0x2
    "00000010", -- 2286 - 0x8ee  :    2 - 0x2
    "00000010", -- 2287 - 0x8ef  :    2 - 0x2
    "11111111", -- 2288 - 0x8f0  :  255 - 0xff -- Sprite 0x8f
    "11111111", -- 2289 - 0x8f1  :  255 - 0xff
    "01111000", -- 2290 - 0x8f2  :  120 - 0x78
    "00111000", -- 2291 - 0x8f3  :   56 - 0x38
    "00011000", -- 2292 - 0x8f4  :   24 - 0x18
    "00001000", -- 2293 - 0x8f5  :    8 - 0x8
    "10000000", -- 2294 - 0x8f6  :  128 - 0x80
    "11000000", -- 2295 - 0x8f7  :  192 - 0xc0
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00000000", -- 2298 - 0x8fa  :    0 - 0x0
    "00000011", -- 2299 - 0x8fb  :    3 - 0x3
    "01000011", -- 2300 - 0x8fc  :   67 - 0x43
    "01100010", -- 2301 - 0x8fd  :   98 - 0x62
    "10110010", -- 2302 - 0x8fe  :  178 - 0xb2
    "11011010", -- 2303 - 0x8ff  :  218 - 0xda
    "11111111", -- 2304 - 0x900  :  255 - 0xff -- Sprite 0x90
    "11111111", -- 2305 - 0x901  :  255 - 0xff
    "00000001", -- 2306 - 0x902  :    1 - 0x1
    "00000001", -- 2307 - 0x903  :    1 - 0x1
    "00000001", -- 2308 - 0x904  :    1 - 0x1
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "11111111", -- 2310 - 0x906  :  255 - 0xff
    "11111111", -- 2311 - 0x907  :  255 - 0xff
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "11111100", -- 2315 - 0x90b  :  252 - 0xfc
    "11111100", -- 2316 - 0x90c  :  252 - 0xfc
    "00000000", -- 2317 - 0x90d  :    0 - 0x0
    "11111111", -- 2318 - 0x90e  :  255 - 0xff
    "11111111", -- 2319 - 0x90f  :  255 - 0xff
    "11111111", -- 2320 - 0x910  :  255 - 0xff -- Sprite 0x91
    "11111111", -- 2321 - 0x911  :  255 - 0xff
    "11111111", -- 2322 - 0x912  :  255 - 0xff
    "11111111", -- 2323 - 0x913  :  255 - 0xff
    "11111111", -- 2324 - 0x914  :  255 - 0xff
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "01111111", -- 2326 - 0x916  :  127 - 0x7f
    "00111111", -- 2327 - 0x917  :   63 - 0x3f
    "00000000", -- 2328 - 0x918  :    0 - 0x0
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "00000000", -- 2330 - 0x91a  :    0 - 0x0
    "00000000", -- 2331 - 0x91b  :    0 - 0x0
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "11000111", -- 2336 - 0x920  :  199 - 0xc7 -- Sprite 0x92
    "11000111", -- 2337 - 0x921  :  199 - 0xc7
    "11000111", -- 2338 - 0x922  :  199 - 0xc7
    "11000111", -- 2339 - 0x923  :  199 - 0xc7
    "11000111", -- 2340 - 0x924  :  199 - 0xc7
    "11000111", -- 2341 - 0x925  :  199 - 0xc7
    "11000111", -- 2342 - 0x926  :  199 - 0xc7
    "11000111", -- 2343 - 0x927  :  199 - 0xc7
    "00010111", -- 2344 - 0x928  :   23 - 0x17
    "00010111", -- 2345 - 0x929  :   23 - 0x17
    "00010111", -- 2346 - 0x92a  :   23 - 0x17
    "00010111", -- 2347 - 0x92b  :   23 - 0x17
    "00010111", -- 2348 - 0x92c  :   23 - 0x17
    "00010111", -- 2349 - 0x92d  :   23 - 0x17
    "00010111", -- 2350 - 0x92e  :   23 - 0x17
    "00010111", -- 2351 - 0x92f  :   23 - 0x17
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Sprite 0x93
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "11111111", -- 2354 - 0x932  :  255 - 0xff
    "11111111", -- 2355 - 0x933  :  255 - 0xff
    "11111001", -- 2356 - 0x934  :  249 - 0xf9
    "11111001", -- 2357 - 0x935  :  249 - 0xf9
    "11111111", -- 2358 - 0x936  :  255 - 0xff
    "11111111", -- 2359 - 0x937  :  255 - 0xff
    "11111111", -- 2360 - 0x938  :  255 - 0xff
    "11111111", -- 2361 - 0x939  :  255 - 0xff
    "11111111", -- 2362 - 0x93a  :  255 - 0xff
    "11111111", -- 2363 - 0x93b  :  255 - 0xff
    "11111001", -- 2364 - 0x93c  :  249 - 0xf9
    "11111001", -- 2365 - 0x93d  :  249 - 0xf9
    "11111111", -- 2366 - 0x93e  :  255 - 0xff
    "11111111", -- 2367 - 0x93f  :  255 - 0xff
    "11110111", -- 2368 - 0x940  :  247 - 0xf7 -- Sprite 0x94
    "11111011", -- 2369 - 0x941  :  251 - 0xfb
    "11111011", -- 2370 - 0x942  :  251 - 0xfb
    "11111101", -- 2371 - 0x943  :  253 - 0xfd
    "11111100", -- 2372 - 0x944  :  252 - 0xfc
    "11111100", -- 2373 - 0x945  :  252 - 0xfc
    "01111100", -- 2374 - 0x946  :  124 - 0x7c
    "01111100", -- 2375 - 0x947  :  124 - 0x7c
    "11110000", -- 2376 - 0x948  :  240 - 0xf0
    "11111000", -- 2377 - 0x949  :  248 - 0xf8
    "11111000", -- 2378 - 0x94a  :  248 - 0xf8
    "11111100", -- 2379 - 0x94b  :  252 - 0xfc
    "11111100", -- 2380 - 0x94c  :  252 - 0xfc
    "11111100", -- 2381 - 0x94d  :  252 - 0xfc
    "01111100", -- 2382 - 0x94e  :  124 - 0x7c
    "01111100", -- 2383 - 0x94f  :  124 - 0x7c
    "11000111", -- 2384 - 0x950  :  199 - 0xc7 -- Sprite 0x95
    "10001111", -- 2385 - 0x951  :  143 - 0x8f
    "10001111", -- 2386 - 0x952  :  143 - 0x8f
    "00011111", -- 2387 - 0x953  :   31 - 0x1f
    "00011111", -- 2388 - 0x954  :   31 - 0x1f
    "00111111", -- 2389 - 0x955  :   63 - 0x3f
    "00111111", -- 2390 - 0x956  :   63 - 0x3f
    "01111111", -- 2391 - 0x957  :  127 - 0x7f
    "00010111", -- 2392 - 0x958  :   23 - 0x17
    "00101111", -- 2393 - 0x959  :   47 - 0x2f
    "00101111", -- 2394 - 0x95a  :   47 - 0x2f
    "01011111", -- 2395 - 0x95b  :   95 - 0x5f
    "01011111", -- 2396 - 0x95c  :   95 - 0x5f
    "10111111", -- 2397 - 0x95d  :  191 - 0xbf
    "10111111", -- 2398 - 0x95e  :  191 - 0xbf
    "01111111", -- 2399 - 0x95f  :  127 - 0x7f
    "00001111", -- 2400 - 0x960  :   15 - 0xf -- Sprite 0x96
    "00001111", -- 2401 - 0x961  :   15 - 0xf
    "10000111", -- 2402 - 0x962  :  135 - 0x87
    "10000111", -- 2403 - 0x963  :  135 - 0x87
    "11000010", -- 2404 - 0x964  :  194 - 0xc2
    "11000010", -- 2405 - 0x965  :  194 - 0xc2
    "11100000", -- 2406 - 0x966  :  224 - 0xe0
    "11100000", -- 2407 - 0x967  :  224 - 0xe0
    "01100000", -- 2408 - 0x968  :   96 - 0x60
    "01100000", -- 2409 - 0x969  :   96 - 0x60
    "10110000", -- 2410 - 0x96a  :  176 - 0xb0
    "10110000", -- 2411 - 0x96b  :  176 - 0xb0
    "11011000", -- 2412 - 0x96c  :  216 - 0xd8
    "11011000", -- 2413 - 0x96d  :  216 - 0xd8
    "11101100", -- 2414 - 0x96e  :  236 - 0xec
    "11101100", -- 2415 - 0x96f  :  236 - 0xec
    "10000011", -- 2416 - 0x970  :  131 - 0x83 -- Sprite 0x97
    "10001111", -- 2417 - 0x971  :  143 - 0x8f
    "00001111", -- 2418 - 0x972  :   15 - 0xf
    "00011111", -- 2419 - 0x973  :   31 - 0x1f
    "00011111", -- 2420 - 0x974  :   31 - 0x1f
    "00111111", -- 2421 - 0x975  :   63 - 0x3f
    "00111111", -- 2422 - 0x976  :   63 - 0x3f
    "00111111", -- 2423 - 0x977  :   63 - 0x3f
    "00110011", -- 2424 - 0x978  :   51 - 0x33
    "00101111", -- 2425 - 0x979  :   47 - 0x2f
    "01101111", -- 2426 - 0x97a  :  111 - 0x6f
    "01011111", -- 2427 - 0x97b  :   95 - 0x5f
    "11011111", -- 2428 - 0x97c  :  223 - 0xdf
    "10111111", -- 2429 - 0x97d  :  191 - 0xbf
    "10111111", -- 2430 - 0x97e  :  191 - 0xbf
    "10111111", -- 2431 - 0x97f  :  191 - 0xbf
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Sprite 0x98
    "11111111", -- 2433 - 0x981  :  255 - 0xff
    "11111111", -- 2434 - 0x982  :  255 - 0xff
    "11111110", -- 2435 - 0x983  :  254 - 0xfe
    "11111001", -- 2436 - 0x984  :  249 - 0xf9
    "11100111", -- 2437 - 0x985  :  231 - 0xe7
    "11111100", -- 2438 - 0x986  :  252 - 0xfc
    "11110000", -- 2439 - 0x987  :  240 - 0xf0
    "11111111", -- 2440 - 0x988  :  255 - 0xff
    "11111111", -- 2441 - 0x989  :  255 - 0xff
    "11111111", -- 2442 - 0x98a  :  255 - 0xff
    "11111110", -- 2443 - 0x98b  :  254 - 0xfe
    "11111001", -- 2444 - 0x98c  :  249 - 0xf9
    "11100111", -- 2445 - 0x98d  :  231 - 0xe7
    "11111100", -- 2446 - 0x98e  :  252 - 0xfc
    "11110011", -- 2447 - 0x98f  :  243 - 0xf3
    "11110111", -- 2448 - 0x990  :  247 - 0xf7 -- Sprite 0x99
    "11111011", -- 2449 - 0x991  :  251 - 0xfb
    "11111011", -- 2450 - 0x992  :  251 - 0xfb
    "01110011", -- 2451 - 0x993  :  115 - 0x73
    "11000001", -- 2452 - 0x994  :  193 - 0xc1
    "00000011", -- 2453 - 0x995  :    3 - 0x3
    "00001111", -- 2454 - 0x996  :   15 - 0xf
    "00111111", -- 2455 - 0x997  :   63 - 0x3f
    "11110000", -- 2456 - 0x998  :  240 - 0xf0
    "11111000", -- 2457 - 0x999  :  248 - 0xf8
    "11111000", -- 2458 - 0x99a  :  248 - 0xf8
    "01110000", -- 2459 - 0x99b  :  112 - 0x70
    "11001100", -- 2460 - 0x99c  :  204 - 0xcc
    "00110000", -- 2461 - 0x99d  :   48 - 0x30
    "11000000", -- 2462 - 0x99e  :  192 - 0xc0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "11111111", -- 2464 - 0x9a0  :  255 - 0xff -- Sprite 0x9a
    "11111111", -- 2465 - 0x9a1  :  255 - 0xff
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "10000000", -- 2467 - 0x9a3  :  128 - 0x80
    "10000000", -- 2468 - 0x9a4  :  128 - 0x80
    "10000000", -- 2469 - 0x9a5  :  128 - 0x80
    "10001111", -- 2470 - 0x9a6  :  143 - 0x8f
    "10001111", -- 2471 - 0x9a7  :  143 - 0x8f
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00111111", -- 2476 - 0x9ac  :   63 - 0x3f
    "00100000", -- 2477 - 0x9ad  :   32 - 0x20
    "00101111", -- 2478 - 0x9ae  :   47 - 0x2f
    "00101111", -- 2479 - 0x9af  :   47 - 0x2f
    "11111111", -- 2480 - 0x9b0  :  255 - 0xff -- Sprite 0x9b
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "11111111", -- 2482 - 0x9b2  :  255 - 0xff
    "00001111", -- 2483 - 0x9b3  :   15 - 0xf
    "00001111", -- 2484 - 0x9b4  :   15 - 0xf
    "00000111", -- 2485 - 0x9b5  :    7 - 0x7
    "11110111", -- 2486 - 0x9b6  :  247 - 0xf7
    "11110001", -- 2487 - 0x9b7  :  241 - 0xf1
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "11100000", -- 2492 - 0x9bc  :  224 - 0xe0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "11110000", -- 2494 - 0x9be  :  240 - 0xf0
    "11110000", -- 2495 - 0x9bf  :  240 - 0xf0
    "00011100", -- 2496 - 0x9c0  :   28 - 0x1c -- Sprite 0x9c
    "00011110", -- 2497 - 0x9c1  :   30 - 0x1e
    "00011111", -- 2498 - 0x9c2  :   31 - 0x1f
    "00011111", -- 2499 - 0x9c3  :   31 - 0x1f
    "00011111", -- 2500 - 0x9c4  :   31 - 0x1f
    "00011111", -- 2501 - 0x9c5  :   31 - 0x1f
    "00011111", -- 2502 - 0x9c6  :   31 - 0x1f
    "00011111", -- 2503 - 0x9c7  :   31 - 0x1f
    "01011101", -- 2504 - 0x9c8  :   93 - 0x5d
    "01011110", -- 2505 - 0x9c9  :   94 - 0x5e
    "01011111", -- 2506 - 0x9ca  :   95 - 0x5f
    "01011111", -- 2507 - 0x9cb  :   95 - 0x5f
    "01011111", -- 2508 - 0x9cc  :   95 - 0x5f
    "01011111", -- 2509 - 0x9cd  :   95 - 0x5f
    "01011111", -- 2510 - 0x9ce  :   95 - 0x5f
    "01011111", -- 2511 - 0x9cf  :   95 - 0x5f
    "00111110", -- 2512 - 0x9d0  :   62 - 0x3e -- Sprite 0x9d
    "00011100", -- 2513 - 0x9d1  :   28 - 0x1c
    "00001000", -- 2514 - 0x9d2  :    8 - 0x8
    "10000000", -- 2515 - 0x9d3  :  128 - 0x80
    "11000001", -- 2516 - 0x9d4  :  193 - 0xc1
    "11100011", -- 2517 - 0x9d5  :  227 - 0xe3
    "11110111", -- 2518 - 0x9d6  :  247 - 0xf7
    "11111111", -- 2519 - 0x9d7  :  255 - 0xff
    "10000000", -- 2520 - 0x9d8  :  128 - 0x80
    "11000001", -- 2521 - 0x9d9  :  193 - 0xc1
    "01100011", -- 2522 - 0x9da  :   99 - 0x63
    "10110110", -- 2523 - 0x9db  :  182 - 0xb6
    "11011001", -- 2524 - 0x9dc  :  217 - 0xd9
    "11101011", -- 2525 - 0x9dd  :  235 - 0xeb
    "11110111", -- 2526 - 0x9de  :  247 - 0xf7
    "11111111", -- 2527 - 0x9df  :  255 - 0xff
    "00011100", -- 2528 - 0x9e0  :   28 - 0x1c -- Sprite 0x9e
    "00111100", -- 2529 - 0x9e1  :   60 - 0x3c
    "01111100", -- 2530 - 0x9e2  :  124 - 0x7c
    "11111100", -- 2531 - 0x9e3  :  252 - 0xfc
    "11111100", -- 2532 - 0x9e4  :  252 - 0xfc
    "11111100", -- 2533 - 0x9e5  :  252 - 0xfc
    "11111100", -- 2534 - 0x9e6  :  252 - 0xfc
    "11111100", -- 2535 - 0x9e7  :  252 - 0xfc
    "11011101", -- 2536 - 0x9e8  :  221 - 0xdd
    "10111101", -- 2537 - 0x9e9  :  189 - 0xbd
    "01111101", -- 2538 - 0x9ea  :  125 - 0x7d
    "11111101", -- 2539 - 0x9eb  :  253 - 0xfd
    "11111101", -- 2540 - 0x9ec  :  253 - 0xfd
    "11111101", -- 2541 - 0x9ed  :  253 - 0xfd
    "11111101", -- 2542 - 0x9ee  :  253 - 0xfd
    "11111101", -- 2543 - 0x9ef  :  253 - 0xfd
    "01111100", -- 2544 - 0x9f0  :  124 - 0x7c -- Sprite 0x9f
    "01111100", -- 2545 - 0x9f1  :  124 - 0x7c
    "01111000", -- 2546 - 0x9f2  :  120 - 0x78
    "01111000", -- 2547 - 0x9f3  :  120 - 0x78
    "01110001", -- 2548 - 0x9f4  :  113 - 0x71
    "01110001", -- 2549 - 0x9f5  :  113 - 0x71
    "01100011", -- 2550 - 0x9f6  :   99 - 0x63
    "01100011", -- 2551 - 0x9f7  :   99 - 0x63
    "00000001", -- 2552 - 0x9f8  :    1 - 0x1
    "00000001", -- 2553 - 0x9f9  :    1 - 0x1
    "00000010", -- 2554 - 0x9fa  :    2 - 0x2
    "00000010", -- 2555 - 0x9fb  :    2 - 0x2
    "00000101", -- 2556 - 0x9fc  :    5 - 0x5
    "00000101", -- 2557 - 0x9fd  :    5 - 0x5
    "00001011", -- 2558 - 0x9fe  :   11 - 0xb
    "00001011", -- 2559 - 0x9ff  :   11 - 0xb
    "01110001", -- 2560 - 0xa00  :  113 - 0x71 -- Sprite 0xa0
    "01110000", -- 2561 - 0xa01  :  112 - 0x70
    "11111000", -- 2562 - 0xa02  :  248 - 0xf8
    "11111000", -- 2563 - 0xa03  :  248 - 0xf8
    "11111100", -- 2564 - 0xa04  :  252 - 0xfc
    "11111100", -- 2565 - 0xa05  :  252 - 0xfc
    "11111110", -- 2566 - 0xa06  :  254 - 0xfe
    "11111110", -- 2567 - 0xa07  :  254 - 0xfe
    "01110100", -- 2568 - 0xa08  :  116 - 0x74
    "01110110", -- 2569 - 0xa09  :  118 - 0x76
    "11111010", -- 2570 - 0xa0a  :  250 - 0xfa
    "11111011", -- 2571 - 0xa0b  :  251 - 0xfb
    "11111101", -- 2572 - 0xa0c  :  253 - 0xfd
    "11111101", -- 2573 - 0xa0d  :  253 - 0xfd
    "11111110", -- 2574 - 0xa0e  :  254 - 0xfe
    "11111110", -- 2575 - 0xa0f  :  254 - 0xfe
    "11111000", -- 2576 - 0xa10  :  248 - 0xf8 -- Sprite 0xa1
    "11111000", -- 2577 - 0xa11  :  248 - 0xf8
    "11111000", -- 2578 - 0xa12  :  248 - 0xf8
    "01111000", -- 2579 - 0xa13  :  120 - 0x78
    "01111000", -- 2580 - 0xa14  :  120 - 0x78
    "00111000", -- 2581 - 0xa15  :   56 - 0x38
    "00111000", -- 2582 - 0xa16  :   56 - 0x38
    "00011000", -- 2583 - 0xa17  :   24 - 0x18
    "00000010", -- 2584 - 0xa18  :    2 - 0x2
    "00000010", -- 2585 - 0xa19  :    2 - 0x2
    "00000010", -- 2586 - 0xa1a  :    2 - 0x2
    "00000010", -- 2587 - 0xa1b  :    2 - 0x2
    "00000010", -- 2588 - 0xa1c  :    2 - 0x2
    "10000010", -- 2589 - 0xa1d  :  130 - 0x82
    "10000010", -- 2590 - 0xa1e  :  130 - 0x82
    "11000010", -- 2591 - 0xa1f  :  194 - 0xc2
    "11100000", -- 2592 - 0xa20  :  224 - 0xe0 -- Sprite 0xa2
    "11110000", -- 2593 - 0xa21  :  240 - 0xf0
    "11111000", -- 2594 - 0xa22  :  248 - 0xf8
    "11111000", -- 2595 - 0xa23  :  248 - 0xf8
    "11111100", -- 2596 - 0xa24  :  252 - 0xfc
    "11111100", -- 2597 - 0xa25  :  252 - 0xfc
    "11111110", -- 2598 - 0xa26  :  254 - 0xfe
    "11111111", -- 2599 - 0xa27  :  255 - 0xff
    "11101010", -- 2600 - 0xa28  :  234 - 0xea
    "11110110", -- 2601 - 0xa29  :  246 - 0xf6
    "11111010", -- 2602 - 0xa2a  :  250 - 0xfa
    "11111010", -- 2603 - 0xa2b  :  250 - 0xfa
    "11111100", -- 2604 - 0xa2c  :  252 - 0xfc
    "11111100", -- 2605 - 0xa2d  :  252 - 0xfc
    "11111110", -- 2606 - 0xa2e  :  254 - 0xfe
    "11111111", -- 2607 - 0xa2f  :  255 - 0xff
    "11111111", -- 2608 - 0xa30  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 2609 - 0xa31  :  255 - 0xff
    "11111111", -- 2610 - 0xa32  :  255 - 0xff
    "11111111", -- 2611 - 0xa33  :  255 - 0xff
    "11111111", -- 2612 - 0xa34  :  255 - 0xff
    "11111111", -- 2613 - 0xa35  :  255 - 0xff
    "11111111", -- 2614 - 0xa36  :  255 - 0xff
    "11111111", -- 2615 - 0xa37  :  255 - 0xff
    "11111111", -- 2616 - 0xa38  :  255 - 0xff
    "11111111", -- 2617 - 0xa39  :  255 - 0xff
    "11111111", -- 2618 - 0xa3a  :  255 - 0xff
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "00011111", -- 2624 - 0xa40  :   31 - 0x1f -- Sprite 0xa4
    "00011111", -- 2625 - 0xa41  :   31 - 0x1f
    "00011111", -- 2626 - 0xa42  :   31 - 0x1f
    "00011111", -- 2627 - 0xa43  :   31 - 0x1f
    "00011111", -- 2628 - 0xa44  :   31 - 0x1f
    "00011111", -- 2629 - 0xa45  :   31 - 0x1f
    "00011111", -- 2630 - 0xa46  :   31 - 0x1f
    "00011111", -- 2631 - 0xa47  :   31 - 0x1f
    "01000000", -- 2632 - 0xa48  :   64 - 0x40
    "01000000", -- 2633 - 0xa49  :   64 - 0x40
    "01000000", -- 2634 - 0xa4a  :   64 - 0x40
    "01000000", -- 2635 - 0xa4b  :   64 - 0x40
    "01000000", -- 2636 - 0xa4c  :   64 - 0x40
    "01000000", -- 2637 - 0xa4d  :   64 - 0x40
    "01000000", -- 2638 - 0xa4e  :   64 - 0x40
    "01000000", -- 2639 - 0xa4f  :   64 - 0x40
    "11111000", -- 2640 - 0xa50  :  248 - 0xf8 -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "11111000", -- 2643 - 0xa53  :  248 - 0xf8
    "11111000", -- 2644 - 0xa54  :  248 - 0xf8
    "11111000", -- 2645 - 0xa55  :  248 - 0xf8
    "11111000", -- 2646 - 0xa56  :  248 - 0xf8
    "11111000", -- 2647 - 0xa57  :  248 - 0xf8
    "11111000", -- 2648 - 0xa58  :  248 - 0xf8
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111000", -- 2651 - 0xa5b  :  248 - 0xf8
    "11111011", -- 2652 - 0xa5c  :  251 - 0xfb
    "11111010", -- 2653 - 0xa5d  :  250 - 0xfa
    "11111010", -- 2654 - 0xa5e  :  250 - 0xfa
    "11111010", -- 2655 - 0xa5f  :  250 - 0xfa
    "11111100", -- 2656 - 0xa60  :  252 - 0xfc -- Sprite 0xa6
    "11111000", -- 2657 - 0xa61  :  248 - 0xf8
    "11110000", -- 2658 - 0xa62  :  240 - 0xf0
    "00000001", -- 2659 - 0xa63  :    1 - 0x1
    "00000001", -- 2660 - 0xa64  :    1 - 0x1
    "00000011", -- 2661 - 0xa65  :    3 - 0x3
    "11000011", -- 2662 - 0xa66  :  195 - 0xc3
    "10000111", -- 2663 - 0xa67  :  135 - 0x87
    "11111100", -- 2664 - 0xa68  :  252 - 0xfc
    "11111010", -- 2665 - 0xa69  :  250 - 0xfa
    "11110110", -- 2666 - 0xa6a  :  246 - 0xf6
    "00001101", -- 2667 - 0xa6b  :   13 - 0xd
    "11111001", -- 2668 - 0xa6c  :  249 - 0xf9
    "00000011", -- 2669 - 0xa6d  :    3 - 0x3
    "00010011", -- 2670 - 0xa6e  :   19 - 0x13
    "00110111", -- 2671 - 0xa6f  :   55 - 0x37
    "01111111", -- 2672 - 0xa70  :  127 - 0x7f -- Sprite 0xa7
    "11111001", -- 2673 - 0xa71  :  249 - 0xf9
    "11111001", -- 2674 - 0xa72  :  249 - 0xf9
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111110", -- 2676 - 0xa74  :  254 - 0xfe
    "11111100", -- 2677 - 0xa75  :  252 - 0xfc
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "01111111", -- 2680 - 0xa78  :  127 - 0x7f
    "11111001", -- 2681 - 0xa79  :  249 - 0xf9
    "11111001", -- 2682 - 0xa7a  :  249 - 0xf9
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111110", -- 2684 - 0xa7c  :  254 - 0xfe
    "11111100", -- 2685 - 0xa7d  :  252 - 0xfc
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "11110000", -- 2688 - 0xa80  :  240 - 0xf0 -- Sprite 0xa8
    "11110000", -- 2689 - 0xa81  :  240 - 0xf0
    "11111000", -- 2690 - 0xa82  :  248 - 0xf8
    "01111000", -- 2691 - 0xa83  :  120 - 0x78
    "11111100", -- 2692 - 0xa84  :  252 - 0xfc
    "11110100", -- 2693 - 0xa85  :  244 - 0xf4
    "11110110", -- 2694 - 0xa86  :  246 - 0xf6
    "11111010", -- 2695 - 0xa87  :  250 - 0xfa
    "11110110", -- 2696 - 0xa88  :  246 - 0xf6
    "11110110", -- 2697 - 0xa89  :  246 - 0xf6
    "11111011", -- 2698 - 0xa8a  :  251 - 0xfb
    "01111011", -- 2699 - 0xa8b  :  123 - 0x7b
    "11111101", -- 2700 - 0xa8c  :  253 - 0xfd
    "11110101", -- 2701 - 0xa8d  :  245 - 0xf5
    "11110110", -- 2702 - 0xa8e  :  246 - 0xf6
    "11111010", -- 2703 - 0xa8f  :  250 - 0xfa
    "00111111", -- 2704 - 0xa90  :   63 - 0x3f -- Sprite 0xa9
    "00111111", -- 2705 - 0xa91  :   63 - 0x3f
    "00111111", -- 2706 - 0xa92  :   63 - 0x3f
    "00111111", -- 2707 - 0xa93  :   63 - 0x3f
    "00111111", -- 2708 - 0xa94  :   63 - 0x3f
    "00011111", -- 2709 - 0xa95  :   31 - 0x1f
    "00001111", -- 2710 - 0xa96  :   15 - 0xf
    "00000111", -- 2711 - 0xa97  :    7 - 0x7
    "10111111", -- 2712 - 0xa98  :  191 - 0xbf
    "10111111", -- 2713 - 0xa99  :  191 - 0xbf
    "00111111", -- 2714 - 0xa9a  :   63 - 0x3f
    "00111111", -- 2715 - 0xa9b  :   63 - 0x3f
    "10111111", -- 2716 - 0xa9c  :  191 - 0xbf
    "10011111", -- 2717 - 0xa9d  :  159 - 0x9f
    "11001111", -- 2718 - 0xa9e  :  207 - 0xcf
    "11010111", -- 2719 - 0xa9f  :  215 - 0xd7
    "11100000", -- 2720 - 0xaa0  :  224 - 0xe0 -- Sprite 0xaa
    "11111000", -- 2721 - 0xaa1  :  248 - 0xf8
    "11111111", -- 2722 - 0xaa2  :  255 - 0xff
    "11110011", -- 2723 - 0xaa3  :  243 - 0xf3
    "11111100", -- 2724 - 0xaa4  :  252 - 0xfc
    "11111111", -- 2725 - 0xaa5  :  255 - 0xff
    "11111111", -- 2726 - 0xaa6  :  255 - 0xff
    "11111111", -- 2727 - 0xaa7  :  255 - 0xff
    "11100100", -- 2728 - 0xaa8  :  228 - 0xe4
    "11111000", -- 2729 - 0xaa9  :  248 - 0xf8
    "11111111", -- 2730 - 0xaaa  :  255 - 0xff
    "11110011", -- 2731 - 0xaab  :  243 - 0xf3
    "11111100", -- 2732 - 0xaac  :  252 - 0xfc
    "11111111", -- 2733 - 0xaad  :  255 - 0xff
    "11111111", -- 2734 - 0xaae  :  255 - 0xff
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "11111111", -- 2736 - 0xab0  :  255 - 0xff -- Sprite 0xab
    "11111111", -- 2737 - 0xab1  :  255 - 0xff
    "00111111", -- 2738 - 0xab2  :   63 - 0x3f
    "11001111", -- 2739 - 0xab3  :  207 - 0xcf
    "11110011", -- 2740 - 0xab4  :  243 - 0xf3
    "00111101", -- 2741 - 0xab5  :   61 - 0x3d
    "11011000", -- 2742 - 0xab6  :  216 - 0xd8
    "10110000", -- 2743 - 0xab7  :  176 - 0xb0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "11000000", -- 2747 - 0xabb  :  192 - 0xc0
    "11110000", -- 2748 - 0xabc  :  240 - 0xf0
    "00111100", -- 2749 - 0xabd  :   60 - 0x3c
    "11011000", -- 2750 - 0xabe  :  216 - 0xd8
    "10110110", -- 2751 - 0xabf  :  182 - 0xb6
    "10001111", -- 2752 - 0xac0  :  143 - 0x8f -- Sprite 0xac
    "11101111", -- 2753 - 0xac1  :  239 - 0xef
    "11100000", -- 2754 - 0xac2  :  224 - 0xe0
    "11111000", -- 2755 - 0xac3  :  248 - 0xf8
    "11111000", -- 2756 - 0xac4  :  248 - 0xf8
    "11111111", -- 2757 - 0xac5  :  255 - 0xff
    "11111111", -- 2758 - 0xac6  :  255 - 0xff
    "11111111", -- 2759 - 0xac7  :  255 - 0xff
    "00001111", -- 2760 - 0xac8  :   15 - 0xf
    "00001111", -- 2761 - 0xac9  :   15 - 0xf
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000011", -- 2763 - 0xacb  :    3 - 0x3
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "11110001", -- 2768 - 0xad0  :  241 - 0xf1 -- Sprite 0xad
    "11110001", -- 2769 - 0xad1  :  241 - 0xf1
    "00000001", -- 2770 - 0xad2  :    1 - 0x1
    "00000001", -- 2771 - 0xad3  :    1 - 0x1
    "00000001", -- 2772 - 0xad4  :    1 - 0x1
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "11110100", -- 2776 - 0xad8  :  244 - 0xf4
    "11110100", -- 2777 - 0xad9  :  244 - 0xf4
    "00000100", -- 2778 - 0xada  :    4 - 0x4
    "11111100", -- 2779 - 0xadb  :  252 - 0xfc
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00011111", -- 2784 - 0xae0  :   31 - 0x1f -- Sprite 0xae
    "00011111", -- 2785 - 0xae1  :   31 - 0x1f
    "00011111", -- 2786 - 0xae2  :   31 - 0x1f
    "00011111", -- 2787 - 0xae3  :   31 - 0x1f
    "00011111", -- 2788 - 0xae4  :   31 - 0x1f
    "00011111", -- 2789 - 0xae5  :   31 - 0x1f
    "00011111", -- 2790 - 0xae6  :   31 - 0x1f
    "00011111", -- 2791 - 0xae7  :   31 - 0x1f
    "01011111", -- 2792 - 0xae8  :   95 - 0x5f
    "01011111", -- 2793 - 0xae9  :   95 - 0x5f
    "01011111", -- 2794 - 0xaea  :   95 - 0x5f
    "01011111", -- 2795 - 0xaeb  :   95 - 0x5f
    "01011111", -- 2796 - 0xaec  :   95 - 0x5f
    "01011111", -- 2797 - 0xaed  :   95 - 0x5f
    "01011111", -- 2798 - 0xaee  :   95 - 0x5f
    "01011111", -- 2799 - 0xaef  :   95 - 0x5f
    "11111100", -- 2800 - 0xaf0  :  252 - 0xfc -- Sprite 0xaf
    "11111100", -- 2801 - 0xaf1  :  252 - 0xfc
    "11111100", -- 2802 - 0xaf2  :  252 - 0xfc
    "11111100", -- 2803 - 0xaf3  :  252 - 0xfc
    "11110100", -- 2804 - 0xaf4  :  244 - 0xf4
    "11110100", -- 2805 - 0xaf5  :  244 - 0xf4
    "11110100", -- 2806 - 0xaf6  :  244 - 0xf4
    "11110100", -- 2807 - 0xaf7  :  244 - 0xf4
    "11111101", -- 2808 - 0xaf8  :  253 - 0xfd
    "11111101", -- 2809 - 0xaf9  :  253 - 0xfd
    "11111101", -- 2810 - 0xafa  :  253 - 0xfd
    "11111101", -- 2811 - 0xafb  :  253 - 0xfd
    "11110101", -- 2812 - 0xafc  :  245 - 0xf5
    "11110101", -- 2813 - 0xafd  :  245 - 0xf5
    "11110101", -- 2814 - 0xafe  :  245 - 0xf5
    "11110101", -- 2815 - 0xaff  :  245 - 0xf5
    "00001100", -- 2816 - 0xb00  :   12 - 0xc -- Sprite 0xb0
    "00011100", -- 2817 - 0xb01  :   28 - 0x1c
    "00001100", -- 2818 - 0xb02  :   12 - 0xc
    "00001100", -- 2819 - 0xb03  :   12 - 0xc
    "00001100", -- 2820 - 0xb04  :   12 - 0xc
    "00001100", -- 2821 - 0xb05  :   12 - 0xc
    "00111111", -- 2822 - 0xb06  :   63 - 0x3f
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00001100", -- 2824 - 0xb08  :   12 - 0xc
    "00011100", -- 2825 - 0xb09  :   28 - 0x1c
    "00001100", -- 2826 - 0xb0a  :   12 - 0xc
    "00001100", -- 2827 - 0xb0b  :   12 - 0xc
    "00001100", -- 2828 - 0xb0c  :   12 - 0xc
    "00001100", -- 2829 - 0xb0d  :   12 - 0xc
    "00111111", -- 2830 - 0xb0e  :   63 - 0x3f
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00111110", -- 2832 - 0xb10  :   62 - 0x3e -- Sprite 0xb1
    "01100011", -- 2833 - 0xb11  :   99 - 0x63
    "00000111", -- 2834 - 0xb12  :    7 - 0x7
    "00011110", -- 2835 - 0xb13  :   30 - 0x1e
    "00111100", -- 2836 - 0xb14  :   60 - 0x3c
    "01110000", -- 2837 - 0xb15  :  112 - 0x70
    "01111111", -- 2838 - 0xb16  :  127 - 0x7f
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00111110", -- 2840 - 0xb18  :   62 - 0x3e
    "01100011", -- 2841 - 0xb19  :   99 - 0x63
    "00000111", -- 2842 - 0xb1a  :    7 - 0x7
    "00011110", -- 2843 - 0xb1b  :   30 - 0x1e
    "00111100", -- 2844 - 0xb1c  :   60 - 0x3c
    "01110000", -- 2845 - 0xb1d  :  112 - 0x70
    "01111111", -- 2846 - 0xb1e  :  127 - 0x7f
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "01111110", -- 2848 - 0xb20  :  126 - 0x7e -- Sprite 0xb2
    "01100011", -- 2849 - 0xb21  :   99 - 0x63
    "01100011", -- 2850 - 0xb22  :   99 - 0x63
    "01100011", -- 2851 - 0xb23  :   99 - 0x63
    "01111110", -- 2852 - 0xb24  :  126 - 0x7e
    "01100000", -- 2853 - 0xb25  :   96 - 0x60
    "01100000", -- 2854 - 0xb26  :   96 - 0x60
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "01111110", -- 2856 - 0xb28  :  126 - 0x7e
    "01100011", -- 2857 - 0xb29  :   99 - 0x63
    "01100011", -- 2858 - 0xb2a  :   99 - 0x63
    "01100011", -- 2859 - 0xb2b  :   99 - 0x63
    "01111110", -- 2860 - 0xb2c  :  126 - 0x7e
    "01100000", -- 2861 - 0xb2d  :   96 - 0x60
    "01100000", -- 2862 - 0xb2e  :   96 - 0x60
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "01100011", -- 2864 - 0xb30  :   99 - 0x63 -- Sprite 0xb3
    "01100011", -- 2865 - 0xb31  :   99 - 0x63
    "01100011", -- 2866 - 0xb32  :   99 - 0x63
    "01100011", -- 2867 - 0xb33  :   99 - 0x63
    "01100011", -- 2868 - 0xb34  :   99 - 0x63
    "01100011", -- 2869 - 0xb35  :   99 - 0x63
    "00111110", -- 2870 - 0xb36  :   62 - 0x3e
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "01100011", -- 2872 - 0xb38  :   99 - 0x63
    "01100011", -- 2873 - 0xb39  :   99 - 0x63
    "01100011", -- 2874 - 0xb3a  :   99 - 0x63
    "01100011", -- 2875 - 0xb3b  :   99 - 0x63
    "01100011", -- 2876 - 0xb3c  :   99 - 0x63
    "01100011", -- 2877 - 0xb3d  :   99 - 0x63
    "00111110", -- 2878 - 0xb3e  :   62 - 0x3e
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "01100011", -- 2880 - 0xb40  :   99 - 0x63 -- Sprite 0xb4
    "01100011", -- 2881 - 0xb41  :   99 - 0x63
    "01100011", -- 2882 - 0xb42  :   99 - 0x63
    "01111111", -- 2883 - 0xb43  :  127 - 0x7f
    "01100011", -- 2884 - 0xb44  :   99 - 0x63
    "01100011", -- 2885 - 0xb45  :   99 - 0x63
    "01100011", -- 2886 - 0xb46  :   99 - 0x63
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "01100011", -- 2888 - 0xb48  :   99 - 0x63
    "01100011", -- 2889 - 0xb49  :   99 - 0x63
    "01100011", -- 2890 - 0xb4a  :   99 - 0x63
    "01111111", -- 2891 - 0xb4b  :  127 - 0x7f
    "01100011", -- 2892 - 0xb4c  :   99 - 0x63
    "01100011", -- 2893 - 0xb4d  :   99 - 0x63
    "01100011", -- 2894 - 0xb4e  :   99 - 0x63
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00111111", -- 2896 - 0xb50  :   63 - 0x3f -- Sprite 0xb5
    "00001100", -- 2897 - 0xb51  :   12 - 0xc
    "00001100", -- 2898 - 0xb52  :   12 - 0xc
    "00001100", -- 2899 - 0xb53  :   12 - 0xc
    "00001100", -- 2900 - 0xb54  :   12 - 0xc
    "00001100", -- 2901 - 0xb55  :   12 - 0xc
    "00111111", -- 2902 - 0xb56  :   63 - 0x3f
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00111111", -- 2904 - 0xb58  :   63 - 0x3f
    "00001100", -- 2905 - 0xb59  :   12 - 0xc
    "00001100", -- 2906 - 0xb5a  :   12 - 0xc
    "00001100", -- 2907 - 0xb5b  :   12 - 0xc
    "00001100", -- 2908 - 0xb5c  :   12 - 0xc
    "00001100", -- 2909 - 0xb5d  :   12 - 0xc
    "00111111", -- 2910 - 0xb5e  :   63 - 0x3f
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Sprite 0xb6
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "01111110", -- 2915 - 0xb63  :  126 - 0x7e
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "01111110", -- 2923 - 0xb6b  :  126 - 0x7e
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00111100", -- 2928 - 0xb70  :   60 - 0x3c -- Sprite 0xb7
    "01100110", -- 2929 - 0xb71  :  102 - 0x66
    "01100000", -- 2930 - 0xb72  :   96 - 0x60
    "00111110", -- 2931 - 0xb73  :   62 - 0x3e
    "00000011", -- 2932 - 0xb74  :    3 - 0x3
    "01100011", -- 2933 - 0xb75  :   99 - 0x63
    "00111110", -- 2934 - 0xb76  :   62 - 0x3e
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00111100", -- 2936 - 0xb78  :   60 - 0x3c
    "01100110", -- 2937 - 0xb79  :  102 - 0x66
    "01100000", -- 2938 - 0xb7a  :   96 - 0x60
    "00111110", -- 2939 - 0xb7b  :   62 - 0x3e
    "00000011", -- 2940 - 0xb7c  :    3 - 0x3
    "01100011", -- 2941 - 0xb7d  :   99 - 0x63
    "00111110", -- 2942 - 0xb7e  :   62 - 0x3e
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00011110", -- 2944 - 0xb80  :   30 - 0x1e -- Sprite 0xb8
    "00110011", -- 2945 - 0xb81  :   51 - 0x33
    "01100000", -- 2946 - 0xb82  :   96 - 0x60
    "01100000", -- 2947 - 0xb83  :   96 - 0x60
    "01100000", -- 2948 - 0xb84  :   96 - 0x60
    "00110011", -- 2949 - 0xb85  :   51 - 0x33
    "00011110", -- 2950 - 0xb86  :   30 - 0x1e
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00011110", -- 2952 - 0xb88  :   30 - 0x1e
    "00110011", -- 2953 - 0xb89  :   51 - 0x33
    "01100000", -- 2954 - 0xb8a  :   96 - 0x60
    "01100000", -- 2955 - 0xb8b  :   96 - 0x60
    "01100000", -- 2956 - 0xb8c  :   96 - 0x60
    "00110011", -- 2957 - 0xb8d  :   51 - 0x33
    "00011110", -- 2958 - 0xb8e  :   30 - 0x1e
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00111110", -- 2960 - 0xb90  :   62 - 0x3e -- Sprite 0xb9
    "01100011", -- 2961 - 0xb91  :   99 - 0x63
    "01100011", -- 2962 - 0xb92  :   99 - 0x63
    "01100011", -- 2963 - 0xb93  :   99 - 0x63
    "01100011", -- 2964 - 0xb94  :   99 - 0x63
    "01100011", -- 2965 - 0xb95  :   99 - 0x63
    "00111110", -- 2966 - 0xb96  :   62 - 0x3e
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00111110", -- 2968 - 0xb98  :   62 - 0x3e
    "01100011", -- 2969 - 0xb99  :   99 - 0x63
    "01100011", -- 2970 - 0xb9a  :   99 - 0x63
    "01100011", -- 2971 - 0xb9b  :   99 - 0x63
    "01100011", -- 2972 - 0xb9c  :   99 - 0x63
    "01100011", -- 2973 - 0xb9d  :   99 - 0x63
    "00111110", -- 2974 - 0xb9e  :   62 - 0x3e
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "01111110", -- 2976 - 0xba0  :  126 - 0x7e -- Sprite 0xba
    "01100011", -- 2977 - 0xba1  :   99 - 0x63
    "01100011", -- 2978 - 0xba2  :   99 - 0x63
    "01100111", -- 2979 - 0xba3  :  103 - 0x67
    "01111100", -- 2980 - 0xba4  :  124 - 0x7c
    "01101110", -- 2981 - 0xba5  :  110 - 0x6e
    "01100111", -- 2982 - 0xba6  :  103 - 0x67
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "01111110", -- 2984 - 0xba8  :  126 - 0x7e
    "01100011", -- 2985 - 0xba9  :   99 - 0x63
    "01100011", -- 2986 - 0xbaa  :   99 - 0x63
    "01100111", -- 2987 - 0xbab  :  103 - 0x67
    "01111100", -- 2988 - 0xbac  :  124 - 0x7c
    "01101110", -- 2989 - 0xbad  :  110 - 0x6e
    "01100111", -- 2990 - 0xbae  :  103 - 0x67
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "01111111", -- 2992 - 0xbb0  :  127 - 0x7f -- Sprite 0xbb
    "01100000", -- 2993 - 0xbb1  :   96 - 0x60
    "01100000", -- 2994 - 0xbb2  :   96 - 0x60
    "01111110", -- 2995 - 0xbb3  :  126 - 0x7e
    "01100000", -- 2996 - 0xbb4  :   96 - 0x60
    "01100000", -- 2997 - 0xbb5  :   96 - 0x60
    "01111111", -- 2998 - 0xbb6  :  127 - 0x7f
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "01111111", -- 3000 - 0xbb8  :  127 - 0x7f
    "01100000", -- 3001 - 0xbb9  :   96 - 0x60
    "01100000", -- 3002 - 0xbba  :   96 - 0x60
    "01111110", -- 3003 - 0xbbb  :  126 - 0x7e
    "01100000", -- 3004 - 0xbbc  :   96 - 0x60
    "01100000", -- 3005 - 0xbbd  :   96 - 0x60
    "01111111", -- 3006 - 0xbbe  :  127 - 0x7f
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Sprite 0xbc
    "00100010", -- 3009 - 0xbc1  :   34 - 0x22
    "01100101", -- 3010 - 0xbc2  :  101 - 0x65
    "00100101", -- 3011 - 0xbc3  :   37 - 0x25
    "00100101", -- 3012 - 0xbc4  :   37 - 0x25
    "01110010", -- 3013 - 0xbc5  :  114 - 0x72
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Sprite 0xbd
    "01110010", -- 3025 - 0xbd1  :  114 - 0x72
    "01000101", -- 3026 - 0xbd2  :   69 - 0x45
    "01100101", -- 3027 - 0xbd3  :  101 - 0x65
    "00010101", -- 3028 - 0xbd4  :   21 - 0x15
    "01100010", -- 3029 - 0xbd5  :   98 - 0x62
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Sprite 0xbe
    "01100111", -- 3041 - 0xbe1  :  103 - 0x67
    "01010010", -- 3042 - 0xbe2  :   82 - 0x52
    "01100010", -- 3043 - 0xbe3  :   98 - 0x62
    "01000010", -- 3044 - 0xbe4  :   66 - 0x42
    "01000010", -- 3045 - 0xbe5  :   66 - 0x42
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "01100000", -- 3057 - 0xbf1  :   96 - 0x60
    "10000000", -- 3058 - 0xbf2  :  128 - 0x80
    "01000000", -- 3059 - 0xbf3  :   64 - 0x40
    "00100000", -- 3060 - 0xbf4  :   32 - 0x20
    "11000110", -- 3061 - 0xbf5  :  198 - 0xc6
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "01100011", -- 3072 - 0xc00  :   99 - 0x63 -- Sprite 0xc0
    "01100110", -- 3073 - 0xc01  :  102 - 0x66
    "01101100", -- 3074 - 0xc02  :  108 - 0x6c
    "01111000", -- 3075 - 0xc03  :  120 - 0x78
    "01111100", -- 3076 - 0xc04  :  124 - 0x7c
    "01100110", -- 3077 - 0xc05  :  102 - 0x66
    "01100011", -- 3078 - 0xc06  :   99 - 0x63
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "01100011", -- 3080 - 0xc08  :   99 - 0x63
    "01100110", -- 3081 - 0xc09  :  102 - 0x66
    "01101100", -- 3082 - 0xc0a  :  108 - 0x6c
    "01111000", -- 3083 - 0xc0b  :  120 - 0x78
    "01111100", -- 3084 - 0xc0c  :  124 - 0x7c
    "01100110", -- 3085 - 0xc0d  :  102 - 0x66
    "01100011", -- 3086 - 0xc0e  :   99 - 0x63
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00111111", -- 3088 - 0xc10  :   63 - 0x3f -- Sprite 0xc1
    "00001100", -- 3089 - 0xc11  :   12 - 0xc
    "00001100", -- 3090 - 0xc12  :   12 - 0xc
    "00001100", -- 3091 - 0xc13  :   12 - 0xc
    "00001100", -- 3092 - 0xc14  :   12 - 0xc
    "00001100", -- 3093 - 0xc15  :   12 - 0xc
    "00111111", -- 3094 - 0xc16  :   63 - 0x3f
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00111111", -- 3096 - 0xc18  :   63 - 0x3f
    "00001100", -- 3097 - 0xc19  :   12 - 0xc
    "00001100", -- 3098 - 0xc1a  :   12 - 0xc
    "00001100", -- 3099 - 0xc1b  :   12 - 0xc
    "00001100", -- 3100 - 0xc1c  :   12 - 0xc
    "00001100", -- 3101 - 0xc1d  :   12 - 0xc
    "00111111", -- 3102 - 0xc1e  :   63 - 0x3f
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "01100011", -- 3104 - 0xc20  :   99 - 0x63 -- Sprite 0xc2
    "01110111", -- 3105 - 0xc21  :  119 - 0x77
    "01111111", -- 3106 - 0xc22  :  127 - 0x7f
    "01111111", -- 3107 - 0xc23  :  127 - 0x7f
    "01101011", -- 3108 - 0xc24  :  107 - 0x6b
    "01100011", -- 3109 - 0xc25  :   99 - 0x63
    "01100011", -- 3110 - 0xc26  :   99 - 0x63
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "01100011", -- 3112 - 0xc28  :   99 - 0x63
    "01110111", -- 3113 - 0xc29  :  119 - 0x77
    "01111111", -- 3114 - 0xc2a  :  127 - 0x7f
    "01111111", -- 3115 - 0xc2b  :  127 - 0x7f
    "01101011", -- 3116 - 0xc2c  :  107 - 0x6b
    "01100011", -- 3117 - 0xc2d  :   99 - 0x63
    "01100011", -- 3118 - 0xc2e  :   99 - 0x63
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00011100", -- 3120 - 0xc30  :   28 - 0x1c -- Sprite 0xc3
    "00110110", -- 3121 - 0xc31  :   54 - 0x36
    "01100011", -- 3122 - 0xc32  :   99 - 0x63
    "01100011", -- 3123 - 0xc33  :   99 - 0x63
    "01111111", -- 3124 - 0xc34  :  127 - 0x7f
    "01100011", -- 3125 - 0xc35  :   99 - 0x63
    "01100011", -- 3126 - 0xc36  :   99 - 0x63
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00011100", -- 3128 - 0xc38  :   28 - 0x1c
    "00110110", -- 3129 - 0xc39  :   54 - 0x36
    "01100011", -- 3130 - 0xc3a  :   99 - 0x63
    "01100011", -- 3131 - 0xc3b  :   99 - 0x63
    "01111111", -- 3132 - 0xc3c  :  127 - 0x7f
    "01100011", -- 3133 - 0xc3d  :   99 - 0x63
    "01100011", -- 3134 - 0xc3e  :   99 - 0x63
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00011111", -- 3136 - 0xc40  :   31 - 0x1f -- Sprite 0xc4
    "00110000", -- 3137 - 0xc41  :   48 - 0x30
    "01100000", -- 3138 - 0xc42  :   96 - 0x60
    "01100111", -- 3139 - 0xc43  :  103 - 0x67
    "01100011", -- 3140 - 0xc44  :   99 - 0x63
    "00110011", -- 3141 - 0xc45  :   51 - 0x33
    "00011111", -- 3142 - 0xc46  :   31 - 0x1f
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00011111", -- 3144 - 0xc48  :   31 - 0x1f
    "00110000", -- 3145 - 0xc49  :   48 - 0x30
    "01100000", -- 3146 - 0xc4a  :   96 - 0x60
    "01100111", -- 3147 - 0xc4b  :  103 - 0x67
    "01100011", -- 3148 - 0xc4c  :   99 - 0x63
    "00110011", -- 3149 - 0xc4d  :   51 - 0x33
    "00011111", -- 3150 - 0xc4e  :   31 - 0x1f
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "01100011", -- 3152 - 0xc50  :   99 - 0x63 -- Sprite 0xc5
    "01100011", -- 3153 - 0xc51  :   99 - 0x63
    "01100011", -- 3154 - 0xc52  :   99 - 0x63
    "01100011", -- 3155 - 0xc53  :   99 - 0x63
    "01100011", -- 3156 - 0xc54  :   99 - 0x63
    "01100011", -- 3157 - 0xc55  :   99 - 0x63
    "00111110", -- 3158 - 0xc56  :   62 - 0x3e
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "01100011", -- 3160 - 0xc58  :   99 - 0x63
    "01100011", -- 3161 - 0xc59  :   99 - 0x63
    "01100011", -- 3162 - 0xc5a  :   99 - 0x63
    "01100011", -- 3163 - 0xc5b  :   99 - 0x63
    "01100011", -- 3164 - 0xc5c  :   99 - 0x63
    "01100011", -- 3165 - 0xc5d  :   99 - 0x63
    "00111110", -- 3166 - 0xc5e  :   62 - 0x3e
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "01111110", -- 3168 - 0xc60  :  126 - 0x7e -- Sprite 0xc6
    "01100011", -- 3169 - 0xc61  :   99 - 0x63
    "01100011", -- 3170 - 0xc62  :   99 - 0x63
    "01100111", -- 3171 - 0xc63  :  103 - 0x67
    "01111100", -- 3172 - 0xc64  :  124 - 0x7c
    "01101110", -- 3173 - 0xc65  :  110 - 0x6e
    "01100111", -- 3174 - 0xc66  :  103 - 0x67
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "01111110", -- 3176 - 0xc68  :  126 - 0x7e
    "01100011", -- 3177 - 0xc69  :   99 - 0x63
    "01100011", -- 3178 - 0xc6a  :   99 - 0x63
    "01100111", -- 3179 - 0xc6b  :  103 - 0x67
    "01111100", -- 3180 - 0xc6c  :  124 - 0x7c
    "01101110", -- 3181 - 0xc6d  :  110 - 0x6e
    "01100111", -- 3182 - 0xc6e  :  103 - 0x67
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "01111111", -- 3184 - 0xc70  :  127 - 0x7f -- Sprite 0xc7
    "01100000", -- 3185 - 0xc71  :   96 - 0x60
    "01100000", -- 3186 - 0xc72  :   96 - 0x60
    "01111110", -- 3187 - 0xc73  :  126 - 0x7e
    "01100000", -- 3188 - 0xc74  :   96 - 0x60
    "01100000", -- 3189 - 0xc75  :   96 - 0x60
    "01111111", -- 3190 - 0xc76  :  127 - 0x7f
    "00000000", -- 3191 - 0xc77  :    0 - 0x0
    "01111111", -- 3192 - 0xc78  :  127 - 0x7f
    "01100000", -- 3193 - 0xc79  :   96 - 0x60
    "01100000", -- 3194 - 0xc7a  :   96 - 0x60
    "01111110", -- 3195 - 0xc7b  :  126 - 0x7e
    "01100000", -- 3196 - 0xc7c  :   96 - 0x60
    "01100000", -- 3197 - 0xc7d  :   96 - 0x60
    "01111111", -- 3198 - 0xc7e  :  127 - 0x7f
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00110110", -- 3200 - 0xc80  :   54 - 0x36 -- Sprite 0xc8
    "00110110", -- 3201 - 0xc81  :   54 - 0x36
    "00010010", -- 3202 - 0xc82  :   18 - 0x12
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00110110", -- 3208 - 0xc88  :   54 - 0x36
    "00110110", -- 3209 - 0xc89  :   54 - 0x36
    "00010010", -- 3210 - 0xc8a  :   18 - 0x12
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00111110", -- 3216 - 0xc90  :   62 - 0x3e -- Sprite 0xc9
    "01100011", -- 3217 - 0xc91  :   99 - 0x63
    "01100011", -- 3218 - 0xc92  :   99 - 0x63
    "01100011", -- 3219 - 0xc93  :   99 - 0x63
    "01100011", -- 3220 - 0xc94  :   99 - 0x63
    "01100011", -- 3221 - 0xc95  :   99 - 0x63
    "00111110", -- 3222 - 0xc96  :   62 - 0x3e
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00111110", -- 3224 - 0xc98  :   62 - 0x3e
    "01100011", -- 3225 - 0xc99  :   99 - 0x63
    "01100011", -- 3226 - 0xc9a  :   99 - 0x63
    "01100011", -- 3227 - 0xc9b  :   99 - 0x63
    "01100011", -- 3228 - 0xc9c  :   99 - 0x63
    "01100011", -- 3229 - 0xc9d  :   99 - 0x63
    "00111110", -- 3230 - 0xc9e  :   62 - 0x3e
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00111100", -- 3232 - 0xca0  :   60 - 0x3c -- Sprite 0xca
    "01100110", -- 3233 - 0xca1  :  102 - 0x66
    "01100000", -- 3234 - 0xca2  :   96 - 0x60
    "00111110", -- 3235 - 0xca3  :   62 - 0x3e
    "00000011", -- 3236 - 0xca4  :    3 - 0x3
    "01100011", -- 3237 - 0xca5  :   99 - 0x63
    "00111110", -- 3238 - 0xca6  :   62 - 0x3e
    "00000000", -- 3239 - 0xca7  :    0 - 0x0
    "00111100", -- 3240 - 0xca8  :   60 - 0x3c
    "01100110", -- 3241 - 0xca9  :  102 - 0x66
    "01100000", -- 3242 - 0xcaa  :   96 - 0x60
    "00111110", -- 3243 - 0xcab  :   62 - 0x3e
    "00000011", -- 3244 - 0xcac  :    3 - 0x3
    "01100011", -- 3245 - 0xcad  :   99 - 0x63
    "00111110", -- 3246 - 0xcae  :   62 - 0x3e
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00000000", -- 3250 - 0xcb2  :    0 - 0x0
    "00000000", -- 3251 - 0xcb3  :    0 - 0x0
    "00000000", -- 3252 - 0xcb4  :    0 - 0x0
    "00000000", -- 3253 - 0xcb5  :    0 - 0x0
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0
    "00111000", -- 3257 - 0xcb9  :   56 - 0x38
    "01111100", -- 3258 - 0xcba  :  124 - 0x7c
    "11111110", -- 3259 - 0xcbb  :  254 - 0xfe
    "11111110", -- 3260 - 0xcbc  :  254 - 0xfe
    "11111110", -- 3261 - 0xcbd  :  254 - 0xfe
    "01111100", -- 3262 - 0xcbe  :  124 - 0x7c
    "00111000", -- 3263 - 0xcbf  :   56 - 0x38
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000000", -- 3268 - 0xcc4  :    0 - 0x0
    "00000000", -- 3269 - 0xcc5  :    0 - 0x0
    "00000000", -- 3270 - 0xcc6  :    0 - 0x0
    "00000000", -- 3271 - 0xcc7  :    0 - 0x0
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "00000000", -- 3277 - 0xccd  :    0 - 0x0
    "00000000", -- 3278 - 0xcce  :    0 - 0x0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00000000", -- 3284 - 0xcd4  :    0 - 0x0
    "00000000", -- 3285 - 0xcd5  :    0 - 0x0
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000000", -- 3300 - 0xce4  :    0 - 0x0
    "00000000", -- 3301 - 0xce5  :    0 - 0x0
    "00000000", -- 3302 - 0xce6  :    0 - 0x0
    "00000000", -- 3303 - 0xce7  :    0 - 0x0
    "00000000", -- 3304 - 0xce8  :    0 - 0x0
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00000000", -- 3308 - 0xcec  :    0 - 0x0
    "00000000", -- 3309 - 0xced  :    0 - 0x0
    "00000000", -- 3310 - 0xcee  :    0 - 0x0
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00000000", -- 3315 - 0xcf3  :    0 - 0x0
    "00000000", -- 3316 - 0xcf4  :    0 - 0x0
    "00000000", -- 3317 - 0xcf5  :    0 - 0x0
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00000000", -- 3324 - 0xcfc  :    0 - 0x0
    "00000000", -- 3325 - 0xcfd  :    0 - 0x0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "01000111", -- 3328 - 0xd00  :   71 - 0x47 -- Sprite 0xd0
    "01000111", -- 3329 - 0xd01  :   71 - 0x47
    "00001111", -- 3330 - 0xd02  :   15 - 0xf
    "00001111", -- 3331 - 0xd03  :   15 - 0xf
    "00011111", -- 3332 - 0xd04  :   31 - 0x1f
    "00011111", -- 3333 - 0xd05  :   31 - 0x1f
    "00111111", -- 3334 - 0xd06  :   63 - 0x3f
    "00111111", -- 3335 - 0xd07  :   63 - 0x3f
    "00010111", -- 3336 - 0xd08  :   23 - 0x17
    "00010111", -- 3337 - 0xd09  :   23 - 0x17
    "00101111", -- 3338 - 0xd0a  :   47 - 0x2f
    "00101111", -- 3339 - 0xd0b  :   47 - 0x2f
    "01011111", -- 3340 - 0xd0c  :   95 - 0x5f
    "01011111", -- 3341 - 0xd0d  :   95 - 0x5f
    "00111111", -- 3342 - 0xd0e  :   63 - 0x3f
    "00111111", -- 3343 - 0xd0f  :   63 - 0x3f
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Sprite 0xd1
    "11001111", -- 3345 - 0xd11  :  207 - 0xcf
    "11001111", -- 3346 - 0xd12  :  207 - 0xcf
    "11111011", -- 3347 - 0xd13  :  251 - 0xfb
    "11110111", -- 3348 - 0xd14  :  247 - 0xf7
    "11100111", -- 3349 - 0xd15  :  231 - 0xe7
    "11111111", -- 3350 - 0xd16  :  255 - 0xff
    "11111111", -- 3351 - 0xd17  :  255 - 0xff
    "11111111", -- 3352 - 0xd18  :  255 - 0xff
    "11001111", -- 3353 - 0xd19  :  207 - 0xcf
    "11001111", -- 3354 - 0xd1a  :  207 - 0xcf
    "11111011", -- 3355 - 0xd1b  :  251 - 0xfb
    "11110111", -- 3356 - 0xd1c  :  247 - 0xf7
    "11100111", -- 3357 - 0xd1d  :  231 - 0xe7
    "11111111", -- 3358 - 0xd1e  :  255 - 0xff
    "11111111", -- 3359 - 0xd1f  :  255 - 0xff
    "00011000", -- 3360 - 0xd20  :   24 - 0x18 -- Sprite 0xd2
    "00001000", -- 3361 - 0xd21  :    8 - 0x8
    "10001000", -- 3362 - 0xd22  :  136 - 0x88
    "10000000", -- 3363 - 0xd23  :  128 - 0x80
    "01000000", -- 3364 - 0xd24  :   64 - 0x40
    "01000000", -- 3365 - 0xd25  :   64 - 0x40
    "10100000", -- 3366 - 0xd26  :  160 - 0xa0
    "10100000", -- 3367 - 0xd27  :  160 - 0xa0
    "01000010", -- 3368 - 0xd28  :   66 - 0x42
    "01100010", -- 3369 - 0xd29  :   98 - 0x62
    "10100010", -- 3370 - 0xd2a  :  162 - 0xa2
    "10110010", -- 3371 - 0xd2b  :  178 - 0xb2
    "01010010", -- 3372 - 0xd2c  :   82 - 0x52
    "01011010", -- 3373 - 0xd2d  :   90 - 0x5a
    "10101010", -- 3374 - 0xd2e  :  170 - 0xaa
    "10101100", -- 3375 - 0xd2f  :  172 - 0xac
    "11111111", -- 3376 - 0xd30  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11111101", -- 3380 - 0xd34  :  253 - 0xfd
    "11111101", -- 3381 - 0xd35  :  253 - 0xfd
    "11111101", -- 3382 - 0xd36  :  253 - 0xfd
    "11111101", -- 3383 - 0xd37  :  253 - 0xfd
    "11111111", -- 3384 - 0xd38  :  255 - 0xff
    "11111111", -- 3385 - 0xd39  :  255 - 0xff
    "11111111", -- 3386 - 0xd3a  :  255 - 0xff
    "11111111", -- 3387 - 0xd3b  :  255 - 0xff
    "11111101", -- 3388 - 0xd3c  :  253 - 0xfd
    "11111101", -- 3389 - 0xd3d  :  253 - 0xfd
    "11111101", -- 3390 - 0xd3e  :  253 - 0xfd
    "11111101", -- 3391 - 0xd3f  :  253 - 0xfd
    "11000111", -- 3392 - 0xd40  :  199 - 0xc7 -- Sprite 0xd4
    "11110111", -- 3393 - 0xd41  :  247 - 0xf7
    "11110000", -- 3394 - 0xd42  :  240 - 0xf0
    "11111000", -- 3395 - 0xd43  :  248 - 0xf8
    "11111000", -- 3396 - 0xd44  :  248 - 0xf8
    "11111111", -- 3397 - 0xd45  :  255 - 0xff
    "11111111", -- 3398 - 0xd46  :  255 - 0xff
    "11111111", -- 3399 - 0xd47  :  255 - 0xff
    "00000111", -- 3400 - 0xd48  :    7 - 0x7
    "00000111", -- 3401 - 0xd49  :    7 - 0x7
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000011", -- 3403 - 0xd4b  :    3 - 0x3
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "11111000", -- 3408 - 0xd50  :  248 - 0xf8 -- Sprite 0xd5
    "11111000", -- 3409 - 0xd51  :  248 - 0xf8
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "11111111", -- 3413 - 0xd55  :  255 - 0xff
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "11111010", -- 3416 - 0xd58  :  250 - 0xfa
    "11111010", -- 3417 - 0xd59  :  250 - 0xfa
    "00000010", -- 3418 - 0xd5a  :    2 - 0x2
    "11111110", -- 3419 - 0xd5b  :  254 - 0xfe
    "00000000", -- 3420 - 0xd5c  :    0 - 0x0
    "00000000", -- 3421 - 0xd5d  :    0 - 0x0
    "00000000", -- 3422 - 0xd5e  :    0 - 0x0
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "10001111", -- 3424 - 0xd60  :  143 - 0x8f -- Sprite 0xd6
    "11101111", -- 3425 - 0xd61  :  239 - 0xef
    "11000000", -- 3426 - 0xd62  :  192 - 0xc0
    "11110000", -- 3427 - 0xd63  :  240 - 0xf0
    "11100000", -- 3428 - 0xd64  :  224 - 0xe0
    "11111111", -- 3429 - 0xd65  :  255 - 0xff
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "00001111", -- 3432 - 0xd68  :   15 - 0xf
    "00001111", -- 3433 - 0xd69  :   15 - 0xf
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "00000111", -- 3435 - 0xd6b  :    7 - 0x7
    "00000000", -- 3436 - 0xd6c  :    0 - 0x0
    "00000000", -- 3437 - 0xd6d  :    0 - 0x0
    "00000000", -- 3438 - 0xd6e  :    0 - 0x0
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "11111111", -- 3440 - 0xd70  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "00000000", -- 3442 - 0xd72  :    0 - 0x0
    "00000000", -- 3443 - 0xd73  :    0 - 0x0
    "00000000", -- 3444 - 0xd74  :    0 - 0x0
    "11111111", -- 3445 - 0xd75  :  255 - 0xff
    "11111111", -- 3446 - 0xd76  :  255 - 0xff
    "11111111", -- 3447 - 0xd77  :  255 - 0xff
    "11111111", -- 3448 - 0xd78  :  255 - 0xff
    "11111111", -- 3449 - 0xd79  :  255 - 0xff
    "00000000", -- 3450 - 0xd7a  :    0 - 0x0
    "11111111", -- 3451 - 0xd7b  :  255 - 0xff
    "00000000", -- 3452 - 0xd7c  :    0 - 0x0
    "00000000", -- 3453 - 0xd7d  :    0 - 0x0
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "11000011", -- 3456 - 0xd80  :  195 - 0xc3 -- Sprite 0xd8
    "11111111", -- 3457 - 0xd81  :  255 - 0xff
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000000", -- 3460 - 0xd84  :    0 - 0x0
    "11111111", -- 3461 - 0xd85  :  255 - 0xff
    "11111111", -- 3462 - 0xd86  :  255 - 0xff
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11000011", -- 3464 - 0xd88  :  195 - 0xc3
    "11111111", -- 3465 - 0xd89  :  255 - 0xff
    "00000000", -- 3466 - 0xd8a  :    0 - 0x0
    "11111111", -- 3467 - 0xd8b  :  255 - 0xff
    "00000000", -- 3468 - 0xd8c  :    0 - 0x0
    "00000000", -- 3469 - 0xd8d  :    0 - 0x0
    "00000000", -- 3470 - 0xd8e  :    0 - 0x0
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00000011", -- 3472 - 0xd90  :    3 - 0x3 -- Sprite 0xd9
    "10000001", -- 3473 - 0xd91  :  129 - 0x81
    "00000000", -- 3474 - 0xd92  :    0 - 0x0
    "00000000", -- 3475 - 0xd93  :    0 - 0x0
    "00000011", -- 3476 - 0xd94  :    3 - 0x3
    "11111111", -- 3477 - 0xd95  :  255 - 0xff
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111111", -- 3479 - 0xd97  :  255 - 0xff
    "01101011", -- 3480 - 0xd98  :  107 - 0x6b
    "10110101", -- 3481 - 0xd99  :  181 - 0xb5
    "00110110", -- 3482 - 0xd9a  :   54 - 0x36
    "11111000", -- 3483 - 0xd9b  :  248 - 0xf8
    "00000000", -- 3484 - 0xd9c  :    0 - 0x0
    "00000000", -- 3485 - 0xd9d  :    0 - 0x0
    "00000000", -- 3486 - 0xd9e  :    0 - 0x0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "11111111", -- 3488 - 0xda0  :  255 - 0xff -- Sprite 0xda
    "11111111", -- 3489 - 0xda1  :  255 - 0xff
    "01111110", -- 3490 - 0xda2  :  126 - 0x7e
    "00000000", -- 3491 - 0xda3  :    0 - 0x0
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "11100000", -- 3493 - 0xda5  :  224 - 0xe0
    "11111111", -- 3494 - 0xda6  :  255 - 0xff
    "11111111", -- 3495 - 0xda7  :  255 - 0xff
    "11111111", -- 3496 - 0xda8  :  255 - 0xff
    "11111111", -- 3497 - 0xda9  :  255 - 0xff
    "01111110", -- 3498 - 0xdaa  :  126 - 0x7e
    "10000001", -- 3499 - 0xdab  :  129 - 0x81
    "00011111", -- 3500 - 0xdac  :   31 - 0x1f
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "01100001", -- 3504 - 0xdb0  :   97 - 0x61 -- Sprite 0xdb
    "11000011", -- 3505 - 0xdb1  :  195 - 0xc3
    "00000111", -- 3506 - 0xdb2  :    7 - 0x7
    "00001111", -- 3507 - 0xdb3  :   15 - 0xf
    "00011111", -- 3508 - 0xdb4  :   31 - 0x1f
    "01111111", -- 3509 - 0xdb5  :  127 - 0x7f
    "11111111", -- 3510 - 0xdb6  :  255 - 0xff
    "11111111", -- 3511 - 0xdb7  :  255 - 0xff
    "01101100", -- 3512 - 0xdb8  :  108 - 0x6c
    "11011000", -- 3513 - 0xdb9  :  216 - 0xd8
    "00110000", -- 3514 - 0xdba  :   48 - 0x30
    "11100000", -- 3515 - 0xdbb  :  224 - 0xe0
    "10000000", -- 3516 - 0xdbc  :  128 - 0x80
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000000", -- 3518 - 0xdbe  :    0 - 0x0
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00011111", -- 3520 - 0xdc0  :   31 - 0x1f -- Sprite 0xdc
    "11011111", -- 3521 - 0xdc1  :  223 - 0xdf
    "11000000", -- 3522 - 0xdc2  :  192 - 0xc0
    "11110000", -- 3523 - 0xdc3  :  240 - 0xf0
    "11110000", -- 3524 - 0xdc4  :  240 - 0xf0
    "11111111", -- 3525 - 0xdc5  :  255 - 0xff
    "11111111", -- 3526 - 0xdc6  :  255 - 0xff
    "11111111", -- 3527 - 0xdc7  :  255 - 0xff
    "00011111", -- 3528 - 0xdc8  :   31 - 0x1f
    "00011111", -- 3529 - 0xdc9  :   31 - 0x1f
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000111", -- 3531 - 0xdcb  :    7 - 0x7
    "00000000", -- 3532 - 0xdcc  :    0 - 0x0
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "00000000", -- 3534 - 0xdce  :    0 - 0x0
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "10000100", -- 3536 - 0xdd0  :  132 - 0x84 -- Sprite 0xdd
    "11111100", -- 3537 - 0xdd1  :  252 - 0xfc
    "00000000", -- 3538 - 0xdd2  :    0 - 0x0
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "11111111", -- 3541 - 0xdd5  :  255 - 0xff
    "11111111", -- 3542 - 0xdd6  :  255 - 0xff
    "11111111", -- 3543 - 0xdd7  :  255 - 0xff
    "10000101", -- 3544 - 0xdd8  :  133 - 0x85
    "11111101", -- 3545 - 0xdd9  :  253 - 0xfd
    "00000001", -- 3546 - 0xdda  :    1 - 0x1
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000000", -- 3550 - 0xdde  :    0 - 0x0
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "01111111", -- 3552 - 0xde0  :  127 - 0x7f -- Sprite 0xde
    "01111111", -- 3553 - 0xde1  :  127 - 0x7f
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "11111111", -- 3557 - 0xde5  :  255 - 0xff
    "11111111", -- 3558 - 0xde6  :  255 - 0xff
    "11111111", -- 3559 - 0xde7  :  255 - 0xff
    "01111111", -- 3560 - 0xde8  :  127 - 0x7f
    "01111111", -- 3561 - 0xde9  :  127 - 0x7f
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "01011111", -- 3563 - 0xdeb  :   95 - 0x5f
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "11111100", -- 3568 - 0xdf0  :  252 - 0xfc -- Sprite 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111111", -- 3575 - 0xdf7  :  255 - 0xff
    "11111100", -- 3576 - 0xdf8  :  252 - 0xfc
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00110000", -- 3584 - 0xe00  :   48 - 0x30 -- Sprite 0xe0
    "11110000", -- 3585 - 0xe01  :  240 - 0xf0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "11111111", -- 3589 - 0xe05  :  255 - 0xff
    "11111111", -- 3590 - 0xe06  :  255 - 0xff
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "00110100", -- 3592 - 0xe08  :   52 - 0x34
    "11110110", -- 3593 - 0xe09  :  246 - 0xf6
    "00000010", -- 3594 - 0xe0a  :    2 - 0x2
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "11111111", -- 3600 - 0xe10  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "11111111", -- 3605 - 0xe15  :  255 - 0xff
    "11111111", -- 3606 - 0xe16  :  255 - 0xff
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "11111111", -- 3608 - 0xe18  :  255 - 0xff
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "01111111", -- 3611 - 0xe1b  :  127 - 0x7f
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "11100001", -- 3616 - 0xe20  :  225 - 0xe1 -- Sprite 0xe2
    "11111111", -- 3617 - 0xe21  :  255 - 0xff
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "11111111", -- 3621 - 0xe25  :  255 - 0xff
    "11111111", -- 3622 - 0xe26  :  255 - 0xff
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11100001", -- 3624 - 0xe28  :  225 - 0xe1
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00011111", -- 3632 - 0xe30  :   31 - 0x1f -- Sprite 0xe3
    "00011111", -- 3633 - 0xe31  :   31 - 0x1f
    "00011111", -- 3634 - 0xe32  :   31 - 0x1f
    "00011111", -- 3635 - 0xe33  :   31 - 0x1f
    "00011111", -- 3636 - 0xe34  :   31 - 0x1f
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "01000000", -- 3640 - 0xe38  :   64 - 0x40
    "01000000", -- 3641 - 0xe39  :   64 - 0x40
    "01000000", -- 3642 - 0xe3a  :   64 - 0x40
    "11000000", -- 3643 - 0xe3b  :  192 - 0xc0
    "00000000", -- 3644 - 0xe3c  :    0 - 0x0
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Sprite 0xe4
    "00011111", -- 3649 - 0xe41  :   31 - 0x1f
    "00111111", -- 3650 - 0xe42  :   63 - 0x3f
    "01111000", -- 3651 - 0xe43  :  120 - 0x78
    "01110111", -- 3652 - 0xe44  :  119 - 0x77
    "01101111", -- 3653 - 0xe45  :  111 - 0x6f
    "01101111", -- 3654 - 0xe46  :  111 - 0x6f
    "01101111", -- 3655 - 0xe47  :  111 - 0x6f
    "00000000", -- 3656 - 0xe48  :    0 - 0x0
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000111", -- 3660 - 0xe4c  :    7 - 0x7
    "00001111", -- 3661 - 0xe4d  :   15 - 0xf
    "00001111", -- 3662 - 0xe4e  :   15 - 0xf
    "00001111", -- 3663 - 0xe4f  :   15 - 0xf
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Sprite 0xe5
    "11111000", -- 3665 - 0xe51  :  248 - 0xf8
    "11111100", -- 3666 - 0xe52  :  252 - 0xfc
    "00011110", -- 3667 - 0xe53  :   30 - 0x1e
    "11101110", -- 3668 - 0xe54  :  238 - 0xee
    "11110110", -- 3669 - 0xe55  :  246 - 0xf6
    "11110110", -- 3670 - 0xe56  :  246 - 0xf6
    "11110110", -- 3671 - 0xe57  :  246 - 0xf6
    "00000000", -- 3672 - 0xe58  :    0 - 0x0
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "11100000", -- 3676 - 0xe5c  :  224 - 0xe0
    "11110000", -- 3677 - 0xe5d  :  240 - 0xf0
    "11110000", -- 3678 - 0xe5e  :  240 - 0xf0
    "11110000", -- 3679 - 0xe5f  :  240 - 0xf0
    "11110110", -- 3680 - 0xe60  :  246 - 0xf6 -- Sprite 0xe6
    "11110110", -- 3681 - 0xe61  :  246 - 0xf6
    "11110110", -- 3682 - 0xe62  :  246 - 0xf6
    "11101110", -- 3683 - 0xe63  :  238 - 0xee
    "00011110", -- 3684 - 0xe64  :   30 - 0x1e
    "11111100", -- 3685 - 0xe65  :  252 - 0xfc
    "11111000", -- 3686 - 0xe66  :  248 - 0xf8
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "11110000", -- 3688 - 0xe68  :  240 - 0xf0
    "11110000", -- 3689 - 0xe69  :  240 - 0xf0
    "11110000", -- 3690 - 0xe6a  :  240 - 0xf0
    "11100000", -- 3691 - 0xe6b  :  224 - 0xe0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "01101111", -- 3696 - 0xe70  :  111 - 0x6f -- Sprite 0xe7
    "01101111", -- 3697 - 0xe71  :  111 - 0x6f
    "01101111", -- 3698 - 0xe72  :  111 - 0x6f
    "01110111", -- 3699 - 0xe73  :  119 - 0x77
    "01111000", -- 3700 - 0xe74  :  120 - 0x78
    "00111111", -- 3701 - 0xe75  :   63 - 0x3f
    "00011111", -- 3702 - 0xe76  :   31 - 0x1f
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00001111", -- 3704 - 0xe78  :   15 - 0xf
    "00001111", -- 3705 - 0xe79  :   15 - 0xf
    "00001111", -- 3706 - 0xe7a  :   15 - 0xf
    "00000111", -- 3707 - 0xe7b  :    7 - 0x7
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Sprite 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "00000000", -- 3720 - 0xe88  :    0 - 0x0
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11110110", -- 3728 - 0xe90  :  246 - 0xf6 -- Sprite 0xe9
    "11110110", -- 3729 - 0xe91  :  246 - 0xf6
    "11110110", -- 3730 - 0xe92  :  246 - 0xf6
    "11110110", -- 3731 - 0xe93  :  246 - 0xf6
    "11110110", -- 3732 - 0xe94  :  246 - 0xf6
    "11110110", -- 3733 - 0xe95  :  246 - 0xf6
    "11110110", -- 3734 - 0xe96  :  246 - 0xf6
    "11110110", -- 3735 - 0xe97  :  246 - 0xf6
    "11110000", -- 3736 - 0xe98  :  240 - 0xf0
    "11110000", -- 3737 - 0xe99  :  240 - 0xf0
    "11110000", -- 3738 - 0xe9a  :  240 - 0xf0
    "11110000", -- 3739 - 0xe9b  :  240 - 0xf0
    "11110000", -- 3740 - 0xe9c  :  240 - 0xf0
    "11110000", -- 3741 - 0xe9d  :  240 - 0xf0
    "11110000", -- 3742 - 0xe9e  :  240 - 0xf0
    "11110000", -- 3743 - 0xe9f  :  240 - 0xf0
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "11111111", -- 3752 - 0xea8  :  255 - 0xff
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "01101111", -- 3760 - 0xeb0  :  111 - 0x6f -- Sprite 0xeb
    "01101111", -- 3761 - 0xeb1  :  111 - 0x6f
    "01101111", -- 3762 - 0xeb2  :  111 - 0x6f
    "01101111", -- 3763 - 0xeb3  :  111 - 0x6f
    "01101111", -- 3764 - 0xeb4  :  111 - 0x6f
    "01101111", -- 3765 - 0xeb5  :  111 - 0x6f
    "01101111", -- 3766 - 0xeb6  :  111 - 0x6f
    "01101111", -- 3767 - 0xeb7  :  111 - 0x6f
    "00001111", -- 3768 - 0xeb8  :   15 - 0xf
    "00001111", -- 3769 - 0xeb9  :   15 - 0xf
    "00001111", -- 3770 - 0xeba  :   15 - 0xf
    "00001111", -- 3771 - 0xebb  :   15 - 0xf
    "00001111", -- 3772 - 0xebc  :   15 - 0xf
    "00001111", -- 3773 - 0xebd  :   15 - 0xf
    "00001111", -- 3774 - 0xebe  :   15 - 0xf
    "00001111", -- 3775 - 0xebf  :   15 - 0xf
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0
    "00000000", -- 3801 - 0xed9  :    0 - 0x0
    "00000000", -- 3802 - 0xeda  :    0 - 0x0
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000000", -- 3816 - 0xee8  :    0 - 0x0
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "00000000", -- 3828 - 0xef4  :    0 - 0x0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "00000000", -- 3830 - 0xef6  :    0 - 0x0
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "00000000", -- 3832 - 0xef8  :    0 - 0x0
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "11111111", -- 3840 - 0xf00  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 3841 - 0xf01  :  255 - 0xff
    "11111111", -- 3842 - 0xf02  :  255 - 0xff
    "11111111", -- 3843 - 0xf03  :  255 - 0xff
    "11111111", -- 3844 - 0xf04  :  255 - 0xff
    "11111111", -- 3845 - 0xf05  :  255 - 0xff
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11111111", -- 3848 - 0xf08  :  255 - 0xff
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "11111111", -- 3850 - 0xf0a  :  255 - 0xff
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "11111111", -- 3860 - 0xf14  :  255 - 0xff
    "11111111", -- 3861 - 0xf15  :  255 - 0xff
    "11111111", -- 3862 - 0xf16  :  255 - 0xff
    "11111111", -- 3863 - 0xf17  :  255 - 0xff
    "11111111", -- 3864 - 0xf18  :  255 - 0xff
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11111111", -- 3867 - 0xf1b  :  255 - 0xff
    "11111111", -- 3868 - 0xf1c  :  255 - 0xff
    "11111111", -- 3869 - 0xf1d  :  255 - 0xff
    "11111111", -- 3870 - 0xf1e  :  255 - 0xff
    "11111111", -- 3871 - 0xf1f  :  255 - 0xff
    "11111111", -- 3872 - 0xf20  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 3873 - 0xf21  :  255 - 0xff
    "11111111", -- 3874 - 0xf22  :  255 - 0xff
    "11111111", -- 3875 - 0xf23  :  255 - 0xff
    "11111111", -- 3876 - 0xf24  :  255 - 0xff
    "11111111", -- 3877 - 0xf25  :  255 - 0xff
    "11111111", -- 3878 - 0xf26  :  255 - 0xff
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11111111", -- 3883 - 0xf2b  :  255 - 0xff
    "11111111", -- 3884 - 0xf2c  :  255 - 0xff
    "11111111", -- 3885 - 0xf2d  :  255 - 0xff
    "11111111", -- 3886 - 0xf2e  :  255 - 0xff
    "11111111", -- 3887 - 0xf2f  :  255 - 0xff
    "11111111", -- 3888 - 0xf30  :  255 - 0xff -- Sprite 0xf3
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "11111111", -- 3891 - 0xf33  :  255 - 0xff
    "11111111", -- 3892 - 0xf34  :  255 - 0xff
    "11111111", -- 3893 - 0xf35  :  255 - 0xff
    "11111111", -- 3894 - 0xf36  :  255 - 0xff
    "11111111", -- 3895 - 0xf37  :  255 - 0xff
    "11111111", -- 3896 - 0xf38  :  255 - 0xff
    "11111111", -- 3897 - 0xf39  :  255 - 0xff
    "11111111", -- 3898 - 0xf3a  :  255 - 0xff
    "11111111", -- 3899 - 0xf3b  :  255 - 0xff
    "11111111", -- 3900 - 0xf3c  :  255 - 0xff
    "11111111", -- 3901 - 0xf3d  :  255 - 0xff
    "11111111", -- 3902 - 0xf3e  :  255 - 0xff
    "11111111", -- 3903 - 0xf3f  :  255 - 0xff
    "11111111", -- 3904 - 0xf40  :  255 - 0xff -- Sprite 0xf4
    "11111111", -- 3905 - 0xf41  :  255 - 0xff
    "11111111", -- 3906 - 0xf42  :  255 - 0xff
    "11111111", -- 3907 - 0xf43  :  255 - 0xff
    "11111111", -- 3908 - 0xf44  :  255 - 0xff
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "11111111", -- 3912 - 0xf48  :  255 - 0xff
    "11111111", -- 3913 - 0xf49  :  255 - 0xff
    "11111111", -- 3914 - 0xf4a  :  255 - 0xff
    "11111111", -- 3915 - 0xf4b  :  255 - 0xff
    "11111111", -- 3916 - 0xf4c  :  255 - 0xff
    "11111111", -- 3917 - 0xf4d  :  255 - 0xff
    "11111111", -- 3918 - 0xf4e  :  255 - 0xff
    "11111111", -- 3919 - 0xf4f  :  255 - 0xff
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Sprite 0xf5
    "11111111", -- 3921 - 0xf51  :  255 - 0xff
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "11111111", -- 3923 - 0xf53  :  255 - 0xff
    "11111111", -- 3924 - 0xf54  :  255 - 0xff
    "11111111", -- 3925 - 0xf55  :  255 - 0xff
    "11111111", -- 3926 - 0xf56  :  255 - 0xff
    "11111111", -- 3927 - 0xf57  :  255 - 0xff
    "11111111", -- 3928 - 0xf58  :  255 - 0xff
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "11111111", -- 3931 - 0xf5b  :  255 - 0xff
    "11111111", -- 3932 - 0xf5c  :  255 - 0xff
    "11111111", -- 3933 - 0xf5d  :  255 - 0xff
    "11111111", -- 3934 - 0xf5e  :  255 - 0xff
    "11111111", -- 3935 - 0xf5f  :  255 - 0xff
    "11111111", -- 3936 - 0xf60  :  255 - 0xff -- Sprite 0xf6
    "11111111", -- 3937 - 0xf61  :  255 - 0xff
    "11111111", -- 3938 - 0xf62  :  255 - 0xff
    "11111111", -- 3939 - 0xf63  :  255 - 0xff
    "11111111", -- 3940 - 0xf64  :  255 - 0xff
    "11111111", -- 3941 - 0xf65  :  255 - 0xff
    "11111111", -- 3942 - 0xf66  :  255 - 0xff
    "11111111", -- 3943 - 0xf67  :  255 - 0xff
    "11111111", -- 3944 - 0xf68  :  255 - 0xff
    "11111111", -- 3945 - 0xf69  :  255 - 0xff
    "11111111", -- 3946 - 0xf6a  :  255 - 0xff
    "11111111", -- 3947 - 0xf6b  :  255 - 0xff
    "11111111", -- 3948 - 0xf6c  :  255 - 0xff
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "11111111", -- 3952 - 0xf70  :  255 - 0xff -- Sprite 0xf7
    "11111111", -- 3953 - 0xf71  :  255 - 0xff
    "11111111", -- 3954 - 0xf72  :  255 - 0xff
    "11111111", -- 3955 - 0xf73  :  255 - 0xff
    "11111111", -- 3956 - 0xf74  :  255 - 0xff
    "11111111", -- 3957 - 0xf75  :  255 - 0xff
    "11111111", -- 3958 - 0xf76  :  255 - 0xff
    "11111111", -- 3959 - 0xf77  :  255 - 0xff
    "11111111", -- 3960 - 0xf78  :  255 - 0xff
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "11111111", -- 3968 - 0xf80  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "11111111", -- 3970 - 0xf82  :  255 - 0xff
    "11111111", -- 3971 - 0xf83  :  255 - 0xff
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "11111111", -- 3974 - 0xf86  :  255 - 0xff
    "11111111", -- 3975 - 0xf87  :  255 - 0xff
    "11111111", -- 3976 - 0xf88  :  255 - 0xff
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111111", -- 3982 - 0xf8e  :  255 - 0xff
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "11111111", -- 3992 - 0xf98  :  255 - 0xff
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111111", -- 3999 - 0xf9f  :  255 - 0xff
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "11111111", -- 4007 - 0xfa7  :  255 - 0xff
    "11111111", -- 4008 - 0xfa8  :  255 - 0xff
    "11111111", -- 4009 - 0xfa9  :  255 - 0xff
    "11111111", -- 4010 - 0xfaa  :  255 - 0xff
    "11111111", -- 4011 - 0xfab  :  255 - 0xff
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "11111111", -- 4015 - 0xfaf  :  255 - 0xff
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "11111111", -- 4024 - 0xfb8  :  255 - 0xff
    "11111111", -- 4025 - 0xfb9  :  255 - 0xff
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "11111111", -- 4031 - 0xfbf  :  255 - 0xff
    "11111111", -- 4032 - 0xfc0  :  255 - 0xff -- Sprite 0xfc
    "11111111", -- 4033 - 0xfc1  :  255 - 0xff
    "11111111", -- 4034 - 0xfc2  :  255 - 0xff
    "11111111", -- 4035 - 0xfc3  :  255 - 0xff
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "11111111", -- 4040 - 0xfc8  :  255 - 0xff
    "11111111", -- 4041 - 0xfc9  :  255 - 0xff
    "11111111", -- 4042 - 0xfca  :  255 - 0xff
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "11111111", -- 4048 - 0xfd0  :  255 - 0xff -- Sprite 0xfd
    "11111111", -- 4049 - 0xfd1  :  255 - 0xff
    "11111111", -- 4050 - 0xfd2  :  255 - 0xff
    "11111111", -- 4051 - 0xfd3  :  255 - 0xff
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "11111111", -- 4064 - 0xfe0  :  255 - 0xff -- Sprite 0xfe
    "11111111", -- 4065 - 0xfe1  :  255 - 0xff
    "11111111", -- 4066 - 0xfe2  :  255 - 0xff
    "11111111", -- 4067 - 0xfe3  :  255 - 0xff
    "11111111", -- 4068 - 0xfe4  :  255 - 0xff
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11111111", -- 4075 - 0xfeb  :  255 - 0xff
    "11111111", -- 4076 - 0xfec  :  255 - 0xff
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111", -- 4095 - 0xfff  :  255 - 0xff
          -- Pattern Table 1---------
    "00000000", -- 4096 - 0x1000  :    0 - 0x0 -- Background 0x0
    "00000011", -- 4097 - 0x1001  :    3 - 0x3
    "00001111", -- 4098 - 0x1002  :   15 - 0xf
    "00011111", -- 4099 - 0x1003  :   31 - 0x1f
    "00111111", -- 4100 - 0x1004  :   63 - 0x3f
    "00111111", -- 4101 - 0x1005  :   63 - 0x3f
    "01111111", -- 4102 - 0x1006  :  127 - 0x7f
    "01111111", -- 4103 - 0x1007  :  127 - 0x7f
    "00000000", -- 4104 - 0x1008  :    0 - 0x0
    "00000000", -- 4105 - 0x1009  :    0 - 0x0
    "00000000", -- 4106 - 0x100a  :    0 - 0x0
    "00000000", -- 4107 - 0x100b  :    0 - 0x0
    "00000000", -- 4108 - 0x100c  :    0 - 0x0
    "00000000", -- 4109 - 0x100d  :    0 - 0x0
    "00000000", -- 4110 - 0x100e  :    0 - 0x0
    "00000000", -- 4111 - 0x100f  :    0 - 0x0
    "00000000", -- 4112 - 0x1010  :    0 - 0x0 -- Background 0x1
    "11000000", -- 4113 - 0x1011  :  192 - 0xc0
    "11110000", -- 4114 - 0x1012  :  240 - 0xf0
    "11111000", -- 4115 - 0x1013  :  248 - 0xf8
    "11111000", -- 4116 - 0x1014  :  248 - 0xf8
    "11111100", -- 4117 - 0x1015  :  252 - 0xfc
    "11111100", -- 4118 - 0x1016  :  252 - 0xfc
    "11111100", -- 4119 - 0x1017  :  252 - 0xfc
    "00000000", -- 4120 - 0x1018  :    0 - 0x0
    "00000000", -- 4121 - 0x1019  :    0 - 0x0
    "00000000", -- 4122 - 0x101a  :    0 - 0x0
    "00000000", -- 4123 - 0x101b  :    0 - 0x0
    "00000000", -- 4124 - 0x101c  :    0 - 0x0
    "00000000", -- 4125 - 0x101d  :    0 - 0x0
    "00000000", -- 4126 - 0x101e  :    0 - 0x0
    "00000000", -- 4127 - 0x101f  :    0 - 0x0
    "00000000", -- 4128 - 0x1020  :    0 - 0x0 -- Background 0x2
    "00000111", -- 4129 - 0x1021  :    7 - 0x7
    "00011111", -- 4130 - 0x1022  :   31 - 0x1f
    "00111111", -- 4131 - 0x1023  :   63 - 0x3f
    "00111111", -- 4132 - 0x1024  :   63 - 0x3f
    "00001111", -- 4133 - 0x1025  :   15 - 0xf
    "00000011", -- 4134 - 0x1026  :    3 - 0x3
    "00000000", -- 4135 - 0x1027  :    0 - 0x0
    "00000000", -- 4136 - 0x1028  :    0 - 0x0
    "00000000", -- 4137 - 0x1029  :    0 - 0x0
    "00000000", -- 4138 - 0x102a  :    0 - 0x0
    "00000000", -- 4139 - 0x102b  :    0 - 0x0
    "00000000", -- 4140 - 0x102c  :    0 - 0x0
    "00000000", -- 4141 - 0x102d  :    0 - 0x0
    "00000000", -- 4142 - 0x102e  :    0 - 0x0
    "00000000", -- 4143 - 0x102f  :    0 - 0x0
    "00000000", -- 4144 - 0x1030  :    0 - 0x0 -- Background 0x3
    "00000000", -- 4145 - 0x1031  :    0 - 0x0
    "00000111", -- 4146 - 0x1032  :    7 - 0x7
    "00011111", -- 4147 - 0x1033  :   31 - 0x1f
    "00111111", -- 4148 - 0x1034  :   63 - 0x3f
    "00111111", -- 4149 - 0x1035  :   63 - 0x3f
    "01111111", -- 4150 - 0x1036  :  127 - 0x7f
    "01111111", -- 4151 - 0x1037  :  127 - 0x7f
    "00000000", -- 4152 - 0x1038  :    0 - 0x0
    "00000000", -- 4153 - 0x1039  :    0 - 0x0
    "00000000", -- 4154 - 0x103a  :    0 - 0x0
    "00000000", -- 4155 - 0x103b  :    0 - 0x0
    "00000000", -- 4156 - 0x103c  :    0 - 0x0
    "00000000", -- 4157 - 0x103d  :    0 - 0x0
    "00000000", -- 4158 - 0x103e  :    0 - 0x0
    "00000000", -- 4159 - 0x103f  :    0 - 0x0
    "01111110", -- 4160 - 0x1040  :  126 - 0x7e -- Background 0x4
    "01111110", -- 4161 - 0x1041  :  126 - 0x7e
    "01111100", -- 4162 - 0x1042  :  124 - 0x7c
    "00111100", -- 4163 - 0x1043  :   60 - 0x3c
    "00111000", -- 4164 - 0x1044  :   56 - 0x38
    "00011000", -- 4165 - 0x1045  :   24 - 0x18
    "00000000", -- 4166 - 0x1046  :    0 - 0x0
    "00000000", -- 4167 - 0x1047  :    0 - 0x0
    "00000000", -- 4168 - 0x1048  :    0 - 0x0
    "00000000", -- 4169 - 0x1049  :    0 - 0x0
    "00000000", -- 4170 - 0x104a  :    0 - 0x0
    "00000000", -- 4171 - 0x104b  :    0 - 0x0
    "00000000", -- 4172 - 0x104c  :    0 - 0x0
    "00000000", -- 4173 - 0x104d  :    0 - 0x0
    "00000000", -- 4174 - 0x104e  :    0 - 0x0
    "00000000", -- 4175 - 0x104f  :    0 - 0x0
    "00000000", -- 4176 - 0x1050  :    0 - 0x0 -- Background 0x5
    "11000000", -- 4177 - 0x1051  :  192 - 0xc0
    "11110000", -- 4178 - 0x1052  :  240 - 0xf0
    "11111000", -- 4179 - 0x1053  :  248 - 0xf8
    "11111000", -- 4180 - 0x1054  :  248 - 0xf8
    "11111100", -- 4181 - 0x1055  :  252 - 0xfc
    "01111100", -- 4182 - 0x1056  :  124 - 0x7c
    "00111100", -- 4183 - 0x1057  :   60 - 0x3c
    "00000000", -- 4184 - 0x1058  :    0 - 0x0
    "00000000", -- 4185 - 0x1059  :    0 - 0x0
    "00000000", -- 4186 - 0x105a  :    0 - 0x0
    "00000000", -- 4187 - 0x105b  :    0 - 0x0
    "00000000", -- 4188 - 0x105c  :    0 - 0x0
    "00000000", -- 4189 - 0x105d  :    0 - 0x0
    "00000000", -- 4190 - 0x105e  :    0 - 0x0
    "00000000", -- 4191 - 0x105f  :    0 - 0x0
    "00000000", -- 4192 - 0x1060  :    0 - 0x0 -- Background 0x6
    "00000111", -- 4193 - 0x1061  :    7 - 0x7
    "00000111", -- 4194 - 0x1062  :    7 - 0x7
    "00000011", -- 4195 - 0x1063  :    3 - 0x3
    "00000001", -- 4196 - 0x1064  :    1 - 0x1
    "00000000", -- 4197 - 0x1065  :    0 - 0x0
    "00000000", -- 4198 - 0x1066  :    0 - 0x0
    "00000000", -- 4199 - 0x1067  :    0 - 0x0
    "00000000", -- 4200 - 0x1068  :    0 - 0x0
    "00000000", -- 4201 - 0x1069  :    0 - 0x0
    "00000000", -- 4202 - 0x106a  :    0 - 0x0
    "00000000", -- 4203 - 0x106b  :    0 - 0x0
    "00000000", -- 4204 - 0x106c  :    0 - 0x0
    "00000000", -- 4205 - 0x106d  :    0 - 0x0
    "00000000", -- 4206 - 0x106e  :    0 - 0x0
    "00000000", -- 4207 - 0x106f  :    0 - 0x0
    "00000000", -- 4208 - 0x1070  :    0 - 0x0 -- Background 0x7
    "00000000", -- 4209 - 0x1071  :    0 - 0x0
    "00000111", -- 4210 - 0x1072  :    7 - 0x7
    "00011111", -- 4211 - 0x1073  :   31 - 0x1f
    "00111111", -- 4212 - 0x1074  :   63 - 0x3f
    "00111111", -- 4213 - 0x1075  :   63 - 0x3f
    "01111110", -- 4214 - 0x1076  :  126 - 0x7e
    "01111100", -- 4215 - 0x1077  :  124 - 0x7c
    "00000000", -- 4216 - 0x1078  :    0 - 0x0
    "00000000", -- 4217 - 0x1079  :    0 - 0x0
    "00000000", -- 4218 - 0x107a  :    0 - 0x0
    "00000000", -- 4219 - 0x107b  :    0 - 0x0
    "00000000", -- 4220 - 0x107c  :    0 - 0x0
    "00000000", -- 4221 - 0x107d  :    0 - 0x0
    "00000000", -- 4222 - 0x107e  :    0 - 0x0
    "00000000", -- 4223 - 0x107f  :    0 - 0x0
    "01111000", -- 4224 - 0x1080  :  120 - 0x78 -- Background 0x8
    "01110000", -- 4225 - 0x1081  :  112 - 0x70
    "01100000", -- 4226 - 0x1082  :   96 - 0x60
    "00000000", -- 4227 - 0x1083  :    0 - 0x0
    "00000000", -- 4228 - 0x1084  :    0 - 0x0
    "00000000", -- 4229 - 0x1085  :    0 - 0x0
    "00000000", -- 4230 - 0x1086  :    0 - 0x0
    "00000000", -- 4231 - 0x1087  :    0 - 0x0
    "00000000", -- 4232 - 0x1088  :    0 - 0x0
    "00000000", -- 4233 - 0x1089  :    0 - 0x0
    "00000000", -- 4234 - 0x108a  :    0 - 0x0
    "00000000", -- 4235 - 0x108b  :    0 - 0x0
    "00000000", -- 4236 - 0x108c  :    0 - 0x0
    "00000000", -- 4237 - 0x108d  :    0 - 0x0
    "00000000", -- 4238 - 0x108e  :    0 - 0x0
    "00000000", -- 4239 - 0x108f  :    0 - 0x0
    "00000000", -- 4240 - 0x1090  :    0 - 0x0 -- Background 0x9
    "00000000", -- 4241 - 0x1091  :    0 - 0x0
    "00000000", -- 4242 - 0x1092  :    0 - 0x0
    "00000000", -- 4243 - 0x1093  :    0 - 0x0
    "00000000", -- 4244 - 0x1094  :    0 - 0x0
    "01000000", -- 4245 - 0x1095  :   64 - 0x40
    "11110000", -- 4246 - 0x1096  :  240 - 0xf0
    "11111000", -- 4247 - 0x1097  :  248 - 0xf8
    "00000000", -- 4248 - 0x1098  :    0 - 0x0
    "00000000", -- 4249 - 0x1099  :    0 - 0x0
    "00000000", -- 4250 - 0x109a  :    0 - 0x0
    "00000000", -- 4251 - 0x109b  :    0 - 0x0
    "00000000", -- 4252 - 0x109c  :    0 - 0x0
    "00000000", -- 4253 - 0x109d  :    0 - 0x0
    "00000000", -- 4254 - 0x109e  :    0 - 0x0
    "00000000", -- 4255 - 0x109f  :    0 - 0x0
    "11111110", -- 4256 - 0x10a0  :  254 - 0xfe -- Background 0xa
    "01111111", -- 4257 - 0x10a1  :  127 - 0x7f
    "01111111", -- 4258 - 0x10a2  :  127 - 0x7f
    "00111111", -- 4259 - 0x10a3  :   63 - 0x3f
    "00001110", -- 4260 - 0x10a4  :   14 - 0xe
    "00000000", -- 4261 - 0x10a5  :    0 - 0x0
    "00000000", -- 4262 - 0x10a6  :    0 - 0x0
    "00000000", -- 4263 - 0x10a7  :    0 - 0x0
    "00000000", -- 4264 - 0x10a8  :    0 - 0x0
    "00000000", -- 4265 - 0x10a9  :    0 - 0x0
    "00000000", -- 4266 - 0x10aa  :    0 - 0x0
    "00000000", -- 4267 - 0x10ab  :    0 - 0x0
    "00000000", -- 4268 - 0x10ac  :    0 - 0x0
    "00000000", -- 4269 - 0x10ad  :    0 - 0x0
    "00000000", -- 4270 - 0x10ae  :    0 - 0x0
    "00000000", -- 4271 - 0x10af  :    0 - 0x0
    "00000000", -- 4272 - 0x10b0  :    0 - 0x0 -- Background 0xb
    "00000000", -- 4273 - 0x10b1  :    0 - 0x0
    "00000000", -- 4274 - 0x10b2  :    0 - 0x0
    "00000000", -- 4275 - 0x10b3  :    0 - 0x0
    "00000000", -- 4276 - 0x10b4  :    0 - 0x0
    "00000000", -- 4277 - 0x10b5  :    0 - 0x0
    "00000000", -- 4278 - 0x10b6  :    0 - 0x0
    "11100000", -- 4279 - 0x10b7  :  224 - 0xe0
    "00000000", -- 4280 - 0x10b8  :    0 - 0x0
    "00000000", -- 4281 - 0x10b9  :    0 - 0x0
    "00000000", -- 4282 - 0x10ba  :    0 - 0x0
    "00000000", -- 4283 - 0x10bb  :    0 - 0x0
    "00000000", -- 4284 - 0x10bc  :    0 - 0x0
    "00000000", -- 4285 - 0x10bd  :    0 - 0x0
    "00000000", -- 4286 - 0x10be  :    0 - 0x0
    "00000000", -- 4287 - 0x10bf  :    0 - 0x0
    "11111100", -- 4288 - 0x10c0  :  252 - 0xfc -- Background 0xc
    "11111111", -- 4289 - 0x10c1  :  255 - 0xff
    "01111111", -- 4290 - 0x10c2  :  127 - 0x7f
    "00111111", -- 4291 - 0x10c3  :   63 - 0x3f
    "00001110", -- 4292 - 0x10c4  :   14 - 0xe
    "00000000", -- 4293 - 0x10c5  :    0 - 0x0
    "00000000", -- 4294 - 0x10c6  :    0 - 0x0
    "00000000", -- 4295 - 0x10c7  :    0 - 0x0
    "00000000", -- 4296 - 0x10c8  :    0 - 0x0
    "00000000", -- 4297 - 0x10c9  :    0 - 0x0
    "00000000", -- 4298 - 0x10ca  :    0 - 0x0
    "00000000", -- 4299 - 0x10cb  :    0 - 0x0
    "00000000", -- 4300 - 0x10cc  :    0 - 0x0
    "00000000", -- 4301 - 0x10cd  :    0 - 0x0
    "00000000", -- 4302 - 0x10ce  :    0 - 0x0
    "00000000", -- 4303 - 0x10cf  :    0 - 0x0
    "11110000", -- 4304 - 0x10d0  :  240 - 0xf0 -- Background 0xd
    "11111111", -- 4305 - 0x10d1  :  255 - 0xff
    "11111111", -- 4306 - 0x10d2  :  255 - 0xff
    "01111111", -- 4307 - 0x10d3  :  127 - 0x7f
    "00011110", -- 4308 - 0x10d4  :   30 - 0x1e
    "00000000", -- 4309 - 0x10d5  :    0 - 0x0
    "00000000", -- 4310 - 0x10d6  :    0 - 0x0
    "00000000", -- 4311 - 0x10d7  :    0 - 0x0
    "00000000", -- 4312 - 0x10d8  :    0 - 0x0
    "00000000", -- 4313 - 0x10d9  :    0 - 0x0
    "00000000", -- 4314 - 0x10da  :    0 - 0x0
    "00000000", -- 4315 - 0x10db  :    0 - 0x0
    "00000000", -- 4316 - 0x10dc  :    0 - 0x0
    "00000000", -- 4317 - 0x10dd  :    0 - 0x0
    "00000000", -- 4318 - 0x10de  :    0 - 0x0
    "00000000", -- 4319 - 0x10df  :    0 - 0x0
    "00000000", -- 4320 - 0x10e0  :    0 - 0x0 -- Background 0xe
    "00001111", -- 4321 - 0x10e1  :   15 - 0xf
    "11111111", -- 4322 - 0x10e2  :  255 - 0xff
    "11111111", -- 4323 - 0x10e3  :  255 - 0xff
    "01111111", -- 4324 - 0x10e4  :  127 - 0x7f
    "00011110", -- 4325 - 0x10e5  :   30 - 0x1e
    "00000000", -- 4326 - 0x10e6  :    0 - 0x0
    "00000000", -- 4327 - 0x10e7  :    0 - 0x0
    "00000000", -- 4328 - 0x10e8  :    0 - 0x0
    "00000000", -- 4329 - 0x10e9  :    0 - 0x0
    "00000000", -- 4330 - 0x10ea  :    0 - 0x0
    "00000000", -- 4331 - 0x10eb  :    0 - 0x0
    "00000000", -- 4332 - 0x10ec  :    0 - 0x0
    "00000000", -- 4333 - 0x10ed  :    0 - 0x0
    "00000000", -- 4334 - 0x10ee  :    0 - 0x0
    "00000000", -- 4335 - 0x10ef  :    0 - 0x0
    "00000000", -- 4336 - 0x10f0  :    0 - 0x0 -- Background 0xf
    "00000011", -- 4337 - 0x10f1  :    3 - 0x3
    "00001111", -- 4338 - 0x10f2  :   15 - 0xf
    "01111111", -- 4339 - 0x10f3  :  127 - 0x7f
    "11111111", -- 4340 - 0x10f4  :  255 - 0xff
    "01111110", -- 4341 - 0x10f5  :  126 - 0x7e
    "00011100", -- 4342 - 0x10f6  :   28 - 0x1c
    "00000000", -- 4343 - 0x10f7  :    0 - 0x0
    "00000000", -- 4344 - 0x10f8  :    0 - 0x0
    "00000000", -- 4345 - 0x10f9  :    0 - 0x0
    "00000000", -- 4346 - 0x10fa  :    0 - 0x0
    "00000000", -- 4347 - 0x10fb  :    0 - 0x0
    "00000000", -- 4348 - 0x10fc  :    0 - 0x0
    "00000000", -- 4349 - 0x10fd  :    0 - 0x0
    "00000000", -- 4350 - 0x10fe  :    0 - 0x0
    "00000000", -- 4351 - 0x10ff  :    0 - 0x0
    "00000000", -- 4352 - 0x1100  :    0 - 0x0 -- Background 0x10
    "00000001", -- 4353 - 0x1101  :    1 - 0x1
    "00000011", -- 4354 - 0x1102  :    3 - 0x3
    "00001111", -- 4355 - 0x1103  :   15 - 0xf
    "00011111", -- 4356 - 0x1104  :   31 - 0x1f
    "01111111", -- 4357 - 0x1105  :  127 - 0x7f
    "01111110", -- 4358 - 0x1106  :  126 - 0x7e
    "00111100", -- 4359 - 0x1107  :   60 - 0x3c
    "00000000", -- 4360 - 0x1108  :    0 - 0x0
    "00000000", -- 4361 - 0x1109  :    0 - 0x0
    "00000000", -- 4362 - 0x110a  :    0 - 0x0
    "00000000", -- 4363 - 0x110b  :    0 - 0x0
    "00000000", -- 4364 - 0x110c  :    0 - 0x0
    "00000000", -- 4365 - 0x110d  :    0 - 0x0
    "00000000", -- 4366 - 0x110e  :    0 - 0x0
    "00000000", -- 4367 - 0x110f  :    0 - 0x0
    "00000000", -- 4368 - 0x1110  :    0 - 0x0 -- Background 0x11
    "00000001", -- 4369 - 0x1111  :    1 - 0x1
    "00000011", -- 4370 - 0x1112  :    3 - 0x3
    "00000111", -- 4371 - 0x1113  :    7 - 0x7
    "00000111", -- 4372 - 0x1114  :    7 - 0x7
    "00001111", -- 4373 - 0x1115  :   15 - 0xf
    "00011111", -- 4374 - 0x1116  :   31 - 0x1f
    "00001110", -- 4375 - 0x1117  :   14 - 0xe
    "00000000", -- 4376 - 0x1118  :    0 - 0x0
    "00000000", -- 4377 - 0x1119  :    0 - 0x0
    "00000000", -- 4378 - 0x111a  :    0 - 0x0
    "00000000", -- 4379 - 0x111b  :    0 - 0x0
    "00000000", -- 4380 - 0x111c  :    0 - 0x0
    "00000000", -- 4381 - 0x111d  :    0 - 0x0
    "00000000", -- 4382 - 0x111e  :    0 - 0x0
    "00000000", -- 4383 - 0x111f  :    0 - 0x0
    "00000000", -- 4384 - 0x1120  :    0 - 0x0 -- Background 0x12
    "00000000", -- 4385 - 0x1121  :    0 - 0x0
    "00000001", -- 4386 - 0x1122  :    1 - 0x1
    "00000011", -- 4387 - 0x1123  :    3 - 0x3
    "00000011", -- 4388 - 0x1124  :    3 - 0x3
    "00000011", -- 4389 - 0x1125  :    3 - 0x3
    "00000111", -- 4390 - 0x1126  :    7 - 0x7
    "00000010", -- 4391 - 0x1127  :    2 - 0x2
    "00000000", -- 4392 - 0x1128  :    0 - 0x0
    "00000000", -- 4393 - 0x1129  :    0 - 0x0
    "00000000", -- 4394 - 0x112a  :    0 - 0x0
    "00000000", -- 4395 - 0x112b  :    0 - 0x0
    "00000000", -- 4396 - 0x112c  :    0 - 0x0
    "00000000", -- 4397 - 0x112d  :    0 - 0x0
    "00000000", -- 4398 - 0x112e  :    0 - 0x0
    "00000000", -- 4399 - 0x112f  :    0 - 0x0
    "00000000", -- 4400 - 0x1130  :    0 - 0x0 -- Background 0x13
    "00000000", -- 4401 - 0x1131  :    0 - 0x0
    "00000001", -- 4402 - 0x1132  :    1 - 0x1
    "00000001", -- 4403 - 0x1133  :    1 - 0x1
    "00000001", -- 4404 - 0x1134  :    1 - 0x1
    "00000001", -- 4405 - 0x1135  :    1 - 0x1
    "00000001", -- 4406 - 0x1136  :    1 - 0x1
    "00000001", -- 4407 - 0x1137  :    1 - 0x1
    "00000000", -- 4408 - 0x1138  :    0 - 0x0
    "00000000", -- 4409 - 0x1139  :    0 - 0x0
    "00000000", -- 4410 - 0x113a  :    0 - 0x0
    "00000000", -- 4411 - 0x113b  :    0 - 0x0
    "00000000", -- 4412 - 0x113c  :    0 - 0x0
    "00000000", -- 4413 - 0x113d  :    0 - 0x0
    "00000000", -- 4414 - 0x113e  :    0 - 0x0
    "00000000", -- 4415 - 0x113f  :    0 - 0x0
    "00000000", -- 4416 - 0x1140  :    0 - 0x0 -- Background 0x14
    "00000000", -- 4417 - 0x1141  :    0 - 0x0
    "00000000", -- 4418 - 0x1142  :    0 - 0x0
    "00000000", -- 4419 - 0x1143  :    0 - 0x0
    "00000000", -- 4420 - 0x1144  :    0 - 0x0
    "00000000", -- 4421 - 0x1145  :    0 - 0x0
    "00000100", -- 4422 - 0x1146  :    4 - 0x4
    "00000010", -- 4423 - 0x1147  :    2 - 0x2
    "00000000", -- 4424 - 0x1148  :    0 - 0x0
    "00000000", -- 4425 - 0x1149  :    0 - 0x0
    "00000000", -- 4426 - 0x114a  :    0 - 0x0
    "00000000", -- 4427 - 0x114b  :    0 - 0x0
    "00000000", -- 4428 - 0x114c  :    0 - 0x0
    "00000000", -- 4429 - 0x114d  :    0 - 0x0
    "00000000", -- 4430 - 0x114e  :    0 - 0x0
    "00000000", -- 4431 - 0x114f  :    0 - 0x0
    "00000000", -- 4432 - 0x1150  :    0 - 0x0 -- Background 0x15
    "00000000", -- 4433 - 0x1151  :    0 - 0x0
    "00000000", -- 4434 - 0x1152  :    0 - 0x0
    "00000000", -- 4435 - 0x1153  :    0 - 0x0
    "00000000", -- 4436 - 0x1154  :    0 - 0x0
    "00000000", -- 4437 - 0x1155  :    0 - 0x0
    "00100000", -- 4438 - 0x1156  :   32 - 0x20
    "01001000", -- 4439 - 0x1157  :   72 - 0x48
    "00000000", -- 4440 - 0x1158  :    0 - 0x0
    "00000000", -- 4441 - 0x1159  :    0 - 0x0
    "00000000", -- 4442 - 0x115a  :    0 - 0x0
    "00000000", -- 4443 - 0x115b  :    0 - 0x0
    "00000000", -- 4444 - 0x115c  :    0 - 0x0
    "00000000", -- 4445 - 0x115d  :    0 - 0x0
    "00000000", -- 4446 - 0x115e  :    0 - 0x0
    "00000000", -- 4447 - 0x115f  :    0 - 0x0
    "00010000", -- 4448 - 0x1160  :   16 - 0x10 -- Background 0x16
    "00001000", -- 4449 - 0x1161  :    8 - 0x8
    "00000000", -- 4450 - 0x1162  :    0 - 0x0
    "00110000", -- 4451 - 0x1163  :   48 - 0x30
    "00000000", -- 4452 - 0x1164  :    0 - 0x0
    "00001000", -- 4453 - 0x1165  :    8 - 0x8
    "00010010", -- 4454 - 0x1166  :   18 - 0x12
    "00000100", -- 4455 - 0x1167  :    4 - 0x4
    "00000000", -- 4456 - 0x1168  :    0 - 0x0
    "00000000", -- 4457 - 0x1169  :    0 - 0x0
    "00000000", -- 4458 - 0x116a  :    0 - 0x0
    "00000000", -- 4459 - 0x116b  :    0 - 0x0
    "00000000", -- 4460 - 0x116c  :    0 - 0x0
    "00000000", -- 4461 - 0x116d  :    0 - 0x0
    "00000000", -- 4462 - 0x116e  :    0 - 0x0
    "00000000", -- 4463 - 0x116f  :    0 - 0x0
    "00010000", -- 4464 - 0x1170  :   16 - 0x10 -- Background 0x17
    "00000000", -- 4465 - 0x1171  :    0 - 0x0
    "00001100", -- 4466 - 0x1172  :   12 - 0xc
    "00000000", -- 4467 - 0x1173  :    0 - 0x0
    "00010000", -- 4468 - 0x1174  :   16 - 0x10
    "00001000", -- 4469 - 0x1175  :    8 - 0x8
    "01000000", -- 4470 - 0x1176  :   64 - 0x40
    "00100000", -- 4471 - 0x1177  :   32 - 0x20
    "00000000", -- 4472 - 0x1178  :    0 - 0x0
    "00000000", -- 4473 - 0x1179  :    0 - 0x0
    "00000000", -- 4474 - 0x117a  :    0 - 0x0
    "00000000", -- 4475 - 0x117b  :    0 - 0x0
    "00000000", -- 4476 - 0x117c  :    0 - 0x0
    "00000000", -- 4477 - 0x117d  :    0 - 0x0
    "00000000", -- 4478 - 0x117e  :    0 - 0x0
    "00000000", -- 4479 - 0x117f  :    0 - 0x0
    "00000000", -- 4480 - 0x1180  :    0 - 0x0 -- Background 0x18
    "00000000", -- 4481 - 0x1181  :    0 - 0x0
    "00000011", -- 4482 - 0x1182  :    3 - 0x3
    "00000011", -- 4483 - 0x1183  :    3 - 0x3
    "00000001", -- 4484 - 0x1184  :    1 - 0x1
    "00100001", -- 4485 - 0x1185  :   33 - 0x21
    "00100001", -- 4486 - 0x1186  :   33 - 0x21
    "01110011", -- 4487 - 0x1187  :  115 - 0x73
    "00000000", -- 4488 - 0x1188  :    0 - 0x0
    "00000000", -- 4489 - 0x1189  :    0 - 0x0
    "00000011", -- 4490 - 0x118a  :    3 - 0x3
    "00000011", -- 4491 - 0x118b  :    3 - 0x3
    "00010011", -- 4492 - 0x118c  :   19 - 0x13
    "00111111", -- 4493 - 0x118d  :   63 - 0x3f
    "00111111", -- 4494 - 0x118e  :   63 - 0x3f
    "01111111", -- 4495 - 0x118f  :  127 - 0x7f
    "01111111", -- 4496 - 0x1190  :  127 - 0x7f -- Background 0x19
    "01111111", -- 4497 - 0x1191  :  127 - 0x7f
    "01111111", -- 4498 - 0x1192  :  127 - 0x7f
    "01111111", -- 4499 - 0x1193  :  127 - 0x7f
    "01101110", -- 4500 - 0x1194  :  110 - 0x6e
    "01000110", -- 4501 - 0x1195  :   70 - 0x46
    "00000000", -- 4502 - 0x1196  :    0 - 0x0
    "00000000", -- 4503 - 0x1197  :    0 - 0x0
    "01111111", -- 4504 - 0x1198  :  127 - 0x7f
    "01111111", -- 4505 - 0x1199  :  127 - 0x7f
    "01111111", -- 4506 - 0x119a  :  127 - 0x7f
    "01111111", -- 4507 - 0x119b  :  127 - 0x7f
    "01101110", -- 4508 - 0x119c  :  110 - 0x6e
    "01000110", -- 4509 - 0x119d  :   70 - 0x46
    "00000000", -- 4510 - 0x119e  :    0 - 0x0
    "00000000", -- 4511 - 0x119f  :    0 - 0x0
    "01111111", -- 4512 - 0x11a0  :  127 - 0x7f -- Background 0x1a
    "01111111", -- 4513 - 0x11a1  :  127 - 0x7f
    "01111111", -- 4514 - 0x11a2  :  127 - 0x7f
    "01111111", -- 4515 - 0x11a3  :  127 - 0x7f
    "01111011", -- 4516 - 0x11a4  :  123 - 0x7b
    "00110001", -- 4517 - 0x11a5  :   49 - 0x31
    "00000000", -- 4518 - 0x11a6  :    0 - 0x0
    "00000000", -- 4519 - 0x11a7  :    0 - 0x0
    "01111111", -- 4520 - 0x11a8  :  127 - 0x7f
    "01111111", -- 4521 - 0x11a9  :  127 - 0x7f
    "01111111", -- 4522 - 0x11aa  :  127 - 0x7f
    "01111111", -- 4523 - 0x11ab  :  127 - 0x7f
    "01111011", -- 4524 - 0x11ac  :  123 - 0x7b
    "00110001", -- 4525 - 0x11ad  :   49 - 0x31
    "00000000", -- 4526 - 0x11ae  :    0 - 0x0
    "00000000", -- 4527 - 0x11af  :    0 - 0x0
    "00000000", -- 4528 - 0x11b0  :    0 - 0x0 -- Background 0x1b
    "00000011", -- 4529 - 0x11b1  :    3 - 0x3
    "00001111", -- 4530 - 0x11b2  :   15 - 0xf
    "00011111", -- 4531 - 0x11b3  :   31 - 0x1f
    "00100111", -- 4532 - 0x11b4  :   39 - 0x27
    "00000011", -- 4533 - 0x11b5  :    3 - 0x3
    "00000011", -- 4534 - 0x11b6  :    3 - 0x3
    "01000011", -- 4535 - 0x11b7  :   67 - 0x43
    "00000000", -- 4536 - 0x11b8  :    0 - 0x0
    "00000011", -- 4537 - 0x11b9  :    3 - 0x3
    "00001111", -- 4538 - 0x11ba  :   15 - 0xf
    "00011111", -- 4539 - 0x11bb  :   31 - 0x1f
    "00111111", -- 4540 - 0x11bc  :   63 - 0x3f
    "00111111", -- 4541 - 0x11bd  :   63 - 0x3f
    "00001111", -- 4542 - 0x11be  :   15 - 0xf
    "01001111", -- 4543 - 0x11bf  :   79 - 0x4f
    "00000000", -- 4544 - 0x11c0  :    0 - 0x0 -- Background 0x1c
    "11000000", -- 4545 - 0x11c1  :  192 - 0xc0
    "11110000", -- 4546 - 0x11c2  :  240 - 0xf0
    "11111000", -- 4547 - 0x11c3  :  248 - 0xf8
    "10011100", -- 4548 - 0x11c4  :  156 - 0x9c
    "00001100", -- 4549 - 0x11c5  :   12 - 0xc
    "00001100", -- 4550 - 0x11c6  :   12 - 0xc
    "00001110", -- 4551 - 0x11c7  :   14 - 0xe
    "00000000", -- 4552 - 0x11c8  :    0 - 0x0
    "11000000", -- 4553 - 0x11c9  :  192 - 0xc0
    "11110000", -- 4554 - 0x11ca  :  240 - 0xf0
    "11111000", -- 4555 - 0x11cb  :  248 - 0xf8
    "11111100", -- 4556 - 0x11cc  :  252 - 0xfc
    "11111100", -- 4557 - 0x11cd  :  252 - 0xfc
    "00111100", -- 4558 - 0x11ce  :   60 - 0x3c
    "00111110", -- 4559 - 0x11cf  :   62 - 0x3e
    "01100111", -- 4560 - 0x11d0  :  103 - 0x67 -- Background 0x1d
    "01111111", -- 4561 - 0x11d1  :  127 - 0x7f
    "01111111", -- 4562 - 0x11d2  :  127 - 0x7f
    "01111111", -- 4563 - 0x11d3  :  127 - 0x7f
    "01101110", -- 4564 - 0x11d4  :  110 - 0x6e
    "01000110", -- 4565 - 0x11d5  :   70 - 0x46
    "00000000", -- 4566 - 0x11d6  :    0 - 0x0
    "00000000", -- 4567 - 0x11d7  :    0 - 0x0
    "01111111", -- 4568 - 0x11d8  :  127 - 0x7f
    "01111111", -- 4569 - 0x11d9  :  127 - 0x7f
    "01111111", -- 4570 - 0x11da  :  127 - 0x7f
    "01111111", -- 4571 - 0x11db  :  127 - 0x7f
    "01101110", -- 4572 - 0x11dc  :  110 - 0x6e
    "01000110", -- 4573 - 0x11dd  :   70 - 0x46
    "00000000", -- 4574 - 0x11de  :    0 - 0x0
    "00000000", -- 4575 - 0x11df  :    0 - 0x0
    "01100111", -- 4576 - 0x11e0  :  103 - 0x67 -- Background 0x1e
    "01111111", -- 4577 - 0x11e1  :  127 - 0x7f
    "01111111", -- 4578 - 0x11e2  :  127 - 0x7f
    "01111111", -- 4579 - 0x11e3  :  127 - 0x7f
    "01111011", -- 4580 - 0x11e4  :  123 - 0x7b
    "00110001", -- 4581 - 0x11e5  :   49 - 0x31
    "00000000", -- 4582 - 0x11e6  :    0 - 0x0
    "00000000", -- 4583 - 0x11e7  :    0 - 0x0
    "01111111", -- 4584 - 0x11e8  :  127 - 0x7f
    "01111111", -- 4585 - 0x11e9  :  127 - 0x7f
    "01111111", -- 4586 - 0x11ea  :  127 - 0x7f
    "01111111", -- 4587 - 0x11eb  :  127 - 0x7f
    "01111011", -- 4588 - 0x11ec  :  123 - 0x7b
    "00110001", -- 4589 - 0x11ed  :   49 - 0x31
    "00000000", -- 4590 - 0x11ee  :    0 - 0x0
    "00000000", -- 4591 - 0x11ef  :    0 - 0x0
    "10011110", -- 4592 - 0x11f0  :  158 - 0x9e -- Background 0x1f
    "11111110", -- 4593 - 0x11f1  :  254 - 0xfe
    "11111110", -- 4594 - 0x11f2  :  254 - 0xfe
    "11111110", -- 4595 - 0x11f3  :  254 - 0xfe
    "01110110", -- 4596 - 0x11f4  :  118 - 0x76
    "01100010", -- 4597 - 0x11f5  :   98 - 0x62
    "00000000", -- 4598 - 0x11f6  :    0 - 0x0
    "00000000", -- 4599 - 0x11f7  :    0 - 0x0
    "11111110", -- 4600 - 0x11f8  :  254 - 0xfe
    "11111110", -- 4601 - 0x11f9  :  254 - 0xfe
    "11111110", -- 4602 - 0x11fa  :  254 - 0xfe
    "11111110", -- 4603 - 0x11fb  :  254 - 0xfe
    "01110110", -- 4604 - 0x11fc  :  118 - 0x76
    "01100010", -- 4605 - 0x11fd  :   98 - 0x62
    "00000000", -- 4606 - 0x11fe  :    0 - 0x0
    "00000000", -- 4607 - 0x11ff  :    0 - 0x0
    "10011110", -- 4608 - 0x1200  :  158 - 0x9e -- Background 0x20
    "11111110", -- 4609 - 0x1201  :  254 - 0xfe
    "11111110", -- 4610 - 0x1202  :  254 - 0xfe
    "11111110", -- 4611 - 0x1203  :  254 - 0xfe
    "11011110", -- 4612 - 0x1204  :  222 - 0xde
    "10001100", -- 4613 - 0x1205  :  140 - 0x8c
    "00000000", -- 4614 - 0x1206  :    0 - 0x0
    "00000000", -- 4615 - 0x1207  :    0 - 0x0
    "11111110", -- 4616 - 0x1208  :  254 - 0xfe
    "11111110", -- 4617 - 0x1209  :  254 - 0xfe
    "11111110", -- 4618 - 0x120a  :  254 - 0xfe
    "11111110", -- 4619 - 0x120b  :  254 - 0xfe
    "11011110", -- 4620 - 0x120c  :  222 - 0xde
    "10001100", -- 4621 - 0x120d  :  140 - 0x8c
    "00000000", -- 4622 - 0x120e  :    0 - 0x0
    "00000000", -- 4623 - 0x120f  :    0 - 0x0
    "00000000", -- 4624 - 0x1210  :    0 - 0x0 -- Background 0x21
    "00000011", -- 4625 - 0x1211  :    3 - 0x3
    "00001111", -- 4626 - 0x1212  :   15 - 0xf
    "00011111", -- 4627 - 0x1213  :   31 - 0x1f
    "00111111", -- 4628 - 0x1214  :   63 - 0x3f
    "00110011", -- 4629 - 0x1215  :   51 - 0x33
    "00100001", -- 4630 - 0x1216  :   33 - 0x21
    "01100001", -- 4631 - 0x1217  :   97 - 0x61
    "00000000", -- 4632 - 0x1218  :    0 - 0x0
    "00000011", -- 4633 - 0x1219  :    3 - 0x3
    "00001111", -- 4634 - 0x121a  :   15 - 0xf
    "00011111", -- 4635 - 0x121b  :   31 - 0x1f
    "00111111", -- 4636 - 0x121c  :   63 - 0x3f
    "00111111", -- 4637 - 0x121d  :   63 - 0x3f
    "00111111", -- 4638 - 0x121e  :   63 - 0x3f
    "01111111", -- 4639 - 0x121f  :  127 - 0x7f
    "01100001", -- 4640 - 0x1220  :   97 - 0x61 -- Background 0x22
    "01110011", -- 4641 - 0x1221  :  115 - 0x73
    "01111111", -- 4642 - 0x1222  :  127 - 0x7f
    "01111111", -- 4643 - 0x1223  :  127 - 0x7f
    "01101110", -- 4644 - 0x1224  :  110 - 0x6e
    "01000110", -- 4645 - 0x1225  :   70 - 0x46
    "00000000", -- 4646 - 0x1226  :    0 - 0x0
    "00000000", -- 4647 - 0x1227  :    0 - 0x0
    "01110011", -- 4648 - 0x1228  :  115 - 0x73
    "01110011", -- 4649 - 0x1229  :  115 - 0x73
    "01111111", -- 4650 - 0x122a  :  127 - 0x7f
    "01111111", -- 4651 - 0x122b  :  127 - 0x7f
    "01101110", -- 4652 - 0x122c  :  110 - 0x6e
    "01000110", -- 4653 - 0x122d  :   70 - 0x46
    "00000000", -- 4654 - 0x122e  :    0 - 0x0
    "00000000", -- 4655 - 0x122f  :    0 - 0x0
    "01100001", -- 4656 - 0x1230  :   97 - 0x61 -- Background 0x23
    "01110011", -- 4657 - 0x1231  :  115 - 0x73
    "01111111", -- 4658 - 0x1232  :  127 - 0x7f
    "01111111", -- 4659 - 0x1233  :  127 - 0x7f
    "01110111", -- 4660 - 0x1234  :  119 - 0x77
    "00100011", -- 4661 - 0x1235  :   35 - 0x23
    "00000000", -- 4662 - 0x1236  :    0 - 0x0
    "00000000", -- 4663 - 0x1237  :    0 - 0x0
    "01110011", -- 4664 - 0x1238  :  115 - 0x73
    "01110011", -- 4665 - 0x1239  :  115 - 0x73
    "01111111", -- 4666 - 0x123a  :  127 - 0x7f
    "01111111", -- 4667 - 0x123b  :  127 - 0x7f
    "01110111", -- 4668 - 0x123c  :  119 - 0x77
    "00100011", -- 4669 - 0x123d  :   35 - 0x23
    "00000000", -- 4670 - 0x123e  :    0 - 0x0
    "00000000", -- 4671 - 0x123f  :    0 - 0x0
    "00000000", -- 4672 - 0x1240  :    0 - 0x0 -- Background 0x24
    "00000011", -- 4673 - 0x1241  :    3 - 0x3
    "00001111", -- 4674 - 0x1242  :   15 - 0xf
    "00011111", -- 4675 - 0x1243  :   31 - 0x1f
    "00111111", -- 4676 - 0x1244  :   63 - 0x3f
    "00111111", -- 4677 - 0x1245  :   63 - 0x3f
    "00111111", -- 4678 - 0x1246  :   63 - 0x3f
    "01111111", -- 4679 - 0x1247  :  127 - 0x7f
    "00000000", -- 4680 - 0x1248  :    0 - 0x0
    "00000000", -- 4681 - 0x1249  :    0 - 0x0
    "00000000", -- 4682 - 0x124a  :    0 - 0x0
    "00000000", -- 4683 - 0x124b  :    0 - 0x0
    "00000000", -- 4684 - 0x124c  :    0 - 0x0
    "00000110", -- 4685 - 0x124d  :    6 - 0x6
    "00000110", -- 4686 - 0x124e  :    6 - 0x6
    "00000000", -- 4687 - 0x124f  :    0 - 0x0
    "01111111", -- 4688 - 0x1250  :  127 - 0x7f -- Background 0x25
    "01111111", -- 4689 - 0x1251  :  127 - 0x7f
    "01111111", -- 4690 - 0x1252  :  127 - 0x7f
    "01111111", -- 4691 - 0x1253  :  127 - 0x7f
    "01101110", -- 4692 - 0x1254  :  110 - 0x6e
    "01000110", -- 4693 - 0x1255  :   70 - 0x46
    "00000000", -- 4694 - 0x1256  :    0 - 0x0
    "00000000", -- 4695 - 0x1257  :    0 - 0x0
    "00000000", -- 4696 - 0x1258  :    0 - 0x0
    "00011001", -- 4697 - 0x1259  :   25 - 0x19
    "00100110", -- 4698 - 0x125a  :   38 - 0x26
    "00000000", -- 4699 - 0x125b  :    0 - 0x0
    "00000000", -- 4700 - 0x125c  :    0 - 0x0
    "00000000", -- 4701 - 0x125d  :    0 - 0x0
    "00000000", -- 4702 - 0x125e  :    0 - 0x0
    "00000000", -- 4703 - 0x125f  :    0 - 0x0
    "01111111", -- 4704 - 0x1260  :  127 - 0x7f -- Background 0x26
    "01111111", -- 4705 - 0x1261  :  127 - 0x7f
    "01111111", -- 4706 - 0x1262  :  127 - 0x7f
    "01111111", -- 4707 - 0x1263  :  127 - 0x7f
    "01111011", -- 4708 - 0x1264  :  123 - 0x7b
    "00110001", -- 4709 - 0x1265  :   49 - 0x31
    "00000000", -- 4710 - 0x1266  :    0 - 0x0
    "00000000", -- 4711 - 0x1267  :    0 - 0x0
    "00000000", -- 4712 - 0x1268  :    0 - 0x0
    "00011001", -- 4713 - 0x1269  :   25 - 0x19
    "00100110", -- 4714 - 0x126a  :   38 - 0x26
    "00000000", -- 4715 - 0x126b  :    0 - 0x0
    "00000000", -- 4716 - 0x126c  :    0 - 0x0
    "00000000", -- 4717 - 0x126d  :    0 - 0x0
    "00000000", -- 4718 - 0x126e  :    0 - 0x0
    "00000000", -- 4719 - 0x126f  :    0 - 0x0
    "00000000", -- 4720 - 0x1270  :    0 - 0x0 -- Background 0x27
    "00000000", -- 4721 - 0x1271  :    0 - 0x0
    "00000000", -- 4722 - 0x1272  :    0 - 0x0
    "00000000", -- 4723 - 0x1273  :    0 - 0x0
    "00000000", -- 4724 - 0x1274  :    0 - 0x0
    "00000000", -- 4725 - 0x1275  :    0 - 0x0
    "00000000", -- 4726 - 0x1276  :    0 - 0x0
    "00000000", -- 4727 - 0x1277  :    0 - 0x0
    "00000000", -- 4728 - 0x1278  :    0 - 0x0
    "00001100", -- 4729 - 0x1279  :   12 - 0xc
    "00010010", -- 4730 - 0x127a  :   18 - 0x12
    "00010010", -- 4731 - 0x127b  :   18 - 0x12
    "00011110", -- 4732 - 0x127c  :   30 - 0x1e
    "00001100", -- 4733 - 0x127d  :   12 - 0xc
    "00000000", -- 4734 - 0x127e  :    0 - 0x0
    "00000000", -- 4735 - 0x127f  :    0 - 0x0
    "00000000", -- 4736 - 0x1280  :    0 - 0x0 -- Background 0x28
    "00000000", -- 4737 - 0x1281  :    0 - 0x0
    "00000000", -- 4738 - 0x1282  :    0 - 0x0
    "00000000", -- 4739 - 0x1283  :    0 - 0x0
    "00000000", -- 4740 - 0x1284  :    0 - 0x0
    "00000000", -- 4741 - 0x1285  :    0 - 0x0
    "00000000", -- 4742 - 0x1286  :    0 - 0x0
    "00000000", -- 4743 - 0x1287  :    0 - 0x0
    "00000000", -- 4744 - 0x1288  :    0 - 0x0
    "00000000", -- 4745 - 0x1289  :    0 - 0x0
    "00000000", -- 4746 - 0x128a  :    0 - 0x0
    "00000000", -- 4747 - 0x128b  :    0 - 0x0
    "00000000", -- 4748 - 0x128c  :    0 - 0x0
    "00111000", -- 4749 - 0x128d  :   56 - 0x38
    "01001101", -- 4750 - 0x128e  :   77 - 0x4d
    "01001101", -- 4751 - 0x128f  :   77 - 0x4d
    "00000000", -- 4752 - 0x1290  :    0 - 0x0 -- Background 0x29
    "00000000", -- 4753 - 0x1291  :    0 - 0x0
    "00000000", -- 4754 - 0x1292  :    0 - 0x0
    "00000000", -- 4755 - 0x1293  :    0 - 0x0
    "00000000", -- 4756 - 0x1294  :    0 - 0x0
    "00000000", -- 4757 - 0x1295  :    0 - 0x0
    "00000000", -- 4758 - 0x1296  :    0 - 0x0
    "00000000", -- 4759 - 0x1297  :    0 - 0x0
    "00000000", -- 4760 - 0x1298  :    0 - 0x0
    "00000000", -- 4761 - 0x1299  :    0 - 0x0
    "00000000", -- 4762 - 0x129a  :    0 - 0x0
    "00000000", -- 4763 - 0x129b  :    0 - 0x0
    "00000000", -- 4764 - 0x129c  :    0 - 0x0
    "11100000", -- 4765 - 0x129d  :  224 - 0xe0
    "00110000", -- 4766 - 0x129e  :   48 - 0x30
    "00110000", -- 4767 - 0x129f  :   48 - 0x30
    "00000000", -- 4768 - 0x12a0  :    0 - 0x0 -- Background 0x2a
    "00000000", -- 4769 - 0x12a1  :    0 - 0x0
    "00000000", -- 4770 - 0x12a2  :    0 - 0x0
    "00000000", -- 4771 - 0x12a3  :    0 - 0x0
    "00000000", -- 4772 - 0x12a4  :    0 - 0x0
    "00000000", -- 4773 - 0x12a5  :    0 - 0x0
    "00000000", -- 4774 - 0x12a6  :    0 - 0x0
    "00000000", -- 4775 - 0x12a7  :    0 - 0x0
    "00111000", -- 4776 - 0x12a8  :   56 - 0x38
    "00000000", -- 4777 - 0x12a9  :    0 - 0x0
    "00000000", -- 4778 - 0x12aa  :    0 - 0x0
    "00000000", -- 4779 - 0x12ab  :    0 - 0x0
    "00000000", -- 4780 - 0x12ac  :    0 - 0x0
    "00000000", -- 4781 - 0x12ad  :    0 - 0x0
    "00000000", -- 4782 - 0x12ae  :    0 - 0x0
    "00000000", -- 4783 - 0x12af  :    0 - 0x0
    "00000000", -- 4784 - 0x12b0  :    0 - 0x0 -- Background 0x2b
    "00000000", -- 4785 - 0x12b1  :    0 - 0x0
    "00000000", -- 4786 - 0x12b2  :    0 - 0x0
    "00000000", -- 4787 - 0x12b3  :    0 - 0x0
    "00000000", -- 4788 - 0x12b4  :    0 - 0x0
    "00000000", -- 4789 - 0x12b5  :    0 - 0x0
    "00000000", -- 4790 - 0x12b6  :    0 - 0x0
    "00000000", -- 4791 - 0x12b7  :    0 - 0x0
    "11100000", -- 4792 - 0x12b8  :  224 - 0xe0
    "00000000", -- 4793 - 0x12b9  :    0 - 0x0
    "00000000", -- 4794 - 0x12ba  :    0 - 0x0
    "00000000", -- 4795 - 0x12bb  :    0 - 0x0
    "00000000", -- 4796 - 0x12bc  :    0 - 0x0
    "00000000", -- 4797 - 0x12bd  :    0 - 0x0
    "00000000", -- 4798 - 0x12be  :    0 - 0x0
    "00000000", -- 4799 - 0x12bf  :    0 - 0x0
    "00000000", -- 4800 - 0x12c0  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 4801 - 0x12c1  :    0 - 0x0
    "00000000", -- 4802 - 0x12c2  :    0 - 0x0
    "00000000", -- 4803 - 0x12c3  :    0 - 0x0
    "00000000", -- 4804 - 0x12c4  :    0 - 0x0
    "00000000", -- 4805 - 0x12c5  :    0 - 0x0
    "00000000", -- 4806 - 0x12c6  :    0 - 0x0
    "00000000", -- 4807 - 0x12c7  :    0 - 0x0
    "00000000", -- 4808 - 0x12c8  :    0 - 0x0
    "00000000", -- 4809 - 0x12c9  :    0 - 0x0
    "00000000", -- 4810 - 0x12ca  :    0 - 0x0
    "00000000", -- 4811 - 0x12cb  :    0 - 0x0
    "00000000", -- 4812 - 0x12cc  :    0 - 0x0
    "00000000", -- 4813 - 0x12cd  :    0 - 0x0
    "00001100", -- 4814 - 0x12ce  :   12 - 0xc
    "00011110", -- 4815 - 0x12cf  :   30 - 0x1e
    "00000000", -- 4816 - 0x12d0  :    0 - 0x0 -- Background 0x2d
    "00000000", -- 4817 - 0x12d1  :    0 - 0x0
    "00000000", -- 4818 - 0x12d2  :    0 - 0x0
    "00000000", -- 4819 - 0x12d3  :    0 - 0x0
    "00000000", -- 4820 - 0x12d4  :    0 - 0x0
    "00000000", -- 4821 - 0x12d5  :    0 - 0x0
    "00000000", -- 4822 - 0x12d6  :    0 - 0x0
    "00000000", -- 4823 - 0x12d7  :    0 - 0x0
    "00010010", -- 4824 - 0x12d8  :   18 - 0x12
    "00010010", -- 4825 - 0x12d9  :   18 - 0x12
    "00001100", -- 4826 - 0x12da  :   12 - 0xc
    "00000000", -- 4827 - 0x12db  :    0 - 0x0
    "00000000", -- 4828 - 0x12dc  :    0 - 0x0
    "00000000", -- 4829 - 0x12dd  :    0 - 0x0
    "00000000", -- 4830 - 0x12de  :    0 - 0x0
    "00000000", -- 4831 - 0x12df  :    0 - 0x0
    "00000000", -- 4832 - 0x12e0  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 4833 - 0x12e1  :    0 - 0x0
    "00000000", -- 4834 - 0x12e2  :    0 - 0x0
    "00000000", -- 4835 - 0x12e3  :    0 - 0x0
    "00000000", -- 4836 - 0x12e4  :    0 - 0x0
    "00000000", -- 4837 - 0x12e5  :    0 - 0x0
    "00000000", -- 4838 - 0x12e6  :    0 - 0x0
    "00000000", -- 4839 - 0x12e7  :    0 - 0x0
    "00000000", -- 4840 - 0x12e8  :    0 - 0x0
    "00000000", -- 4841 - 0x12e9  :    0 - 0x0
    "00000000", -- 4842 - 0x12ea  :    0 - 0x0
    "00010001", -- 4843 - 0x12eb  :   17 - 0x11
    "00110010", -- 4844 - 0x12ec  :   50 - 0x32
    "00010010", -- 4845 - 0x12ed  :   18 - 0x12
    "00010010", -- 4846 - 0x12ee  :   18 - 0x12
    "00010010", -- 4847 - 0x12ef  :   18 - 0x12
    "00000000", -- 4848 - 0x12f0  :    0 - 0x0 -- Background 0x2f
    "00000000", -- 4849 - 0x12f1  :    0 - 0x0
    "00000000", -- 4850 - 0x12f2  :    0 - 0x0
    "00000000", -- 4851 - 0x12f3  :    0 - 0x0
    "00000000", -- 4852 - 0x12f4  :    0 - 0x0
    "00000000", -- 4853 - 0x12f5  :    0 - 0x0
    "00000000", -- 4854 - 0x12f6  :    0 - 0x0
    "00000000", -- 4855 - 0x12f7  :    0 - 0x0
    "00000000", -- 4856 - 0x12f8  :    0 - 0x0
    "00000000", -- 4857 - 0x12f9  :    0 - 0x0
    "00000000", -- 4858 - 0x12fa  :    0 - 0x0
    "10001100", -- 4859 - 0x12fb  :  140 - 0x8c
    "01010010", -- 4860 - 0x12fc  :   82 - 0x52
    "01010010", -- 4861 - 0x12fd  :   82 - 0x52
    "01010010", -- 4862 - 0x12fe  :   82 - 0x52
    "01010010", -- 4863 - 0x12ff  :   82 - 0x52
    "00000000", -- 4864 - 0x1300  :    0 - 0x0 -- Background 0x30
    "00000000", -- 4865 - 0x1301  :    0 - 0x0
    "00000000", -- 4866 - 0x1302  :    0 - 0x0
    "00000000", -- 4867 - 0x1303  :    0 - 0x0
    "00000000", -- 4868 - 0x1304  :    0 - 0x0
    "00000000", -- 4869 - 0x1305  :    0 - 0x0
    "00000000", -- 4870 - 0x1306  :    0 - 0x0
    "00000000", -- 4871 - 0x1307  :    0 - 0x0
    "00010010", -- 4872 - 0x1308  :   18 - 0x12
    "00111001", -- 4873 - 0x1309  :   57 - 0x39
    "00000000", -- 4874 - 0x130a  :    0 - 0x0
    "00000000", -- 4875 - 0x130b  :    0 - 0x0
    "00000000", -- 4876 - 0x130c  :    0 - 0x0
    "00000000", -- 4877 - 0x130d  :    0 - 0x0
    "00000000", -- 4878 - 0x130e  :    0 - 0x0
    "00000000", -- 4879 - 0x130f  :    0 - 0x0
    "00000000", -- 4880 - 0x1310  :    0 - 0x0 -- Background 0x31
    "00000000", -- 4881 - 0x1311  :    0 - 0x0
    "00000000", -- 4882 - 0x1312  :    0 - 0x0
    "00000000", -- 4883 - 0x1313  :    0 - 0x0
    "00000000", -- 4884 - 0x1314  :    0 - 0x0
    "00000000", -- 4885 - 0x1315  :    0 - 0x0
    "00000000", -- 4886 - 0x1316  :    0 - 0x0
    "00000000", -- 4887 - 0x1317  :    0 - 0x0
    "01010010", -- 4888 - 0x1318  :   82 - 0x52
    "10001100", -- 4889 - 0x1319  :  140 - 0x8c
    "00000000", -- 4890 - 0x131a  :    0 - 0x0
    "00000000", -- 4891 - 0x131b  :    0 - 0x0
    "00000000", -- 4892 - 0x131c  :    0 - 0x0
    "00000000", -- 4893 - 0x131d  :    0 - 0x0
    "00000000", -- 4894 - 0x131e  :    0 - 0x0
    "00000000", -- 4895 - 0x131f  :    0 - 0x0
    "00000000", -- 4896 - 0x1320  :    0 - 0x0 -- Background 0x32
    "00000000", -- 4897 - 0x1321  :    0 - 0x0
    "00000000", -- 4898 - 0x1322  :    0 - 0x0
    "00000000", -- 4899 - 0x1323  :    0 - 0x0
    "00000000", -- 4900 - 0x1324  :    0 - 0x0
    "00000000", -- 4901 - 0x1325  :    0 - 0x0
    "00000000", -- 4902 - 0x1326  :    0 - 0x0
    "00000000", -- 4903 - 0x1327  :    0 - 0x0
    "00000000", -- 4904 - 0x1328  :    0 - 0x0
    "00000000", -- 4905 - 0x1329  :    0 - 0x0
    "00000000", -- 4906 - 0x132a  :    0 - 0x0
    "01110001", -- 4907 - 0x132b  :  113 - 0x71
    "10001010", -- 4908 - 0x132c  :  138 - 0x8a
    "00001010", -- 4909 - 0x132d  :   10 - 0xa
    "00010010", -- 4910 - 0x132e  :   18 - 0x12
    "00100010", -- 4911 - 0x132f  :   34 - 0x22
    "00000000", -- 4912 - 0x1330  :    0 - 0x0 -- Background 0x33
    "00000000", -- 4913 - 0x1331  :    0 - 0x0
    "00000000", -- 4914 - 0x1332  :    0 - 0x0
    "00000000", -- 4915 - 0x1333  :    0 - 0x0
    "00000000", -- 4916 - 0x1334  :    0 - 0x0
    "00000000", -- 4917 - 0x1335  :    0 - 0x0
    "00000000", -- 4918 - 0x1336  :    0 - 0x0
    "00000000", -- 4919 - 0x1337  :    0 - 0x0
    "01000010", -- 4920 - 0x1338  :   66 - 0x42
    "11111001", -- 4921 - 0x1339  :  249 - 0xf9
    "00000000", -- 4922 - 0x133a  :    0 - 0x0
    "00000000", -- 4923 - 0x133b  :    0 - 0x0
    "00000000", -- 4924 - 0x133c  :    0 - 0x0
    "00000000", -- 4925 - 0x133d  :    0 - 0x0
    "00000000", -- 4926 - 0x133e  :    0 - 0x0
    "00000000", -- 4927 - 0x133f  :    0 - 0x0
    "00000000", -- 4928 - 0x1340  :    0 - 0x0 -- Background 0x34
    "00000000", -- 4929 - 0x1341  :    0 - 0x0
    "00000000", -- 4930 - 0x1342  :    0 - 0x0
    "00000000", -- 4931 - 0x1343  :    0 - 0x0
    "00000000", -- 4932 - 0x1344  :    0 - 0x0
    "00000000", -- 4933 - 0x1345  :    0 - 0x0
    "00000000", -- 4934 - 0x1346  :    0 - 0x0
    "00000000", -- 4935 - 0x1347  :    0 - 0x0
    "00000000", -- 4936 - 0x1348  :    0 - 0x0
    "00000000", -- 4937 - 0x1349  :    0 - 0x0
    "00000000", -- 4938 - 0x134a  :    0 - 0x0
    "00110001", -- 4939 - 0x134b  :   49 - 0x31
    "01001010", -- 4940 - 0x134c  :   74 - 0x4a
    "00001010", -- 4941 - 0x134d  :   10 - 0xa
    "00110010", -- 4942 - 0x134e  :   50 - 0x32
    "00001010", -- 4943 - 0x134f  :   10 - 0xa
    "00000000", -- 4944 - 0x1350  :    0 - 0x0 -- Background 0x35
    "00000000", -- 4945 - 0x1351  :    0 - 0x0
    "00000000", -- 4946 - 0x1352  :    0 - 0x0
    "00000000", -- 4947 - 0x1353  :    0 - 0x0
    "00000000", -- 4948 - 0x1354  :    0 - 0x0
    "00000000", -- 4949 - 0x1355  :    0 - 0x0
    "00000000", -- 4950 - 0x1356  :    0 - 0x0
    "00000000", -- 4951 - 0x1357  :    0 - 0x0
    "01001010", -- 4952 - 0x1358  :   74 - 0x4a
    "00110001", -- 4953 - 0x1359  :   49 - 0x31
    "00000000", -- 4954 - 0x135a  :    0 - 0x0
    "00000000", -- 4955 - 0x135b  :    0 - 0x0
    "00000000", -- 4956 - 0x135c  :    0 - 0x0
    "00000000", -- 4957 - 0x135d  :    0 - 0x0
    "00000000", -- 4958 - 0x135e  :    0 - 0x0
    "00000000", -- 4959 - 0x135f  :    0 - 0x0
    "00000000", -- 4960 - 0x1360  :    0 - 0x0 -- Background 0x36
    "00000000", -- 4961 - 0x1361  :    0 - 0x0
    "00000000", -- 4962 - 0x1362  :    0 - 0x0
    "00000000", -- 4963 - 0x1363  :    0 - 0x0
    "00000000", -- 4964 - 0x1364  :    0 - 0x0
    "00000000", -- 4965 - 0x1365  :    0 - 0x0
    "00000000", -- 4966 - 0x1366  :    0 - 0x0
    "00000000", -- 4967 - 0x1367  :    0 - 0x0
    "00000000", -- 4968 - 0x1368  :    0 - 0x0
    "00000000", -- 4969 - 0x1369  :    0 - 0x0
    "00000000", -- 4970 - 0x136a  :    0 - 0x0
    "00010001", -- 4971 - 0x136b  :   17 - 0x11
    "00110010", -- 4972 - 0x136c  :   50 - 0x32
    "01010010", -- 4973 - 0x136d  :   82 - 0x52
    "10010010", -- 4974 - 0x136e  :  146 - 0x92
    "11111010", -- 4975 - 0x136f  :  250 - 0xfa
    "00000000", -- 4976 - 0x1370  :    0 - 0x0 -- Background 0x37
    "00000000", -- 4977 - 0x1371  :    0 - 0x0
    "00000000", -- 4978 - 0x1372  :    0 - 0x0
    "00000000", -- 4979 - 0x1373  :    0 - 0x0
    "00000000", -- 4980 - 0x1374  :    0 - 0x0
    "00000000", -- 4981 - 0x1375  :    0 - 0x0
    "00000000", -- 4982 - 0x1376  :    0 - 0x0
    "00000000", -- 4983 - 0x1377  :    0 - 0x0
    "00010010", -- 4984 - 0x1378  :   18 - 0x12
    "00010001", -- 4985 - 0x1379  :   17 - 0x11
    "00000000", -- 4986 - 0x137a  :    0 - 0x0
    "00000000", -- 4987 - 0x137b  :    0 - 0x0
    "00000000", -- 4988 - 0x137c  :    0 - 0x0
    "00000000", -- 4989 - 0x137d  :    0 - 0x0
    "00000000", -- 4990 - 0x137e  :    0 - 0x0
    "00000000", -- 4991 - 0x137f  :    0 - 0x0
    "00000000", -- 4992 - 0x1380  :    0 - 0x0 -- Background 0x38
    "00000000", -- 4993 - 0x1381  :    0 - 0x0
    "00000000", -- 4994 - 0x1382  :    0 - 0x0
    "00000000", -- 4995 - 0x1383  :    0 - 0x0
    "00000000", -- 4996 - 0x1384  :    0 - 0x0
    "00000000", -- 4997 - 0x1385  :    0 - 0x0
    "00000000", -- 4998 - 0x1386  :    0 - 0x0
    "00000000", -- 4999 - 0x1387  :    0 - 0x0
    "00000000", -- 5000 - 0x1388  :    0 - 0x0
    "00000000", -- 5001 - 0x1389  :    0 - 0x0
    "00000000", -- 5002 - 0x138a  :    0 - 0x0
    "01110001", -- 5003 - 0x138b  :  113 - 0x71
    "01000010", -- 5004 - 0x138c  :   66 - 0x42
    "01000010", -- 5005 - 0x138d  :   66 - 0x42
    "01110010", -- 5006 - 0x138e  :  114 - 0x72
    "00001010", -- 5007 - 0x138f  :   10 - 0xa
    "00000000", -- 5008 - 0x1390  :    0 - 0x0 -- Background 0x39
    "00000000", -- 5009 - 0x1391  :    0 - 0x0
    "00000000", -- 5010 - 0x1392  :    0 - 0x0
    "00000000", -- 5011 - 0x1393  :    0 - 0x0
    "00000000", -- 5012 - 0x1394  :    0 - 0x0
    "00000000", -- 5013 - 0x1395  :    0 - 0x0
    "00000000", -- 5014 - 0x1396  :    0 - 0x0
    "00000000", -- 5015 - 0x1397  :    0 - 0x0
    "00001010", -- 5016 - 0x1398  :   10 - 0xa
    "01110001", -- 5017 - 0x1399  :  113 - 0x71
    "00000000", -- 5018 - 0x139a  :    0 - 0x0
    "00000000", -- 5019 - 0x139b  :    0 - 0x0
    "00000000", -- 5020 - 0x139c  :    0 - 0x0
    "00000000", -- 5021 - 0x139d  :    0 - 0x0
    "00000000", -- 5022 - 0x139e  :    0 - 0x0
    "00000000", -- 5023 - 0x139f  :    0 - 0x0
    "00000000", -- 5024 - 0x13a0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 5025 - 0x13a1  :    0 - 0x0
    "00000000", -- 5026 - 0x13a2  :    0 - 0x0
    "00000000", -- 5027 - 0x13a3  :    0 - 0x0
    "00000000", -- 5028 - 0x13a4  :    0 - 0x0
    "00000000", -- 5029 - 0x13a5  :    0 - 0x0
    "00000000", -- 5030 - 0x13a6  :    0 - 0x0
    "00000000", -- 5031 - 0x13a7  :    0 - 0x0
    "00000000", -- 5032 - 0x13a8  :    0 - 0x0
    "00000000", -- 5033 - 0x13a9  :    0 - 0x0
    "00000000", -- 5034 - 0x13aa  :    0 - 0x0
    "01110001", -- 5035 - 0x13ab  :  113 - 0x71
    "00001010", -- 5036 - 0x13ac  :   10 - 0xa
    "00010010", -- 5037 - 0x13ad  :   18 - 0x12
    "00010010", -- 5038 - 0x13ae  :   18 - 0x12
    "00100010", -- 5039 - 0x13af  :   34 - 0x22
    "00000000", -- 5040 - 0x13b0  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 5041 - 0x13b1  :    0 - 0x0
    "00000000", -- 5042 - 0x13b2  :    0 - 0x0
    "00000000", -- 5043 - 0x13b3  :    0 - 0x0
    "00000000", -- 5044 - 0x13b4  :    0 - 0x0
    "00000000", -- 5045 - 0x13b5  :    0 - 0x0
    "00000000", -- 5046 - 0x13b6  :    0 - 0x0
    "00000000", -- 5047 - 0x13b7  :    0 - 0x0
    "00100010", -- 5048 - 0x13b8  :   34 - 0x22
    "00100001", -- 5049 - 0x13b9  :   33 - 0x21
    "00000000", -- 5050 - 0x13ba  :    0 - 0x0
    "00000000", -- 5051 - 0x13bb  :    0 - 0x0
    "00000000", -- 5052 - 0x13bc  :    0 - 0x0
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "00000000", -- 5054 - 0x13be  :    0 - 0x0
    "00000000", -- 5055 - 0x13bf  :    0 - 0x0
    "00000000", -- 5056 - 0x13c0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 5057 - 0x13c1  :    0 - 0x0
    "00000000", -- 5058 - 0x13c2  :    0 - 0x0
    "00000000", -- 5059 - 0x13c3  :    0 - 0x0
    "00000000", -- 5060 - 0x13c4  :    0 - 0x0
    "00000000", -- 5061 - 0x13c5  :    0 - 0x0
    "00000000", -- 5062 - 0x13c6  :    0 - 0x0
    "00000000", -- 5063 - 0x13c7  :    0 - 0x0
    "00000000", -- 5064 - 0x13c8  :    0 - 0x0
    "00000000", -- 5065 - 0x13c9  :    0 - 0x0
    "00000000", -- 5066 - 0x13ca  :    0 - 0x0
    "01110001", -- 5067 - 0x13cb  :  113 - 0x71
    "10001010", -- 5068 - 0x13cc  :  138 - 0x8a
    "10001010", -- 5069 - 0x13cd  :  138 - 0x8a
    "01110010", -- 5070 - 0x13ce  :  114 - 0x72
    "10001010", -- 5071 - 0x13cf  :  138 - 0x8a
    "00000000", -- 5072 - 0x13d0  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 5073 - 0x13d1  :    0 - 0x0
    "00000000", -- 5074 - 0x13d2  :    0 - 0x0
    "00000000", -- 5075 - 0x13d3  :    0 - 0x0
    "00000000", -- 5076 - 0x13d4  :    0 - 0x0
    "00000000", -- 5077 - 0x13d5  :    0 - 0x0
    "00000000", -- 5078 - 0x13d6  :    0 - 0x0
    "00000000", -- 5079 - 0x13d7  :    0 - 0x0
    "10001010", -- 5080 - 0x13d8  :  138 - 0x8a
    "01110001", -- 5081 - 0x13d9  :  113 - 0x71
    "00000000", -- 5082 - 0x13da  :    0 - 0x0
    "00000000", -- 5083 - 0x13db  :    0 - 0x0
    "00000000", -- 5084 - 0x13dc  :    0 - 0x0
    "00000000", -- 5085 - 0x13dd  :    0 - 0x0
    "00000000", -- 5086 - 0x13de  :    0 - 0x0
    "00000000", -- 5087 - 0x13df  :    0 - 0x0
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 5089 - 0x13e1  :    0 - 0x0
    "00000000", -- 5090 - 0x13e2  :    0 - 0x0
    "00000000", -- 5091 - 0x13e3  :    0 - 0x0
    "00000000", -- 5092 - 0x13e4  :    0 - 0x0
    "00000000", -- 5093 - 0x13e5  :    0 - 0x0
    "00000000", -- 5094 - 0x13e6  :    0 - 0x0
    "00000000", -- 5095 - 0x13e7  :    0 - 0x0
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000000", -- 5097 - 0x13e9  :    0 - 0x0
    "00000000", -- 5098 - 0x13ea  :    0 - 0x0
    "10011000", -- 5099 - 0x13eb  :  152 - 0x98
    "10100101", -- 5100 - 0x13ec  :  165 - 0xa5
    "10100101", -- 5101 - 0x13ed  :  165 - 0xa5
    "10100101", -- 5102 - 0x13ee  :  165 - 0xa5
    "10100101", -- 5103 - 0x13ef  :  165 - 0xa5
    "00000000", -- 5104 - 0x13f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 5105 - 0x13f1  :    0 - 0x0
    "00000000", -- 5106 - 0x13f2  :    0 - 0x0
    "00000000", -- 5107 - 0x13f3  :    0 - 0x0
    "00000000", -- 5108 - 0x13f4  :    0 - 0x0
    "00000000", -- 5109 - 0x13f5  :    0 - 0x0
    "00000000", -- 5110 - 0x13f6  :    0 - 0x0
    "00000000", -- 5111 - 0x13f7  :    0 - 0x0
    "00000000", -- 5112 - 0x13f8  :    0 - 0x0
    "00000000", -- 5113 - 0x13f9  :    0 - 0x0
    "00000000", -- 5114 - 0x13fa  :    0 - 0x0
    "11000110", -- 5115 - 0x13fb  :  198 - 0xc6
    "00101001", -- 5116 - 0x13fc  :   41 - 0x29
    "00101001", -- 5117 - 0x13fd  :   41 - 0x29
    "00101001", -- 5118 - 0x13fe  :   41 - 0x29
    "00101001", -- 5119 - 0x13ff  :   41 - 0x29
    "00000000", -- 5120 - 0x1400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 5121 - 0x1401  :    0 - 0x0
    "00000000", -- 5122 - 0x1402  :    0 - 0x0
    "00000000", -- 5123 - 0x1403  :    0 - 0x0
    "00000000", -- 5124 - 0x1404  :    0 - 0x0
    "00000000", -- 5125 - 0x1405  :    0 - 0x0
    "00000000", -- 5126 - 0x1406  :    0 - 0x0
    "00000000", -- 5127 - 0x1407  :    0 - 0x0
    "10100101", -- 5128 - 0x1408  :  165 - 0xa5
    "10011000", -- 5129 - 0x1409  :  152 - 0x98
    "00000000", -- 5130 - 0x140a  :    0 - 0x0
    "00000000", -- 5131 - 0x140b  :    0 - 0x0
    "00000000", -- 5132 - 0x140c  :    0 - 0x0
    "00000000", -- 5133 - 0x140d  :    0 - 0x0
    "00000000", -- 5134 - 0x140e  :    0 - 0x0
    "00000000", -- 5135 - 0x140f  :    0 - 0x0
    "00000000", -- 5136 - 0x1410  :    0 - 0x0 -- Background 0x41
    "00000000", -- 5137 - 0x1411  :    0 - 0x0
    "00000000", -- 5138 - 0x1412  :    0 - 0x0
    "00000000", -- 5139 - 0x1413  :    0 - 0x0
    "00000000", -- 5140 - 0x1414  :    0 - 0x0
    "00000000", -- 5141 - 0x1415  :    0 - 0x0
    "00000000", -- 5142 - 0x1416  :    0 - 0x0
    "00000000", -- 5143 - 0x1417  :    0 - 0x0
    "00101001", -- 5144 - 0x1418  :   41 - 0x29
    "11000110", -- 5145 - 0x1419  :  198 - 0xc6
    "00000000", -- 5146 - 0x141a  :    0 - 0x0
    "00000000", -- 5147 - 0x141b  :    0 - 0x0
    "00000000", -- 5148 - 0x141c  :    0 - 0x0
    "00000000", -- 5149 - 0x141d  :    0 - 0x0
    "00000000", -- 5150 - 0x141e  :    0 - 0x0
    "00000000", -- 5151 - 0x141f  :    0 - 0x0
    "00000000", -- 5152 - 0x1420  :    0 - 0x0 -- Background 0x42
    "00000000", -- 5153 - 0x1421  :    0 - 0x0
    "00000000", -- 5154 - 0x1422  :    0 - 0x0
    "00000000", -- 5155 - 0x1423  :    0 - 0x0
    "00000000", -- 5156 - 0x1424  :    0 - 0x0
    "00000000", -- 5157 - 0x1425  :    0 - 0x0
    "00000000", -- 5158 - 0x1426  :    0 - 0x0
    "00000000", -- 5159 - 0x1427  :    0 - 0x0
    "00000000", -- 5160 - 0x1428  :    0 - 0x0
    "00000000", -- 5161 - 0x1429  :    0 - 0x0
    "00000000", -- 5162 - 0x142a  :    0 - 0x0
    "10011100", -- 5163 - 0x142b  :  156 - 0x9c
    "10100001", -- 5164 - 0x142c  :  161 - 0xa1
    "10100001", -- 5165 - 0x142d  :  161 - 0xa1
    "10111101", -- 5166 - 0x142e  :  189 - 0xbd
    "10100101", -- 5167 - 0x142f  :  165 - 0xa5
    "00000000", -- 5168 - 0x1430  :    0 - 0x0 -- Background 0x43
    "00000000", -- 5169 - 0x1431  :    0 - 0x0
    "00000000", -- 5170 - 0x1432  :    0 - 0x0
    "00000000", -- 5171 - 0x1433  :    0 - 0x0
    "00000000", -- 5172 - 0x1434  :    0 - 0x0
    "00000000", -- 5173 - 0x1435  :    0 - 0x0
    "00000000", -- 5174 - 0x1436  :    0 - 0x0
    "00000000", -- 5175 - 0x1437  :    0 - 0x0
    "10100101", -- 5176 - 0x1438  :  165 - 0xa5
    "10011000", -- 5177 - 0x1439  :  152 - 0x98
    "00000000", -- 5178 - 0x143a  :    0 - 0x0
    "00000000", -- 5179 - 0x143b  :    0 - 0x0
    "00000000", -- 5180 - 0x143c  :    0 - 0x0
    "00000000", -- 5181 - 0x143d  :    0 - 0x0
    "00000000", -- 5182 - 0x143e  :    0 - 0x0
    "00000000", -- 5183 - 0x143f  :    0 - 0x0
    "00000000", -- 5184 - 0x1440  :    0 - 0x0 -- Background 0x44
    "00000000", -- 5185 - 0x1441  :    0 - 0x0
    "00000000", -- 5186 - 0x1442  :    0 - 0x0
    "00000000", -- 5187 - 0x1443  :    0 - 0x0
    "00000000", -- 5188 - 0x1444  :    0 - 0x0
    "00000000", -- 5189 - 0x1445  :    0 - 0x0
    "00000000", -- 5190 - 0x1446  :    0 - 0x0
    "00000000", -- 5191 - 0x1447  :    0 - 0x0
    "00000000", -- 5192 - 0x1448  :    0 - 0x0
    "00000000", -- 5193 - 0x1449  :    0 - 0x0
    "00000000", -- 5194 - 0x144a  :    0 - 0x0
    "01100010", -- 5195 - 0x144b  :   98 - 0x62
    "10010101", -- 5196 - 0x144c  :  149 - 0x95
    "00010101", -- 5197 - 0x144d  :   21 - 0x15
    "00100101", -- 5198 - 0x144e  :   37 - 0x25
    "01000101", -- 5199 - 0x144f  :   69 - 0x45
    "00000000", -- 5200 - 0x1450  :    0 - 0x0 -- Background 0x45
    "00000000", -- 5201 - 0x1451  :    0 - 0x0
    "00000000", -- 5202 - 0x1452  :    0 - 0x0
    "00000000", -- 5203 - 0x1453  :    0 - 0x0
    "00000000", -- 5204 - 0x1454  :    0 - 0x0
    "00000000", -- 5205 - 0x1455  :    0 - 0x0
    "00000000", -- 5206 - 0x1456  :    0 - 0x0
    "00000000", -- 5207 - 0x1457  :    0 - 0x0
    "00000000", -- 5208 - 0x1458  :    0 - 0x0
    "00000000", -- 5209 - 0x1459  :    0 - 0x0
    "00000000", -- 5210 - 0x145a  :    0 - 0x0
    "00100010", -- 5211 - 0x145b  :   34 - 0x22
    "01010101", -- 5212 - 0x145c  :   85 - 0x55
    "01010101", -- 5213 - 0x145d  :   85 - 0x55
    "01010101", -- 5214 - 0x145e  :   85 - 0x55
    "01010101", -- 5215 - 0x145f  :   85 - 0x55
    "00000000", -- 5216 - 0x1460  :    0 - 0x0 -- Background 0x46
    "00000000", -- 5217 - 0x1461  :    0 - 0x0
    "00000000", -- 5218 - 0x1462  :    0 - 0x0
    "00000000", -- 5219 - 0x1463  :    0 - 0x0
    "00000000", -- 5220 - 0x1464  :    0 - 0x0
    "00000000", -- 5221 - 0x1465  :    0 - 0x0
    "00000000", -- 5222 - 0x1466  :    0 - 0x0
    "00000000", -- 5223 - 0x1467  :    0 - 0x0
    "10000101", -- 5224 - 0x1468  :  133 - 0x85
    "11110010", -- 5225 - 0x1469  :  242 - 0xf2
    "00000000", -- 5226 - 0x146a  :    0 - 0x0
    "00000000", -- 5227 - 0x146b  :    0 - 0x0
    "00000000", -- 5228 - 0x146c  :    0 - 0x0
    "00000000", -- 5229 - 0x146d  :    0 - 0x0
    "00000000", -- 5230 - 0x146e  :    0 - 0x0
    "00000000", -- 5231 - 0x146f  :    0 - 0x0
    "00000000", -- 5232 - 0x1470  :    0 - 0x0 -- Background 0x47
    "00000000", -- 5233 - 0x1471  :    0 - 0x0
    "00000000", -- 5234 - 0x1472  :    0 - 0x0
    "00000000", -- 5235 - 0x1473  :    0 - 0x0
    "00000000", -- 5236 - 0x1474  :    0 - 0x0
    "00000000", -- 5237 - 0x1475  :    0 - 0x0
    "00000000", -- 5238 - 0x1476  :    0 - 0x0
    "00000000", -- 5239 - 0x1477  :    0 - 0x0
    "01010101", -- 5240 - 0x1478  :   85 - 0x55
    "00100010", -- 5241 - 0x1479  :   34 - 0x22
    "00000000", -- 5242 - 0x147a  :    0 - 0x0
    "00000000", -- 5243 - 0x147b  :    0 - 0x0
    "00000000", -- 5244 - 0x147c  :    0 - 0x0
    "00000000", -- 5245 - 0x147d  :    0 - 0x0
    "00000000", -- 5246 - 0x147e  :    0 - 0x0
    "00000000", -- 5247 - 0x147f  :    0 - 0x0
    "00000000", -- 5248 - 0x1480  :    0 - 0x0 -- Background 0x48
    "00000000", -- 5249 - 0x1481  :    0 - 0x0
    "00000000", -- 5250 - 0x1482  :    0 - 0x0
    "00000000", -- 5251 - 0x1483  :    0 - 0x0
    "00000000", -- 5252 - 0x1484  :    0 - 0x0
    "00000000", -- 5253 - 0x1485  :    0 - 0x0
    "00000000", -- 5254 - 0x1486  :    0 - 0x0
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "00000000", -- 5257 - 0x1489  :    0 - 0x0
    "00000000", -- 5258 - 0x148a  :    0 - 0x0
    "01100010", -- 5259 - 0x148b  :   98 - 0x62
    "10010101", -- 5260 - 0x148c  :  149 - 0x95
    "00010101", -- 5261 - 0x148d  :   21 - 0x15
    "01100101", -- 5262 - 0x148e  :  101 - 0x65
    "00010101", -- 5263 - 0x148f  :   21 - 0x15
    "00000000", -- 5264 - 0x1490  :    0 - 0x0 -- Background 0x49
    "00000000", -- 5265 - 0x1491  :    0 - 0x0
    "00000000", -- 5266 - 0x1492  :    0 - 0x0
    "00000000", -- 5267 - 0x1493  :    0 - 0x0
    "00000000", -- 5268 - 0x1494  :    0 - 0x0
    "00000000", -- 5269 - 0x1495  :    0 - 0x0
    "00000000", -- 5270 - 0x1496  :    0 - 0x0
    "00000000", -- 5271 - 0x1497  :    0 - 0x0
    "10010101", -- 5272 - 0x1498  :  149 - 0x95
    "01100010", -- 5273 - 0x1499  :   98 - 0x62
    "00000000", -- 5274 - 0x149a  :    0 - 0x0
    "00000000", -- 5275 - 0x149b  :    0 - 0x0
    "00000000", -- 5276 - 0x149c  :    0 - 0x0
    "00000000", -- 5277 - 0x149d  :    0 - 0x0
    "00000000", -- 5278 - 0x149e  :    0 - 0x0
    "00000000", -- 5279 - 0x149f  :    0 - 0x0
    "00000000", -- 5280 - 0x14a0  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 5281 - 0x14a1  :    0 - 0x0
    "00000000", -- 5282 - 0x14a2  :    0 - 0x0
    "00000000", -- 5283 - 0x14a3  :    0 - 0x0
    "00000000", -- 5284 - 0x14a4  :    0 - 0x0
    "00000000", -- 5285 - 0x14a5  :    0 - 0x0
    "00000000", -- 5286 - 0x14a6  :    0 - 0x0
    "00000000", -- 5287 - 0x14a7  :    0 - 0x0
    "00000000", -- 5288 - 0x14a8  :    0 - 0x0
    "00000000", -- 5289 - 0x14a9  :    0 - 0x0
    "00000000", -- 5290 - 0x14aa  :    0 - 0x0
    "11100010", -- 5291 - 0x14ab  :  226 - 0xe2
    "10000101", -- 5292 - 0x14ac  :  133 - 0x85
    "10000101", -- 5293 - 0x14ad  :  133 - 0x85
    "11100101", -- 5294 - 0x14ae  :  229 - 0xe5
    "00010101", -- 5295 - 0x14af  :   21 - 0x15
    "00000000", -- 5296 - 0x14b0  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 5297 - 0x14b1  :    0 - 0x0
    "00000000", -- 5298 - 0x14b2  :    0 - 0x0
    "00000000", -- 5299 - 0x14b3  :    0 - 0x0
    "00000000", -- 5300 - 0x14b4  :    0 - 0x0
    "00000000", -- 5301 - 0x14b5  :    0 - 0x0
    "00000000", -- 5302 - 0x14b6  :    0 - 0x0
    "00000000", -- 5303 - 0x14b7  :    0 - 0x0
    "00010101", -- 5304 - 0x14b8  :   21 - 0x15
    "11100010", -- 5305 - 0x14b9  :  226 - 0xe2
    "00000000", -- 5306 - 0x14ba  :    0 - 0x0
    "00000000", -- 5307 - 0x14bb  :    0 - 0x0
    "00000000", -- 5308 - 0x14bc  :    0 - 0x0
    "00000000", -- 5309 - 0x14bd  :    0 - 0x0
    "00000000", -- 5310 - 0x14be  :    0 - 0x0
    "00000000", -- 5311 - 0x14bf  :    0 - 0x0
    "00000000", -- 5312 - 0x14c0  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 5313 - 0x14c1  :    0 - 0x0
    "00000000", -- 5314 - 0x14c2  :    0 - 0x0
    "00000000", -- 5315 - 0x14c3  :    0 - 0x0
    "00000000", -- 5316 - 0x14c4  :    0 - 0x0
    "00000000", -- 5317 - 0x14c5  :    0 - 0x0
    "00000000", -- 5318 - 0x14c6  :    0 - 0x0
    "00000000", -- 5319 - 0x14c7  :    0 - 0x0
    "00000000", -- 5320 - 0x14c8  :    0 - 0x0
    "00000000", -- 5321 - 0x14c9  :    0 - 0x0
    "00000000", -- 5322 - 0x14ca  :    0 - 0x0
    "00000000", -- 5323 - 0x14cb  :    0 - 0x0
    "00000000", -- 5324 - 0x14cc  :    0 - 0x0
    "00000000", -- 5325 - 0x14cd  :    0 - 0x0
    "00000000", -- 5326 - 0x14ce  :    0 - 0x0
    "00000000", -- 5327 - 0x14cf  :    0 - 0x0
    "00000000", -- 5328 - 0x14d0  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 5329 - 0x14d1  :    0 - 0x0
    "00000000", -- 5330 - 0x14d2  :    0 - 0x0
    "00000001", -- 5331 - 0x14d3  :    1 - 0x1
    "00000011", -- 5332 - 0x14d4  :    3 - 0x3
    "00000111", -- 5333 - 0x14d5  :    7 - 0x7
    "00001111", -- 5334 - 0x14d6  :   15 - 0xf
    "00011111", -- 5335 - 0x14d7  :   31 - 0x1f
    "00000000", -- 5336 - 0x14d8  :    0 - 0x0
    "00000000", -- 5337 - 0x14d9  :    0 - 0x0
    "00000000", -- 5338 - 0x14da  :    0 - 0x0
    "00000000", -- 5339 - 0x14db  :    0 - 0x0
    "00000000", -- 5340 - 0x14dc  :    0 - 0x0
    "00000000", -- 5341 - 0x14dd  :    0 - 0x0
    "00000000", -- 5342 - 0x14de  :    0 - 0x0
    "00000000", -- 5343 - 0x14df  :    0 - 0x0
    "00000000", -- 5344 - 0x14e0  :    0 - 0x0 -- Background 0x4e
    "00001111", -- 5345 - 0x14e1  :   15 - 0xf
    "01111111", -- 5346 - 0x14e2  :  127 - 0x7f
    "11111111", -- 5347 - 0x14e3  :  255 - 0xff
    "11111111", -- 5348 - 0x14e4  :  255 - 0xff
    "11111111", -- 5349 - 0x14e5  :  255 - 0xff
    "11111111", -- 5350 - 0x14e6  :  255 - 0xff
    "11111111", -- 5351 - 0x14e7  :  255 - 0xff
    "00000000", -- 5352 - 0x14e8  :    0 - 0x0
    "00000000", -- 5353 - 0x14e9  :    0 - 0x0
    "00000000", -- 5354 - 0x14ea  :    0 - 0x0
    "00000000", -- 5355 - 0x14eb  :    0 - 0x0
    "00000000", -- 5356 - 0x14ec  :    0 - 0x0
    "00000000", -- 5357 - 0x14ed  :    0 - 0x0
    "00000000", -- 5358 - 0x14ee  :    0 - 0x0
    "00000000", -- 5359 - 0x14ef  :    0 - 0x0
    "00011111", -- 5360 - 0x14f0  :   31 - 0x1f -- Background 0x4f
    "00111111", -- 5361 - 0x14f1  :   63 - 0x3f
    "00111111", -- 5362 - 0x14f2  :   63 - 0x3f
    "00111111", -- 5363 - 0x14f3  :   63 - 0x3f
    "01111111", -- 5364 - 0x14f4  :  127 - 0x7f
    "01111111", -- 5365 - 0x14f5  :  127 - 0x7f
    "01111111", -- 5366 - 0x14f6  :  127 - 0x7f
    "01111111", -- 5367 - 0x14f7  :  127 - 0x7f
    "00000000", -- 5368 - 0x14f8  :    0 - 0x0
    "00000000", -- 5369 - 0x14f9  :    0 - 0x0
    "00000000", -- 5370 - 0x14fa  :    0 - 0x0
    "00000000", -- 5371 - 0x14fb  :    0 - 0x0
    "00000000", -- 5372 - 0x14fc  :    0 - 0x0
    "00000000", -- 5373 - 0x14fd  :    0 - 0x0
    "00000000", -- 5374 - 0x14fe  :    0 - 0x0
    "00000000", -- 5375 - 0x14ff  :    0 - 0x0
    "11111111", -- 5376 - 0x1500  :  255 - 0xff -- Background 0x50
    "11111111", -- 5377 - 0x1501  :  255 - 0xff
    "11111111", -- 5378 - 0x1502  :  255 - 0xff
    "11111111", -- 5379 - 0x1503  :  255 - 0xff
    "11111111", -- 5380 - 0x1504  :  255 - 0xff
    "11111111", -- 5381 - 0x1505  :  255 - 0xff
    "11111111", -- 5382 - 0x1506  :  255 - 0xff
    "11111111", -- 5383 - 0x1507  :  255 - 0xff
    "00000000", -- 5384 - 0x1508  :    0 - 0x0
    "00000000", -- 5385 - 0x1509  :    0 - 0x0
    "00000000", -- 5386 - 0x150a  :    0 - 0x0
    "00000000", -- 5387 - 0x150b  :    0 - 0x0
    "00000000", -- 5388 - 0x150c  :    0 - 0x0
    "00000000", -- 5389 - 0x150d  :    0 - 0x0
    "00000000", -- 5390 - 0x150e  :    0 - 0x0
    "00000000", -- 5391 - 0x150f  :    0 - 0x0
    "11111111", -- 5392 - 0x1510  :  255 - 0xff -- Background 0x51
    "11111111", -- 5393 - 0x1511  :  255 - 0xff
    "11111111", -- 5394 - 0x1512  :  255 - 0xff
    "11111111", -- 5395 - 0x1513  :  255 - 0xff
    "11111111", -- 5396 - 0x1514  :  255 - 0xff
    "11111111", -- 5397 - 0x1515  :  255 - 0xff
    "11111111", -- 5398 - 0x1516  :  255 - 0xff
    "11111110", -- 5399 - 0x1517  :  254 - 0xfe
    "00000000", -- 5400 - 0x1518  :    0 - 0x0
    "00000000", -- 5401 - 0x1519  :    0 - 0x0
    "00000000", -- 5402 - 0x151a  :    0 - 0x0
    "00000000", -- 5403 - 0x151b  :    0 - 0x0
    "00000000", -- 5404 - 0x151c  :    0 - 0x0
    "00000000", -- 5405 - 0x151d  :    0 - 0x0
    "00000000", -- 5406 - 0x151e  :    0 - 0x0
    "00000000", -- 5407 - 0x151f  :    0 - 0x0
    "00000000", -- 5408 - 0x1520  :    0 - 0x0 -- Background 0x52
    "00000000", -- 5409 - 0x1521  :    0 - 0x0
    "00000000", -- 5410 - 0x1522  :    0 - 0x0
    "10000000", -- 5411 - 0x1523  :  128 - 0x80
    "11000000", -- 5412 - 0x1524  :  192 - 0xc0
    "11100000", -- 5413 - 0x1525  :  224 - 0xe0
    "11110000", -- 5414 - 0x1526  :  240 - 0xf0
    "11110000", -- 5415 - 0x1527  :  240 - 0xf0
    "00000000", -- 5416 - 0x1528  :    0 - 0x0
    "00000000", -- 5417 - 0x1529  :    0 - 0x0
    "00000000", -- 5418 - 0x152a  :    0 - 0x0
    "00000000", -- 5419 - 0x152b  :    0 - 0x0
    "00000000", -- 5420 - 0x152c  :    0 - 0x0
    "00000000", -- 5421 - 0x152d  :    0 - 0x0
    "00000000", -- 5422 - 0x152e  :    0 - 0x0
    "00000000", -- 5423 - 0x152f  :    0 - 0x0
    "11111111", -- 5424 - 0x1530  :  255 - 0xff -- Background 0x53
    "11111111", -- 5425 - 0x1531  :  255 - 0xff
    "11111110", -- 5426 - 0x1532  :  254 - 0xfe
    "11111100", -- 5427 - 0x1533  :  252 - 0xfc
    "11110000", -- 5428 - 0x1534  :  240 - 0xf0
    "11100000", -- 5429 - 0x1535  :  224 - 0xe0
    "10000000", -- 5430 - 0x1536  :  128 - 0x80
    "00000000", -- 5431 - 0x1537  :    0 - 0x0
    "00000000", -- 5432 - 0x1538  :    0 - 0x0
    "00000000", -- 5433 - 0x1539  :    0 - 0x0
    "00000000", -- 5434 - 0x153a  :    0 - 0x0
    "00000000", -- 5435 - 0x153b  :    0 - 0x0
    "00000000", -- 5436 - 0x153c  :    0 - 0x0
    "00000000", -- 5437 - 0x153d  :    0 - 0x0
    "00000000", -- 5438 - 0x153e  :    0 - 0x0
    "00000000", -- 5439 - 0x153f  :    0 - 0x0
    "11000000", -- 5440 - 0x1540  :  192 - 0xc0 -- Background 0x54
    "10000000", -- 5441 - 0x1541  :  128 - 0x80
    "00000000", -- 5442 - 0x1542  :    0 - 0x0
    "00000000", -- 5443 - 0x1543  :    0 - 0x0
    "00000000", -- 5444 - 0x1544  :    0 - 0x0
    "00000000", -- 5445 - 0x1545  :    0 - 0x0
    "00000000", -- 5446 - 0x1546  :    0 - 0x0
    "00000000", -- 5447 - 0x1547  :    0 - 0x0
    "00000000", -- 5448 - 0x1548  :    0 - 0x0
    "00000000", -- 5449 - 0x1549  :    0 - 0x0
    "00000000", -- 5450 - 0x154a  :    0 - 0x0
    "00000000", -- 5451 - 0x154b  :    0 - 0x0
    "00000000", -- 5452 - 0x154c  :    0 - 0x0
    "00000000", -- 5453 - 0x154d  :    0 - 0x0
    "00000000", -- 5454 - 0x154e  :    0 - 0x0
    "00000000", -- 5455 - 0x154f  :    0 - 0x0
    "00000000", -- 5456 - 0x1550  :    0 - 0x0 -- Background 0x55
    "11110000", -- 5457 - 0x1551  :  240 - 0xf0
    "11111110", -- 5458 - 0x1552  :  254 - 0xfe
    "11111110", -- 5459 - 0x1553  :  254 - 0xfe
    "11111110", -- 5460 - 0x1554  :  254 - 0xfe
    "11111100", -- 5461 - 0x1555  :  252 - 0xfc
    "11111000", -- 5462 - 0x1556  :  248 - 0xf8
    "11111000", -- 5463 - 0x1557  :  248 - 0xf8
    "00000000", -- 5464 - 0x1558  :    0 - 0x0
    "00000000", -- 5465 - 0x1559  :    0 - 0x0
    "00000000", -- 5466 - 0x155a  :    0 - 0x0
    "00000000", -- 5467 - 0x155b  :    0 - 0x0
    "00000000", -- 5468 - 0x155c  :    0 - 0x0
    "00000000", -- 5469 - 0x155d  :    0 - 0x0
    "00000000", -- 5470 - 0x155e  :    0 - 0x0
    "00000000", -- 5471 - 0x155f  :    0 - 0x0
    "11110000", -- 5472 - 0x1560  :  240 - 0xf0 -- Background 0x56
    "11100000", -- 5473 - 0x1561  :  224 - 0xe0
    "11100000", -- 5474 - 0x1562  :  224 - 0xe0
    "11000000", -- 5475 - 0x1563  :  192 - 0xc0
    "10000000", -- 5476 - 0x1564  :  128 - 0x80
    "10000000", -- 5477 - 0x1565  :  128 - 0x80
    "00000000", -- 5478 - 0x1566  :    0 - 0x0
    "00000000", -- 5479 - 0x1567  :    0 - 0x0
    "00000000", -- 5480 - 0x1568  :    0 - 0x0
    "00000000", -- 5481 - 0x1569  :    0 - 0x0
    "00000000", -- 5482 - 0x156a  :    0 - 0x0
    "00000000", -- 5483 - 0x156b  :    0 - 0x0
    "00000000", -- 5484 - 0x156c  :    0 - 0x0
    "00000000", -- 5485 - 0x156d  :    0 - 0x0
    "00000000", -- 5486 - 0x156e  :    0 - 0x0
    "00000000", -- 5487 - 0x156f  :    0 - 0x0
    "00000000", -- 5488 - 0x1570  :    0 - 0x0 -- Background 0x57
    "00000000", -- 5489 - 0x1571  :    0 - 0x0
    "00000000", -- 5490 - 0x1572  :    0 - 0x0
    "00000000", -- 5491 - 0x1573  :    0 - 0x0
    "00000000", -- 5492 - 0x1574  :    0 - 0x0
    "00000000", -- 5493 - 0x1575  :    0 - 0x0
    "00000000", -- 5494 - 0x1576  :    0 - 0x0
    "00000100", -- 5495 - 0x1577  :    4 - 0x4
    "00000000", -- 5496 - 0x1578  :    0 - 0x0
    "00000000", -- 5497 - 0x1579  :    0 - 0x0
    "00000000", -- 5498 - 0x157a  :    0 - 0x0
    "00000000", -- 5499 - 0x157b  :    0 - 0x0
    "00000000", -- 5500 - 0x157c  :    0 - 0x0
    "00000000", -- 5501 - 0x157d  :    0 - 0x0
    "00000000", -- 5502 - 0x157e  :    0 - 0x0
    "00000100", -- 5503 - 0x157f  :    4 - 0x4
    "00000110", -- 5504 - 0x1580  :    6 - 0x6 -- Background 0x58
    "00000110", -- 5505 - 0x1581  :    6 - 0x6
    "00000111", -- 5506 - 0x1582  :    7 - 0x7
    "00000111", -- 5507 - 0x1583  :    7 - 0x7
    "00000111", -- 5508 - 0x1584  :    7 - 0x7
    "00000111", -- 5509 - 0x1585  :    7 - 0x7
    "00000000", -- 5510 - 0x1586  :    0 - 0x0
    "00000000", -- 5511 - 0x1587  :    0 - 0x0
    "00000110", -- 5512 - 0x1588  :    6 - 0x6
    "00000110", -- 5513 - 0x1589  :    6 - 0x6
    "00000111", -- 5514 - 0x158a  :    7 - 0x7
    "00000111", -- 5515 - 0x158b  :    7 - 0x7
    "00000111", -- 5516 - 0x158c  :    7 - 0x7
    "00000111", -- 5517 - 0x158d  :    7 - 0x7
    "00000000", -- 5518 - 0x158e  :    0 - 0x0
    "00000000", -- 5519 - 0x158f  :    0 - 0x0
    "00000000", -- 5520 - 0x1590  :    0 - 0x0 -- Background 0x59
    "00000000", -- 5521 - 0x1591  :    0 - 0x0
    "00000000", -- 5522 - 0x1592  :    0 - 0x0
    "00000000", -- 5523 - 0x1593  :    0 - 0x0
    "00000000", -- 5524 - 0x1594  :    0 - 0x0
    "00000000", -- 5525 - 0x1595  :    0 - 0x0
    "00000000", -- 5526 - 0x1596  :    0 - 0x0
    "00010000", -- 5527 - 0x1597  :   16 - 0x10
    "00000000", -- 5528 - 0x1598  :    0 - 0x0
    "00000000", -- 5529 - 0x1599  :    0 - 0x0
    "00000000", -- 5530 - 0x159a  :    0 - 0x0
    "00000000", -- 5531 - 0x159b  :    0 - 0x0
    "00000000", -- 5532 - 0x159c  :    0 - 0x0
    "00000000", -- 5533 - 0x159d  :    0 - 0x0
    "00000000", -- 5534 - 0x159e  :    0 - 0x0
    "00010000", -- 5535 - 0x159f  :   16 - 0x10
    "00011100", -- 5536 - 0x15a0  :   28 - 0x1c -- Background 0x5a
    "00011110", -- 5537 - 0x15a1  :   30 - 0x1e
    "00011111", -- 5538 - 0x15a2  :   31 - 0x1f
    "00011111", -- 5539 - 0x15a3  :   31 - 0x1f
    "00011111", -- 5540 - 0x15a4  :   31 - 0x1f
    "00011111", -- 5541 - 0x15a5  :   31 - 0x1f
    "00000000", -- 5542 - 0x15a6  :    0 - 0x0
    "00000000", -- 5543 - 0x15a7  :    0 - 0x0
    "00011100", -- 5544 - 0x15a8  :   28 - 0x1c
    "00011110", -- 5545 - 0x15a9  :   30 - 0x1e
    "00011111", -- 5546 - 0x15aa  :   31 - 0x1f
    "00011111", -- 5547 - 0x15ab  :   31 - 0x1f
    "00011111", -- 5548 - 0x15ac  :   31 - 0x1f
    "00011111", -- 5549 - 0x15ad  :   31 - 0x1f
    "00000000", -- 5550 - 0x15ae  :    0 - 0x0
    "00000000", -- 5551 - 0x15af  :    0 - 0x0
    "00000000", -- 5552 - 0x15b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 5553 - 0x15b1  :    0 - 0x0
    "00000000", -- 5554 - 0x15b2  :    0 - 0x0
    "00000000", -- 5555 - 0x15b3  :    0 - 0x0
    "00000000", -- 5556 - 0x15b4  :    0 - 0x0
    "00000000", -- 5557 - 0x15b5  :    0 - 0x0
    "00000000", -- 5558 - 0x15b6  :    0 - 0x0
    "11000000", -- 5559 - 0x15b7  :  192 - 0xc0
    "00000000", -- 5560 - 0x15b8  :    0 - 0x0
    "00000000", -- 5561 - 0x15b9  :    0 - 0x0
    "00000000", -- 5562 - 0x15ba  :    0 - 0x0
    "00000000", -- 5563 - 0x15bb  :    0 - 0x0
    "00000000", -- 5564 - 0x15bc  :    0 - 0x0
    "00000000", -- 5565 - 0x15bd  :    0 - 0x0
    "00000000", -- 5566 - 0x15be  :    0 - 0x0
    "11000000", -- 5567 - 0x15bf  :  192 - 0xc0
    "11110000", -- 5568 - 0x15c0  :  240 - 0xf0 -- Background 0x5c
    "11111100", -- 5569 - 0x15c1  :  252 - 0xfc
    "11111111", -- 5570 - 0x15c2  :  255 - 0xff
    "11111111", -- 5571 - 0x15c3  :  255 - 0xff
    "11111111", -- 5572 - 0x15c4  :  255 - 0xff
    "11111111", -- 5573 - 0x15c5  :  255 - 0xff
    "00000000", -- 5574 - 0x15c6  :    0 - 0x0
    "00000000", -- 5575 - 0x15c7  :    0 - 0x0
    "11110000", -- 5576 - 0x15c8  :  240 - 0xf0
    "11111100", -- 5577 - 0x15c9  :  252 - 0xfc
    "11111111", -- 5578 - 0x15ca  :  255 - 0xff
    "11111111", -- 5579 - 0x15cb  :  255 - 0xff
    "11111111", -- 5580 - 0x15cc  :  255 - 0xff
    "11111111", -- 5581 - 0x15cd  :  255 - 0xff
    "00000000", -- 5582 - 0x15ce  :    0 - 0x0
    "00000000", -- 5583 - 0x15cf  :    0 - 0x0
    "00000000", -- 5584 - 0x15d0  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 5585 - 0x15d1  :    0 - 0x0
    "00000001", -- 5586 - 0x15d2  :    1 - 0x1
    "00000011", -- 5587 - 0x15d3  :    3 - 0x3
    "00001111", -- 5588 - 0x15d4  :   15 - 0xf
    "00001111", -- 5589 - 0x15d5  :   15 - 0xf
    "00000000", -- 5590 - 0x15d6  :    0 - 0x0
    "00000000", -- 5591 - 0x15d7  :    0 - 0x0
    "00000000", -- 5592 - 0x15d8  :    0 - 0x0
    "00000000", -- 5593 - 0x15d9  :    0 - 0x0
    "00000001", -- 5594 - 0x15da  :    1 - 0x1
    "00000011", -- 5595 - 0x15db  :    3 - 0x3
    "00001111", -- 5596 - 0x15dc  :   15 - 0xf
    "00001111", -- 5597 - 0x15dd  :   15 - 0xf
    "00000000", -- 5598 - 0x15de  :    0 - 0x0
    "00000000", -- 5599 - 0x15df  :    0 - 0x0
    "11111100", -- 5600 - 0x15e0  :  252 - 0xfc -- Background 0x5e
    "11111100", -- 5601 - 0x15e1  :  252 - 0xfc
    "11111100", -- 5602 - 0x15e2  :  252 - 0xfc
    "11111100", -- 5603 - 0x15e3  :  252 - 0xfc
    "11111000", -- 5604 - 0x15e4  :  248 - 0xf8
    "11111100", -- 5605 - 0x15e5  :  252 - 0xfc
    "00111100", -- 5606 - 0x15e6  :   60 - 0x3c
    "00000000", -- 5607 - 0x15e7  :    0 - 0x0
    "11111000", -- 5608 - 0x15e8  :  248 - 0xf8
    "11110000", -- 5609 - 0x15e9  :  240 - 0xf0
    "11100000", -- 5610 - 0x15ea  :  224 - 0xe0
    "11110000", -- 5611 - 0x15eb  :  240 - 0xf0
    "11100000", -- 5612 - 0x15ec  :  224 - 0xe0
    "11000000", -- 5613 - 0x15ed  :  192 - 0xc0
    "00000000", -- 5614 - 0x15ee  :    0 - 0x0
    "00000000", -- 5615 - 0x15ef  :    0 - 0x0
    "00000100", -- 5616 - 0x15f0  :    4 - 0x4 -- Background 0x5f
    "00001100", -- 5617 - 0x15f1  :   12 - 0xc
    "00011100", -- 5618 - 0x15f2  :   28 - 0x1c
    "00001100", -- 5619 - 0x15f3  :   12 - 0xc
    "00011000", -- 5620 - 0x15f4  :   24 - 0x18
    "00111100", -- 5621 - 0x15f5  :   60 - 0x3c
    "00111100", -- 5622 - 0x15f6  :   60 - 0x3c
    "00000000", -- 5623 - 0x15f7  :    0 - 0x0
    "00000000", -- 5624 - 0x15f8  :    0 - 0x0
    "00000000", -- 5625 - 0x15f9  :    0 - 0x0
    "00000000", -- 5626 - 0x15fa  :    0 - 0x0
    "00000000", -- 5627 - 0x15fb  :    0 - 0x0
    "00000000", -- 5628 - 0x15fc  :    0 - 0x0
    "00000000", -- 5629 - 0x15fd  :    0 - 0x0
    "00000000", -- 5630 - 0x15fe  :    0 - 0x0
    "00000000", -- 5631 - 0x15ff  :    0 - 0x0
    "00000000", -- 5632 - 0x1600  :    0 - 0x0 -- Background 0x60
    "00000011", -- 5633 - 0x1601  :    3 - 0x3
    "00001111", -- 5634 - 0x1602  :   15 - 0xf
    "00010011", -- 5635 - 0x1603  :   19 - 0x13
    "00100001", -- 5636 - 0x1604  :   33 - 0x21
    "00100001", -- 5637 - 0x1605  :   33 - 0x21
    "00100001", -- 5638 - 0x1606  :   33 - 0x21
    "01110011", -- 5639 - 0x1607  :  115 - 0x73
    "00000000", -- 5640 - 0x1608  :    0 - 0x0
    "00000011", -- 5641 - 0x1609  :    3 - 0x3
    "00001111", -- 5642 - 0x160a  :   15 - 0xf
    "00011111", -- 5643 - 0x160b  :   31 - 0x1f
    "00111111", -- 5644 - 0x160c  :   63 - 0x3f
    "00111111", -- 5645 - 0x160d  :   63 - 0x3f
    "00111001", -- 5646 - 0x160e  :   57 - 0x39
    "01111011", -- 5647 - 0x160f  :  123 - 0x7b
    "00000000", -- 5648 - 0x1610  :    0 - 0x0 -- Background 0x61
    "11000000", -- 5649 - 0x1611  :  192 - 0xc0
    "11110000", -- 5650 - 0x1612  :  240 - 0xf0
    "11001000", -- 5651 - 0x1613  :  200 - 0xc8
    "10000100", -- 5652 - 0x1614  :  132 - 0x84
    "10000100", -- 5653 - 0x1615  :  132 - 0x84
    "10000100", -- 5654 - 0x1616  :  132 - 0x84
    "11001110", -- 5655 - 0x1617  :  206 - 0xce
    "00000000", -- 5656 - 0x1618  :    0 - 0x0
    "11000000", -- 5657 - 0x1619  :  192 - 0xc0
    "11110000", -- 5658 - 0x161a  :  240 - 0xf0
    "11111000", -- 5659 - 0x161b  :  248 - 0xf8
    "11111100", -- 5660 - 0x161c  :  252 - 0xfc
    "11111100", -- 5661 - 0x161d  :  252 - 0xfc
    "11100100", -- 5662 - 0x161e  :  228 - 0xe4
    "11101110", -- 5663 - 0x161f  :  238 - 0xee
    "10010100", -- 5664 - 0x1620  :  148 - 0x94 -- Background 0x62
    "11101010", -- 5665 - 0x1621  :  234 - 0xea
    "11011110", -- 5666 - 0x1622  :  222 - 0xde
    "11101110", -- 5667 - 0x1623  :  238 - 0xee
    "11011110", -- 5668 - 0x1624  :  222 - 0xde
    "01100110", -- 5669 - 0x1625  :  102 - 0x66
    "01000010", -- 5670 - 0x1626  :   66 - 0x42
    "00000000", -- 5671 - 0x1627  :    0 - 0x0
    "11111110", -- 5672 - 0x1628  :  254 - 0xfe
    "11111110", -- 5673 - 0x1629  :  254 - 0xfe
    "11111110", -- 5674 - 0x162a  :  254 - 0xfe
    "11111110", -- 5675 - 0x162b  :  254 - 0xfe
    "11111110", -- 5676 - 0x162c  :  254 - 0xfe
    "01100110", -- 5677 - 0x162d  :  102 - 0x66
    "01000010", -- 5678 - 0x162e  :   66 - 0x42
    "00000000", -- 5679 - 0x162f  :    0 - 0x0
    "10010100", -- 5680 - 0x1630  :  148 - 0x94 -- Background 0x63
    "11101010", -- 5681 - 0x1631  :  234 - 0xea
    "11011110", -- 5682 - 0x1632  :  222 - 0xde
    "11101110", -- 5683 - 0x1633  :  238 - 0xee
    "11011110", -- 5684 - 0x1634  :  222 - 0xde
    "11001110", -- 5685 - 0x1635  :  206 - 0xce
    "10001100", -- 5686 - 0x1636  :  140 - 0x8c
    "00000000", -- 5687 - 0x1637  :    0 - 0x0
    "11111110", -- 5688 - 0x1638  :  254 - 0xfe
    "11111110", -- 5689 - 0x1639  :  254 - 0xfe
    "11111110", -- 5690 - 0x163a  :  254 - 0xfe
    "11111110", -- 5691 - 0x163b  :  254 - 0xfe
    "11111110", -- 5692 - 0x163c  :  254 - 0xfe
    "11011110", -- 5693 - 0x163d  :  222 - 0xde
    "10001100", -- 5694 - 0x163e  :  140 - 0x8c
    "00000000", -- 5695 - 0x163f  :    0 - 0x0
    "00000000", -- 5696 - 0x1640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 5697 - 0x1641  :    0 - 0x0
    "00000000", -- 5698 - 0x1642  :    0 - 0x0
    "00000000", -- 5699 - 0x1643  :    0 - 0x0
    "00000000", -- 5700 - 0x1644  :    0 - 0x0
    "00000000", -- 5701 - 0x1645  :    0 - 0x0
    "00000000", -- 5702 - 0x1646  :    0 - 0x0
    "00000001", -- 5703 - 0x1647  :    1 - 0x1
    "00000000", -- 5704 - 0x1648  :    0 - 0x0
    "00000000", -- 5705 - 0x1649  :    0 - 0x0
    "00000000", -- 5706 - 0x164a  :    0 - 0x0
    "00000000", -- 5707 - 0x164b  :    0 - 0x0
    "00000000", -- 5708 - 0x164c  :    0 - 0x0
    "00000000", -- 5709 - 0x164d  :    0 - 0x0
    "00000000", -- 5710 - 0x164e  :    0 - 0x0
    "00000000", -- 5711 - 0x164f  :    0 - 0x0
    "00000000", -- 5712 - 0x1650  :    0 - 0x0 -- Background 0x65
    "00000000", -- 5713 - 0x1651  :    0 - 0x0
    "00000000", -- 5714 - 0x1652  :    0 - 0x0
    "00000000", -- 5715 - 0x1653  :    0 - 0x0
    "00000000", -- 5716 - 0x1654  :    0 - 0x0
    "00110110", -- 5717 - 0x1655  :   54 - 0x36
    "00110110", -- 5718 - 0x1656  :   54 - 0x36
    "10010000", -- 5719 - 0x1657  :  144 - 0x90
    "00000000", -- 5720 - 0x1658  :    0 - 0x0
    "00000000", -- 5721 - 0x1659  :    0 - 0x0
    "00000000", -- 5722 - 0x165a  :    0 - 0x0
    "00000000", -- 5723 - 0x165b  :    0 - 0x0
    "01101100", -- 5724 - 0x165c  :  108 - 0x6c
    "11111110", -- 5725 - 0x165d  :  254 - 0xfe
    "11111110", -- 5726 - 0x165e  :  254 - 0xfe
    "11111100", -- 5727 - 0x165f  :  252 - 0xfc
    "00000001", -- 5728 - 0x1660  :    1 - 0x1 -- Background 0x66
    "00000011", -- 5729 - 0x1661  :    3 - 0x3
    "00000111", -- 5730 - 0x1662  :    7 - 0x7
    "00000111", -- 5731 - 0x1663  :    7 - 0x7
    "00011111", -- 5732 - 0x1664  :   31 - 0x1f
    "00011111", -- 5733 - 0x1665  :   31 - 0x1f
    "00011100", -- 5734 - 0x1666  :   28 - 0x1c
    "00000000", -- 5735 - 0x1667  :    0 - 0x0
    "00000000", -- 5736 - 0x1668  :    0 - 0x0
    "00000000", -- 5737 - 0x1669  :    0 - 0x0
    "00000000", -- 5738 - 0x166a  :    0 - 0x0
    "00000000", -- 5739 - 0x166b  :    0 - 0x0
    "00000000", -- 5740 - 0x166c  :    0 - 0x0
    "00000000", -- 5741 - 0x166d  :    0 - 0x0
    "00000000", -- 5742 - 0x166e  :    0 - 0x0
    "00000000", -- 5743 - 0x166f  :    0 - 0x0
    "11111000", -- 5744 - 0x1670  :  248 - 0xf8 -- Background 0x67
    "11111000", -- 5745 - 0x1671  :  248 - 0xf8
    "11111000", -- 5746 - 0x1672  :  248 - 0xf8
    "11111000", -- 5747 - 0x1673  :  248 - 0xf8
    "11111110", -- 5748 - 0x1674  :  254 - 0xfe
    "11111110", -- 5749 - 0x1675  :  254 - 0xfe
    "00001110", -- 5750 - 0x1676  :   14 - 0xe
    "00000000", -- 5751 - 0x1677  :    0 - 0x0
    "00000000", -- 5752 - 0x1678  :    0 - 0x0
    "00000000", -- 5753 - 0x1679  :    0 - 0x0
    "00000000", -- 5754 - 0x167a  :    0 - 0x0
    "00000000", -- 5755 - 0x167b  :    0 - 0x0
    "00000000", -- 5756 - 0x167c  :    0 - 0x0
    "00000000", -- 5757 - 0x167d  :    0 - 0x0
    "00000000", -- 5758 - 0x167e  :    0 - 0x0
    "00000000", -- 5759 - 0x167f  :    0 - 0x0
    "00000111", -- 5760 - 0x1680  :    7 - 0x7 -- Background 0x68
    "00001111", -- 5761 - 0x1681  :   15 - 0xf
    "00011111", -- 5762 - 0x1682  :   31 - 0x1f
    "00011111", -- 5763 - 0x1683  :   31 - 0x1f
    "00111111", -- 5764 - 0x1684  :   63 - 0x3f
    "00111111", -- 5765 - 0x1685  :   63 - 0x3f
    "00111000", -- 5766 - 0x1686  :   56 - 0x38
    "00000000", -- 5767 - 0x1687  :    0 - 0x0
    "00000000", -- 5768 - 0x1688  :    0 - 0x0
    "00000000", -- 5769 - 0x1689  :    0 - 0x0
    "00000000", -- 5770 - 0x168a  :    0 - 0x0
    "00000000", -- 5771 - 0x168b  :    0 - 0x0
    "00000000", -- 5772 - 0x168c  :    0 - 0x0
    "00000000", -- 5773 - 0x168d  :    0 - 0x0
    "00000000", -- 5774 - 0x168e  :    0 - 0x0
    "00000000", -- 5775 - 0x168f  :    0 - 0x0
    "11111000", -- 5776 - 0x1690  :  248 - 0xf8 -- Background 0x69
    "11110000", -- 5777 - 0x1691  :  240 - 0xf0
    "11110000", -- 5778 - 0x1692  :  240 - 0xf0
    "11100000", -- 5779 - 0x1693  :  224 - 0xe0
    "11111000", -- 5780 - 0x1694  :  248 - 0xf8
    "11111000", -- 5781 - 0x1695  :  248 - 0xf8
    "00111000", -- 5782 - 0x1696  :   56 - 0x38
    "00000000", -- 5783 - 0x1697  :    0 - 0x0
    "00000000", -- 5784 - 0x1698  :    0 - 0x0
    "00000000", -- 5785 - 0x1699  :    0 - 0x0
    "00000000", -- 5786 - 0x169a  :    0 - 0x0
    "00000000", -- 5787 - 0x169b  :    0 - 0x0
    "00000000", -- 5788 - 0x169c  :    0 - 0x0
    "00000000", -- 5789 - 0x169d  :    0 - 0x0
    "00000000", -- 5790 - 0x169e  :    0 - 0x0
    "00000000", -- 5791 - 0x169f  :    0 - 0x0
    "00000000", -- 5792 - 0x16a0  :    0 - 0x0 -- Background 0x6a
    "00011111", -- 5793 - 0x16a1  :   31 - 0x1f
    "01111111", -- 5794 - 0x16a2  :  127 - 0x7f
    "00111111", -- 5795 - 0x16a3  :   63 - 0x3f
    "00001111", -- 5796 - 0x16a4  :   15 - 0xf
    "00000111", -- 5797 - 0x16a5  :    7 - 0x7
    "00000000", -- 5798 - 0x16a6  :    0 - 0x0
    "00000000", -- 5799 - 0x16a7  :    0 - 0x0
    "00000000", -- 5800 - 0x16a8  :    0 - 0x0
    "00011111", -- 5801 - 0x16a9  :   31 - 0x1f
    "01111111", -- 5802 - 0x16aa  :  127 - 0x7f
    "00111111", -- 5803 - 0x16ab  :   63 - 0x3f
    "00001111", -- 5804 - 0x16ac  :   15 - 0xf
    "00000111", -- 5805 - 0x16ad  :    7 - 0x7
    "00000000", -- 5806 - 0x16ae  :    0 - 0x0
    "00000000", -- 5807 - 0x16af  :    0 - 0x0
    "00000000", -- 5808 - 0x16b0  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 5809 - 0x16b1  :    0 - 0x0
    "11000000", -- 5810 - 0x16b2  :  192 - 0xc0
    "11110000", -- 5811 - 0x16b3  :  240 - 0xf0
    "11111000", -- 5812 - 0x16b4  :  248 - 0xf8
    "11111000", -- 5813 - 0x16b5  :  248 - 0xf8
    "11100000", -- 5814 - 0x16b6  :  224 - 0xe0
    "00000000", -- 5815 - 0x16b7  :    0 - 0x0
    "00000000", -- 5816 - 0x16b8  :    0 - 0x0
    "00000000", -- 5817 - 0x16b9  :    0 - 0x0
    "11000000", -- 5818 - 0x16ba  :  192 - 0xc0
    "11110000", -- 5819 - 0x16bb  :  240 - 0xf0
    "11111000", -- 5820 - 0x16bc  :  248 - 0xf8
    "11111000", -- 5821 - 0x16bd  :  248 - 0xf8
    "11100000", -- 5822 - 0x16be  :  224 - 0xe0
    "00000000", -- 5823 - 0x16bf  :    0 - 0x0
    "00000000", -- 5824 - 0x16c0  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 5825 - 0x16c1  :    0 - 0x0
    "00000000", -- 5826 - 0x16c2  :    0 - 0x0
    "00000000", -- 5827 - 0x16c3  :    0 - 0x0
    "00000000", -- 5828 - 0x16c4  :    0 - 0x0
    "00000000", -- 5829 - 0x16c5  :    0 - 0x0
    "00000000", -- 5830 - 0x16c6  :    0 - 0x0
    "00000000", -- 5831 - 0x16c7  :    0 - 0x0
    "00000000", -- 5832 - 0x16c8  :    0 - 0x0
    "00000000", -- 5833 - 0x16c9  :    0 - 0x0
    "00000000", -- 5834 - 0x16ca  :    0 - 0x0
    "00000000", -- 5835 - 0x16cb  :    0 - 0x0
    "00000000", -- 5836 - 0x16cc  :    0 - 0x0
    "00000000", -- 5837 - 0x16cd  :    0 - 0x0
    "00000000", -- 5838 - 0x16ce  :    0 - 0x0
    "00000000", -- 5839 - 0x16cf  :    0 - 0x0
    "00000000", -- 5840 - 0x16d0  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 5841 - 0x16d1  :    0 - 0x0
    "00000000", -- 5842 - 0x16d2  :    0 - 0x0
    "00000000", -- 5843 - 0x16d3  :    0 - 0x0
    "00000000", -- 5844 - 0x16d4  :    0 - 0x0
    "00000000", -- 5845 - 0x16d5  :    0 - 0x0
    "00000000", -- 5846 - 0x16d6  :    0 - 0x0
    "00000000", -- 5847 - 0x16d7  :    0 - 0x0
    "00000000", -- 5848 - 0x16d8  :    0 - 0x0
    "00000000", -- 5849 - 0x16d9  :    0 - 0x0
    "00000000", -- 5850 - 0x16da  :    0 - 0x0
    "00000000", -- 5851 - 0x16db  :    0 - 0x0
    "00000000", -- 5852 - 0x16dc  :    0 - 0x0
    "00000000", -- 5853 - 0x16dd  :    0 - 0x0
    "00000000", -- 5854 - 0x16de  :    0 - 0x0
    "00000000", -- 5855 - 0x16df  :    0 - 0x0
    "00000000", -- 5856 - 0x16e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 5857 - 0x16e1  :    0 - 0x0
    "00000000", -- 5858 - 0x16e2  :    0 - 0x0
    "00000000", -- 5859 - 0x16e3  :    0 - 0x0
    "00000000", -- 5860 - 0x16e4  :    0 - 0x0
    "00000000", -- 5861 - 0x16e5  :    0 - 0x0
    "00000000", -- 5862 - 0x16e6  :    0 - 0x0
    "00000000", -- 5863 - 0x16e7  :    0 - 0x0
    "00000000", -- 5864 - 0x16e8  :    0 - 0x0
    "00000000", -- 5865 - 0x16e9  :    0 - 0x0
    "00000000", -- 5866 - 0x16ea  :    0 - 0x0
    "00000000", -- 5867 - 0x16eb  :    0 - 0x0
    "00000000", -- 5868 - 0x16ec  :    0 - 0x0
    "00000000", -- 5869 - 0x16ed  :    0 - 0x0
    "00000000", -- 5870 - 0x16ee  :    0 - 0x0
    "00000000", -- 5871 - 0x16ef  :    0 - 0x0
    "00000000", -- 5872 - 0x16f0  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 5873 - 0x16f1  :    0 - 0x0
    "00000000", -- 5874 - 0x16f2  :    0 - 0x0
    "00000000", -- 5875 - 0x16f3  :    0 - 0x0
    "00000000", -- 5876 - 0x16f4  :    0 - 0x0
    "00000000", -- 5877 - 0x16f5  :    0 - 0x0
    "00000000", -- 5878 - 0x16f6  :    0 - 0x0
    "00000000", -- 5879 - 0x16f7  :    0 - 0x0
    "00000000", -- 5880 - 0x16f8  :    0 - 0x0
    "00000000", -- 5881 - 0x16f9  :    0 - 0x0
    "00000000", -- 5882 - 0x16fa  :    0 - 0x0
    "00000000", -- 5883 - 0x16fb  :    0 - 0x0
    "00000000", -- 5884 - 0x16fc  :    0 - 0x0
    "00000000", -- 5885 - 0x16fd  :    0 - 0x0
    "00000000", -- 5886 - 0x16fe  :    0 - 0x0
    "00000000", -- 5887 - 0x16ff  :    0 - 0x0
    "11111111", -- 5888 - 0x1700  :  255 - 0xff -- Background 0x70
    "11111111", -- 5889 - 0x1701  :  255 - 0xff
    "11111111", -- 5890 - 0x1702  :  255 - 0xff
    "11111111", -- 5891 - 0x1703  :  255 - 0xff
    "11111111", -- 5892 - 0x1704  :  255 - 0xff
    "11111111", -- 5893 - 0x1705  :  255 - 0xff
    "11111111", -- 5894 - 0x1706  :  255 - 0xff
    "11111111", -- 5895 - 0x1707  :  255 - 0xff
    "11111111", -- 5896 - 0x1708  :  255 - 0xff
    "11111111", -- 5897 - 0x1709  :  255 - 0xff
    "11111111", -- 5898 - 0x170a  :  255 - 0xff
    "11111111", -- 5899 - 0x170b  :  255 - 0xff
    "11111111", -- 5900 - 0x170c  :  255 - 0xff
    "11111111", -- 5901 - 0x170d  :  255 - 0xff
    "11111111", -- 5902 - 0x170e  :  255 - 0xff
    "11111111", -- 5903 - 0x170f  :  255 - 0xff
    "11111111", -- 5904 - 0x1710  :  255 - 0xff -- Background 0x71
    "11111111", -- 5905 - 0x1711  :  255 - 0xff
    "11111111", -- 5906 - 0x1712  :  255 - 0xff
    "11111111", -- 5907 - 0x1713  :  255 - 0xff
    "11111111", -- 5908 - 0x1714  :  255 - 0xff
    "11111111", -- 5909 - 0x1715  :  255 - 0xff
    "11111111", -- 5910 - 0x1716  :  255 - 0xff
    "11111111", -- 5911 - 0x1717  :  255 - 0xff
    "11111111", -- 5912 - 0x1718  :  255 - 0xff
    "11111111", -- 5913 - 0x1719  :  255 - 0xff
    "11111111", -- 5914 - 0x171a  :  255 - 0xff
    "11111111", -- 5915 - 0x171b  :  255 - 0xff
    "11111111", -- 5916 - 0x171c  :  255 - 0xff
    "11111111", -- 5917 - 0x171d  :  255 - 0xff
    "11111111", -- 5918 - 0x171e  :  255 - 0xff
    "11111111", -- 5919 - 0x171f  :  255 - 0xff
    "11111111", -- 5920 - 0x1720  :  255 - 0xff -- Background 0x72
    "11111111", -- 5921 - 0x1721  :  255 - 0xff
    "11111111", -- 5922 - 0x1722  :  255 - 0xff
    "11111111", -- 5923 - 0x1723  :  255 - 0xff
    "11111111", -- 5924 - 0x1724  :  255 - 0xff
    "11111111", -- 5925 - 0x1725  :  255 - 0xff
    "11111111", -- 5926 - 0x1726  :  255 - 0xff
    "11111111", -- 5927 - 0x1727  :  255 - 0xff
    "11111111", -- 5928 - 0x1728  :  255 - 0xff
    "11111111", -- 5929 - 0x1729  :  255 - 0xff
    "11111111", -- 5930 - 0x172a  :  255 - 0xff
    "11111111", -- 5931 - 0x172b  :  255 - 0xff
    "11111111", -- 5932 - 0x172c  :  255 - 0xff
    "11111111", -- 5933 - 0x172d  :  255 - 0xff
    "11111111", -- 5934 - 0x172e  :  255 - 0xff
    "11111111", -- 5935 - 0x172f  :  255 - 0xff
    "11111111", -- 5936 - 0x1730  :  255 - 0xff -- Background 0x73
    "11111111", -- 5937 - 0x1731  :  255 - 0xff
    "11111111", -- 5938 - 0x1732  :  255 - 0xff
    "11111111", -- 5939 - 0x1733  :  255 - 0xff
    "11111111", -- 5940 - 0x1734  :  255 - 0xff
    "11111111", -- 5941 - 0x1735  :  255 - 0xff
    "11111111", -- 5942 - 0x1736  :  255 - 0xff
    "11111111", -- 5943 - 0x1737  :  255 - 0xff
    "11111111", -- 5944 - 0x1738  :  255 - 0xff
    "11111111", -- 5945 - 0x1739  :  255 - 0xff
    "11111111", -- 5946 - 0x173a  :  255 - 0xff
    "11111111", -- 5947 - 0x173b  :  255 - 0xff
    "11111111", -- 5948 - 0x173c  :  255 - 0xff
    "11111111", -- 5949 - 0x173d  :  255 - 0xff
    "11111111", -- 5950 - 0x173e  :  255 - 0xff
    "11111111", -- 5951 - 0x173f  :  255 - 0xff
    "11111111", -- 5952 - 0x1740  :  255 - 0xff -- Background 0x74
    "11111111", -- 5953 - 0x1741  :  255 - 0xff
    "11111111", -- 5954 - 0x1742  :  255 - 0xff
    "11111111", -- 5955 - 0x1743  :  255 - 0xff
    "11111111", -- 5956 - 0x1744  :  255 - 0xff
    "11111111", -- 5957 - 0x1745  :  255 - 0xff
    "11111111", -- 5958 - 0x1746  :  255 - 0xff
    "11111111", -- 5959 - 0x1747  :  255 - 0xff
    "11111111", -- 5960 - 0x1748  :  255 - 0xff
    "11111111", -- 5961 - 0x1749  :  255 - 0xff
    "11111111", -- 5962 - 0x174a  :  255 - 0xff
    "11111111", -- 5963 - 0x174b  :  255 - 0xff
    "11111111", -- 5964 - 0x174c  :  255 - 0xff
    "11111111", -- 5965 - 0x174d  :  255 - 0xff
    "11111111", -- 5966 - 0x174e  :  255 - 0xff
    "11111111", -- 5967 - 0x174f  :  255 - 0xff
    "11111111", -- 5968 - 0x1750  :  255 - 0xff -- Background 0x75
    "11111111", -- 5969 - 0x1751  :  255 - 0xff
    "11111111", -- 5970 - 0x1752  :  255 - 0xff
    "11111111", -- 5971 - 0x1753  :  255 - 0xff
    "11111111", -- 5972 - 0x1754  :  255 - 0xff
    "11111111", -- 5973 - 0x1755  :  255 - 0xff
    "11111111", -- 5974 - 0x1756  :  255 - 0xff
    "11111111", -- 5975 - 0x1757  :  255 - 0xff
    "11111111", -- 5976 - 0x1758  :  255 - 0xff
    "11111111", -- 5977 - 0x1759  :  255 - 0xff
    "11111111", -- 5978 - 0x175a  :  255 - 0xff
    "11111111", -- 5979 - 0x175b  :  255 - 0xff
    "11111111", -- 5980 - 0x175c  :  255 - 0xff
    "11111111", -- 5981 - 0x175d  :  255 - 0xff
    "11111111", -- 5982 - 0x175e  :  255 - 0xff
    "11111111", -- 5983 - 0x175f  :  255 - 0xff
    "11111111", -- 5984 - 0x1760  :  255 - 0xff -- Background 0x76
    "11111111", -- 5985 - 0x1761  :  255 - 0xff
    "11111111", -- 5986 - 0x1762  :  255 - 0xff
    "11111111", -- 5987 - 0x1763  :  255 - 0xff
    "11111111", -- 5988 - 0x1764  :  255 - 0xff
    "11111111", -- 5989 - 0x1765  :  255 - 0xff
    "11111111", -- 5990 - 0x1766  :  255 - 0xff
    "11111111", -- 5991 - 0x1767  :  255 - 0xff
    "11111111", -- 5992 - 0x1768  :  255 - 0xff
    "11111111", -- 5993 - 0x1769  :  255 - 0xff
    "11111111", -- 5994 - 0x176a  :  255 - 0xff
    "11111111", -- 5995 - 0x176b  :  255 - 0xff
    "11111111", -- 5996 - 0x176c  :  255 - 0xff
    "11111111", -- 5997 - 0x176d  :  255 - 0xff
    "11111111", -- 5998 - 0x176e  :  255 - 0xff
    "11111111", -- 5999 - 0x176f  :  255 - 0xff
    "11111111", -- 6000 - 0x1770  :  255 - 0xff -- Background 0x77
    "11111111", -- 6001 - 0x1771  :  255 - 0xff
    "11111111", -- 6002 - 0x1772  :  255 - 0xff
    "11111111", -- 6003 - 0x1773  :  255 - 0xff
    "11111111", -- 6004 - 0x1774  :  255 - 0xff
    "11111111", -- 6005 - 0x1775  :  255 - 0xff
    "11111111", -- 6006 - 0x1776  :  255 - 0xff
    "11111111", -- 6007 - 0x1777  :  255 - 0xff
    "11111111", -- 6008 - 0x1778  :  255 - 0xff
    "11111111", -- 6009 - 0x1779  :  255 - 0xff
    "11111111", -- 6010 - 0x177a  :  255 - 0xff
    "11111111", -- 6011 - 0x177b  :  255 - 0xff
    "11111111", -- 6012 - 0x177c  :  255 - 0xff
    "11111111", -- 6013 - 0x177d  :  255 - 0xff
    "11111111", -- 6014 - 0x177e  :  255 - 0xff
    "11111111", -- 6015 - 0x177f  :  255 - 0xff
    "11111111", -- 6016 - 0x1780  :  255 - 0xff -- Background 0x78
    "11111111", -- 6017 - 0x1781  :  255 - 0xff
    "11111111", -- 6018 - 0x1782  :  255 - 0xff
    "11111111", -- 6019 - 0x1783  :  255 - 0xff
    "11111111", -- 6020 - 0x1784  :  255 - 0xff
    "11111111", -- 6021 - 0x1785  :  255 - 0xff
    "11111111", -- 6022 - 0x1786  :  255 - 0xff
    "11111111", -- 6023 - 0x1787  :  255 - 0xff
    "11111111", -- 6024 - 0x1788  :  255 - 0xff
    "11111111", -- 6025 - 0x1789  :  255 - 0xff
    "11111111", -- 6026 - 0x178a  :  255 - 0xff
    "11111111", -- 6027 - 0x178b  :  255 - 0xff
    "11111111", -- 6028 - 0x178c  :  255 - 0xff
    "11111111", -- 6029 - 0x178d  :  255 - 0xff
    "11111111", -- 6030 - 0x178e  :  255 - 0xff
    "11111111", -- 6031 - 0x178f  :  255 - 0xff
    "11111111", -- 6032 - 0x1790  :  255 - 0xff -- Background 0x79
    "11111111", -- 6033 - 0x1791  :  255 - 0xff
    "11111111", -- 6034 - 0x1792  :  255 - 0xff
    "11111111", -- 6035 - 0x1793  :  255 - 0xff
    "11111111", -- 6036 - 0x1794  :  255 - 0xff
    "11111111", -- 6037 - 0x1795  :  255 - 0xff
    "11111111", -- 6038 - 0x1796  :  255 - 0xff
    "11111111", -- 6039 - 0x1797  :  255 - 0xff
    "11111111", -- 6040 - 0x1798  :  255 - 0xff
    "11111111", -- 6041 - 0x1799  :  255 - 0xff
    "11111111", -- 6042 - 0x179a  :  255 - 0xff
    "11111111", -- 6043 - 0x179b  :  255 - 0xff
    "11111111", -- 6044 - 0x179c  :  255 - 0xff
    "11111111", -- 6045 - 0x179d  :  255 - 0xff
    "11111111", -- 6046 - 0x179e  :  255 - 0xff
    "11111111", -- 6047 - 0x179f  :  255 - 0xff
    "11111111", -- 6048 - 0x17a0  :  255 - 0xff -- Background 0x7a
    "11111111", -- 6049 - 0x17a1  :  255 - 0xff
    "11111111", -- 6050 - 0x17a2  :  255 - 0xff
    "11111111", -- 6051 - 0x17a3  :  255 - 0xff
    "11111111", -- 6052 - 0x17a4  :  255 - 0xff
    "11111111", -- 6053 - 0x17a5  :  255 - 0xff
    "11111111", -- 6054 - 0x17a6  :  255 - 0xff
    "11111111", -- 6055 - 0x17a7  :  255 - 0xff
    "11111111", -- 6056 - 0x17a8  :  255 - 0xff
    "11111111", -- 6057 - 0x17a9  :  255 - 0xff
    "11111111", -- 6058 - 0x17aa  :  255 - 0xff
    "11111111", -- 6059 - 0x17ab  :  255 - 0xff
    "11111111", -- 6060 - 0x17ac  :  255 - 0xff
    "11111111", -- 6061 - 0x17ad  :  255 - 0xff
    "11111111", -- 6062 - 0x17ae  :  255 - 0xff
    "11111111", -- 6063 - 0x17af  :  255 - 0xff
    "11111111", -- 6064 - 0x17b0  :  255 - 0xff -- Background 0x7b
    "11111111", -- 6065 - 0x17b1  :  255 - 0xff
    "11111111", -- 6066 - 0x17b2  :  255 - 0xff
    "11111111", -- 6067 - 0x17b3  :  255 - 0xff
    "11111111", -- 6068 - 0x17b4  :  255 - 0xff
    "11111111", -- 6069 - 0x17b5  :  255 - 0xff
    "11111111", -- 6070 - 0x17b6  :  255 - 0xff
    "11111111", -- 6071 - 0x17b7  :  255 - 0xff
    "11111111", -- 6072 - 0x17b8  :  255 - 0xff
    "11111111", -- 6073 - 0x17b9  :  255 - 0xff
    "11111111", -- 6074 - 0x17ba  :  255 - 0xff
    "11111111", -- 6075 - 0x17bb  :  255 - 0xff
    "11111111", -- 6076 - 0x17bc  :  255 - 0xff
    "11111111", -- 6077 - 0x17bd  :  255 - 0xff
    "11111111", -- 6078 - 0x17be  :  255 - 0xff
    "11111111", -- 6079 - 0x17bf  :  255 - 0xff
    "11111111", -- 6080 - 0x17c0  :  255 - 0xff -- Background 0x7c
    "11111111", -- 6081 - 0x17c1  :  255 - 0xff
    "11111111", -- 6082 - 0x17c2  :  255 - 0xff
    "11111111", -- 6083 - 0x17c3  :  255 - 0xff
    "11111111", -- 6084 - 0x17c4  :  255 - 0xff
    "11111111", -- 6085 - 0x17c5  :  255 - 0xff
    "11111111", -- 6086 - 0x17c6  :  255 - 0xff
    "11111111", -- 6087 - 0x17c7  :  255 - 0xff
    "11111111", -- 6088 - 0x17c8  :  255 - 0xff
    "11111111", -- 6089 - 0x17c9  :  255 - 0xff
    "11111111", -- 6090 - 0x17ca  :  255 - 0xff
    "11111111", -- 6091 - 0x17cb  :  255 - 0xff
    "11111111", -- 6092 - 0x17cc  :  255 - 0xff
    "11111111", -- 6093 - 0x17cd  :  255 - 0xff
    "11111111", -- 6094 - 0x17ce  :  255 - 0xff
    "11111111", -- 6095 - 0x17cf  :  255 - 0xff
    "11111111", -- 6096 - 0x17d0  :  255 - 0xff -- Background 0x7d
    "11111111", -- 6097 - 0x17d1  :  255 - 0xff
    "11111111", -- 6098 - 0x17d2  :  255 - 0xff
    "11111111", -- 6099 - 0x17d3  :  255 - 0xff
    "11111111", -- 6100 - 0x17d4  :  255 - 0xff
    "11111111", -- 6101 - 0x17d5  :  255 - 0xff
    "11111111", -- 6102 - 0x17d6  :  255 - 0xff
    "11111111", -- 6103 - 0x17d7  :  255 - 0xff
    "11111111", -- 6104 - 0x17d8  :  255 - 0xff
    "11111111", -- 6105 - 0x17d9  :  255 - 0xff
    "11111111", -- 6106 - 0x17da  :  255 - 0xff
    "11111111", -- 6107 - 0x17db  :  255 - 0xff
    "11111111", -- 6108 - 0x17dc  :  255 - 0xff
    "11111111", -- 6109 - 0x17dd  :  255 - 0xff
    "11111111", -- 6110 - 0x17de  :  255 - 0xff
    "11111111", -- 6111 - 0x17df  :  255 - 0xff
    "11111111", -- 6112 - 0x17e0  :  255 - 0xff -- Background 0x7e
    "11111111", -- 6113 - 0x17e1  :  255 - 0xff
    "11111111", -- 6114 - 0x17e2  :  255 - 0xff
    "11111111", -- 6115 - 0x17e3  :  255 - 0xff
    "11111111", -- 6116 - 0x17e4  :  255 - 0xff
    "11111111", -- 6117 - 0x17e5  :  255 - 0xff
    "11111111", -- 6118 - 0x17e6  :  255 - 0xff
    "11111111", -- 6119 - 0x17e7  :  255 - 0xff
    "11111111", -- 6120 - 0x17e8  :  255 - 0xff
    "11111111", -- 6121 - 0x17e9  :  255 - 0xff
    "11111111", -- 6122 - 0x17ea  :  255 - 0xff
    "11111111", -- 6123 - 0x17eb  :  255 - 0xff
    "11111111", -- 6124 - 0x17ec  :  255 - 0xff
    "11111111", -- 6125 - 0x17ed  :  255 - 0xff
    "11111111", -- 6126 - 0x17ee  :  255 - 0xff
    "11111111", -- 6127 - 0x17ef  :  255 - 0xff
    "11111111", -- 6128 - 0x17f0  :  255 - 0xff -- Background 0x7f
    "11111111", -- 6129 - 0x17f1  :  255 - 0xff
    "11111111", -- 6130 - 0x17f2  :  255 - 0xff
    "11111111", -- 6131 - 0x17f3  :  255 - 0xff
    "11111111", -- 6132 - 0x17f4  :  255 - 0xff
    "11111111", -- 6133 - 0x17f5  :  255 - 0xff
    "11111111", -- 6134 - 0x17f6  :  255 - 0xff
    "11111111", -- 6135 - 0x17f7  :  255 - 0xff
    "11111111", -- 6136 - 0x17f8  :  255 - 0xff
    "11111111", -- 6137 - 0x17f9  :  255 - 0xff
    "11111111", -- 6138 - 0x17fa  :  255 - 0xff
    "11111111", -- 6139 - 0x17fb  :  255 - 0xff
    "11111111", -- 6140 - 0x17fc  :  255 - 0xff
    "11111111", -- 6141 - 0x17fd  :  255 - 0xff
    "11111111", -- 6142 - 0x17fe  :  255 - 0xff
    "11111111", -- 6143 - 0x17ff  :  255 - 0xff
    "11111111", -- 6144 - 0x1800  :  255 - 0xff -- Background 0x80
    "11111111", -- 6145 - 0x1801  :  255 - 0xff
    "11111111", -- 6146 - 0x1802  :  255 - 0xff
    "11111111", -- 6147 - 0x1803  :  255 - 0xff
    "11111111", -- 6148 - 0x1804  :  255 - 0xff
    "11111111", -- 6149 - 0x1805  :  255 - 0xff
    "11111111", -- 6150 - 0x1806  :  255 - 0xff
    "11111111", -- 6151 - 0x1807  :  255 - 0xff
    "11111111", -- 6152 - 0x1808  :  255 - 0xff
    "11111111", -- 6153 - 0x1809  :  255 - 0xff
    "11111111", -- 6154 - 0x180a  :  255 - 0xff
    "11111111", -- 6155 - 0x180b  :  255 - 0xff
    "11111111", -- 6156 - 0x180c  :  255 - 0xff
    "11111111", -- 6157 - 0x180d  :  255 - 0xff
    "11111111", -- 6158 - 0x180e  :  255 - 0xff
    "11111111", -- 6159 - 0x180f  :  255 - 0xff
    "11111111", -- 6160 - 0x1810  :  255 - 0xff -- Background 0x81
    "11111111", -- 6161 - 0x1811  :  255 - 0xff
    "11111111", -- 6162 - 0x1812  :  255 - 0xff
    "11111111", -- 6163 - 0x1813  :  255 - 0xff
    "11111111", -- 6164 - 0x1814  :  255 - 0xff
    "11111111", -- 6165 - 0x1815  :  255 - 0xff
    "11111111", -- 6166 - 0x1816  :  255 - 0xff
    "11111111", -- 6167 - 0x1817  :  255 - 0xff
    "11111111", -- 6168 - 0x1818  :  255 - 0xff
    "11111111", -- 6169 - 0x1819  :  255 - 0xff
    "11111111", -- 6170 - 0x181a  :  255 - 0xff
    "11111111", -- 6171 - 0x181b  :  255 - 0xff
    "11111111", -- 6172 - 0x181c  :  255 - 0xff
    "11111111", -- 6173 - 0x181d  :  255 - 0xff
    "11111111", -- 6174 - 0x181e  :  255 - 0xff
    "11111111", -- 6175 - 0x181f  :  255 - 0xff
    "11111111", -- 6176 - 0x1820  :  255 - 0xff -- Background 0x82
    "11111111", -- 6177 - 0x1821  :  255 - 0xff
    "11111111", -- 6178 - 0x1822  :  255 - 0xff
    "11111111", -- 6179 - 0x1823  :  255 - 0xff
    "11111111", -- 6180 - 0x1824  :  255 - 0xff
    "11111111", -- 6181 - 0x1825  :  255 - 0xff
    "11111111", -- 6182 - 0x1826  :  255 - 0xff
    "11111111", -- 6183 - 0x1827  :  255 - 0xff
    "11111111", -- 6184 - 0x1828  :  255 - 0xff
    "11111111", -- 6185 - 0x1829  :  255 - 0xff
    "11111111", -- 6186 - 0x182a  :  255 - 0xff
    "11111111", -- 6187 - 0x182b  :  255 - 0xff
    "11111111", -- 6188 - 0x182c  :  255 - 0xff
    "11111111", -- 6189 - 0x182d  :  255 - 0xff
    "11111111", -- 6190 - 0x182e  :  255 - 0xff
    "11111111", -- 6191 - 0x182f  :  255 - 0xff
    "11111111", -- 6192 - 0x1830  :  255 - 0xff -- Background 0x83
    "11111111", -- 6193 - 0x1831  :  255 - 0xff
    "11111111", -- 6194 - 0x1832  :  255 - 0xff
    "11111111", -- 6195 - 0x1833  :  255 - 0xff
    "11111111", -- 6196 - 0x1834  :  255 - 0xff
    "11111111", -- 6197 - 0x1835  :  255 - 0xff
    "11111111", -- 6198 - 0x1836  :  255 - 0xff
    "11111111", -- 6199 - 0x1837  :  255 - 0xff
    "11111111", -- 6200 - 0x1838  :  255 - 0xff
    "11111111", -- 6201 - 0x1839  :  255 - 0xff
    "11111111", -- 6202 - 0x183a  :  255 - 0xff
    "11111111", -- 6203 - 0x183b  :  255 - 0xff
    "11111111", -- 6204 - 0x183c  :  255 - 0xff
    "11111111", -- 6205 - 0x183d  :  255 - 0xff
    "11111111", -- 6206 - 0x183e  :  255 - 0xff
    "11111111", -- 6207 - 0x183f  :  255 - 0xff
    "11111111", -- 6208 - 0x1840  :  255 - 0xff -- Background 0x84
    "11111111", -- 6209 - 0x1841  :  255 - 0xff
    "11111111", -- 6210 - 0x1842  :  255 - 0xff
    "11111111", -- 6211 - 0x1843  :  255 - 0xff
    "11111111", -- 6212 - 0x1844  :  255 - 0xff
    "11111111", -- 6213 - 0x1845  :  255 - 0xff
    "11111111", -- 6214 - 0x1846  :  255 - 0xff
    "11111111", -- 6215 - 0x1847  :  255 - 0xff
    "11111111", -- 6216 - 0x1848  :  255 - 0xff
    "11111111", -- 6217 - 0x1849  :  255 - 0xff
    "11111111", -- 6218 - 0x184a  :  255 - 0xff
    "11111111", -- 6219 - 0x184b  :  255 - 0xff
    "11111111", -- 6220 - 0x184c  :  255 - 0xff
    "11111111", -- 6221 - 0x184d  :  255 - 0xff
    "11111111", -- 6222 - 0x184e  :  255 - 0xff
    "11111111", -- 6223 - 0x184f  :  255 - 0xff
    "11111111", -- 6224 - 0x1850  :  255 - 0xff -- Background 0x85
    "11111111", -- 6225 - 0x1851  :  255 - 0xff
    "11111111", -- 6226 - 0x1852  :  255 - 0xff
    "11111111", -- 6227 - 0x1853  :  255 - 0xff
    "11111111", -- 6228 - 0x1854  :  255 - 0xff
    "11111111", -- 6229 - 0x1855  :  255 - 0xff
    "11111111", -- 6230 - 0x1856  :  255 - 0xff
    "11111111", -- 6231 - 0x1857  :  255 - 0xff
    "11111111", -- 6232 - 0x1858  :  255 - 0xff
    "11111111", -- 6233 - 0x1859  :  255 - 0xff
    "11111111", -- 6234 - 0x185a  :  255 - 0xff
    "11111111", -- 6235 - 0x185b  :  255 - 0xff
    "11111111", -- 6236 - 0x185c  :  255 - 0xff
    "11111111", -- 6237 - 0x185d  :  255 - 0xff
    "11111111", -- 6238 - 0x185e  :  255 - 0xff
    "11111111", -- 6239 - 0x185f  :  255 - 0xff
    "11111111", -- 6240 - 0x1860  :  255 - 0xff -- Background 0x86
    "11111111", -- 6241 - 0x1861  :  255 - 0xff
    "11111111", -- 6242 - 0x1862  :  255 - 0xff
    "11111111", -- 6243 - 0x1863  :  255 - 0xff
    "11111111", -- 6244 - 0x1864  :  255 - 0xff
    "11111111", -- 6245 - 0x1865  :  255 - 0xff
    "11111111", -- 6246 - 0x1866  :  255 - 0xff
    "11111111", -- 6247 - 0x1867  :  255 - 0xff
    "11111111", -- 6248 - 0x1868  :  255 - 0xff
    "11111111", -- 6249 - 0x1869  :  255 - 0xff
    "11111111", -- 6250 - 0x186a  :  255 - 0xff
    "11111111", -- 6251 - 0x186b  :  255 - 0xff
    "11111111", -- 6252 - 0x186c  :  255 - 0xff
    "11111111", -- 6253 - 0x186d  :  255 - 0xff
    "11111111", -- 6254 - 0x186e  :  255 - 0xff
    "11111111", -- 6255 - 0x186f  :  255 - 0xff
    "11111111", -- 6256 - 0x1870  :  255 - 0xff -- Background 0x87
    "11111111", -- 6257 - 0x1871  :  255 - 0xff
    "11111111", -- 6258 - 0x1872  :  255 - 0xff
    "11111111", -- 6259 - 0x1873  :  255 - 0xff
    "11111111", -- 6260 - 0x1874  :  255 - 0xff
    "11111111", -- 6261 - 0x1875  :  255 - 0xff
    "11111111", -- 6262 - 0x1876  :  255 - 0xff
    "11111111", -- 6263 - 0x1877  :  255 - 0xff
    "11111111", -- 6264 - 0x1878  :  255 - 0xff
    "11111111", -- 6265 - 0x1879  :  255 - 0xff
    "11111111", -- 6266 - 0x187a  :  255 - 0xff
    "11111111", -- 6267 - 0x187b  :  255 - 0xff
    "11111111", -- 6268 - 0x187c  :  255 - 0xff
    "11111111", -- 6269 - 0x187d  :  255 - 0xff
    "11111111", -- 6270 - 0x187e  :  255 - 0xff
    "11111111", -- 6271 - 0x187f  :  255 - 0xff
    "11111111", -- 6272 - 0x1880  :  255 - 0xff -- Background 0x88
    "11111111", -- 6273 - 0x1881  :  255 - 0xff
    "11111111", -- 6274 - 0x1882  :  255 - 0xff
    "11111111", -- 6275 - 0x1883  :  255 - 0xff
    "11111111", -- 6276 - 0x1884  :  255 - 0xff
    "11111111", -- 6277 - 0x1885  :  255 - 0xff
    "11111111", -- 6278 - 0x1886  :  255 - 0xff
    "11111111", -- 6279 - 0x1887  :  255 - 0xff
    "11111111", -- 6280 - 0x1888  :  255 - 0xff
    "11111111", -- 6281 - 0x1889  :  255 - 0xff
    "11111111", -- 6282 - 0x188a  :  255 - 0xff
    "11111111", -- 6283 - 0x188b  :  255 - 0xff
    "11111111", -- 6284 - 0x188c  :  255 - 0xff
    "11111111", -- 6285 - 0x188d  :  255 - 0xff
    "11111111", -- 6286 - 0x188e  :  255 - 0xff
    "11111111", -- 6287 - 0x188f  :  255 - 0xff
    "11111111", -- 6288 - 0x1890  :  255 - 0xff -- Background 0x89
    "11111111", -- 6289 - 0x1891  :  255 - 0xff
    "11111111", -- 6290 - 0x1892  :  255 - 0xff
    "11111111", -- 6291 - 0x1893  :  255 - 0xff
    "11111111", -- 6292 - 0x1894  :  255 - 0xff
    "11111111", -- 6293 - 0x1895  :  255 - 0xff
    "11111111", -- 6294 - 0x1896  :  255 - 0xff
    "11111111", -- 6295 - 0x1897  :  255 - 0xff
    "11111111", -- 6296 - 0x1898  :  255 - 0xff
    "11111111", -- 6297 - 0x1899  :  255 - 0xff
    "11111111", -- 6298 - 0x189a  :  255 - 0xff
    "11111111", -- 6299 - 0x189b  :  255 - 0xff
    "11111111", -- 6300 - 0x189c  :  255 - 0xff
    "11111111", -- 6301 - 0x189d  :  255 - 0xff
    "11111111", -- 6302 - 0x189e  :  255 - 0xff
    "11111111", -- 6303 - 0x189f  :  255 - 0xff
    "11111111", -- 6304 - 0x18a0  :  255 - 0xff -- Background 0x8a
    "11111111", -- 6305 - 0x18a1  :  255 - 0xff
    "11111111", -- 6306 - 0x18a2  :  255 - 0xff
    "11111111", -- 6307 - 0x18a3  :  255 - 0xff
    "11111111", -- 6308 - 0x18a4  :  255 - 0xff
    "11111111", -- 6309 - 0x18a5  :  255 - 0xff
    "11111111", -- 6310 - 0x18a6  :  255 - 0xff
    "11111111", -- 6311 - 0x18a7  :  255 - 0xff
    "11111111", -- 6312 - 0x18a8  :  255 - 0xff
    "11111111", -- 6313 - 0x18a9  :  255 - 0xff
    "11111111", -- 6314 - 0x18aa  :  255 - 0xff
    "11111111", -- 6315 - 0x18ab  :  255 - 0xff
    "11111111", -- 6316 - 0x18ac  :  255 - 0xff
    "11111111", -- 6317 - 0x18ad  :  255 - 0xff
    "11111111", -- 6318 - 0x18ae  :  255 - 0xff
    "11111111", -- 6319 - 0x18af  :  255 - 0xff
    "11111111", -- 6320 - 0x18b0  :  255 - 0xff -- Background 0x8b
    "11111111", -- 6321 - 0x18b1  :  255 - 0xff
    "11111111", -- 6322 - 0x18b2  :  255 - 0xff
    "11111111", -- 6323 - 0x18b3  :  255 - 0xff
    "11111111", -- 6324 - 0x18b4  :  255 - 0xff
    "11111111", -- 6325 - 0x18b5  :  255 - 0xff
    "11111111", -- 6326 - 0x18b6  :  255 - 0xff
    "11111111", -- 6327 - 0x18b7  :  255 - 0xff
    "11111111", -- 6328 - 0x18b8  :  255 - 0xff
    "11111111", -- 6329 - 0x18b9  :  255 - 0xff
    "11111111", -- 6330 - 0x18ba  :  255 - 0xff
    "11111111", -- 6331 - 0x18bb  :  255 - 0xff
    "11111111", -- 6332 - 0x18bc  :  255 - 0xff
    "11111111", -- 6333 - 0x18bd  :  255 - 0xff
    "11111111", -- 6334 - 0x18be  :  255 - 0xff
    "11111111", -- 6335 - 0x18bf  :  255 - 0xff
    "11111111", -- 6336 - 0x18c0  :  255 - 0xff -- Background 0x8c
    "11111111", -- 6337 - 0x18c1  :  255 - 0xff
    "11111111", -- 6338 - 0x18c2  :  255 - 0xff
    "11111111", -- 6339 - 0x18c3  :  255 - 0xff
    "11111111", -- 6340 - 0x18c4  :  255 - 0xff
    "11111111", -- 6341 - 0x18c5  :  255 - 0xff
    "11111111", -- 6342 - 0x18c6  :  255 - 0xff
    "11111111", -- 6343 - 0x18c7  :  255 - 0xff
    "11111111", -- 6344 - 0x18c8  :  255 - 0xff
    "11111111", -- 6345 - 0x18c9  :  255 - 0xff
    "11111111", -- 6346 - 0x18ca  :  255 - 0xff
    "11111111", -- 6347 - 0x18cb  :  255 - 0xff
    "11111111", -- 6348 - 0x18cc  :  255 - 0xff
    "11111111", -- 6349 - 0x18cd  :  255 - 0xff
    "11111111", -- 6350 - 0x18ce  :  255 - 0xff
    "11111111", -- 6351 - 0x18cf  :  255 - 0xff
    "11111111", -- 6352 - 0x18d0  :  255 - 0xff -- Background 0x8d
    "11111111", -- 6353 - 0x18d1  :  255 - 0xff
    "11111111", -- 6354 - 0x18d2  :  255 - 0xff
    "11111111", -- 6355 - 0x18d3  :  255 - 0xff
    "11111111", -- 6356 - 0x18d4  :  255 - 0xff
    "11111111", -- 6357 - 0x18d5  :  255 - 0xff
    "11111111", -- 6358 - 0x18d6  :  255 - 0xff
    "11111111", -- 6359 - 0x18d7  :  255 - 0xff
    "11111111", -- 6360 - 0x18d8  :  255 - 0xff
    "11111111", -- 6361 - 0x18d9  :  255 - 0xff
    "11111111", -- 6362 - 0x18da  :  255 - 0xff
    "11111111", -- 6363 - 0x18db  :  255 - 0xff
    "11111111", -- 6364 - 0x18dc  :  255 - 0xff
    "11111111", -- 6365 - 0x18dd  :  255 - 0xff
    "11111111", -- 6366 - 0x18de  :  255 - 0xff
    "11111111", -- 6367 - 0x18df  :  255 - 0xff
    "11111111", -- 6368 - 0x18e0  :  255 - 0xff -- Background 0x8e
    "11111111", -- 6369 - 0x18e1  :  255 - 0xff
    "11111111", -- 6370 - 0x18e2  :  255 - 0xff
    "11111111", -- 6371 - 0x18e3  :  255 - 0xff
    "11111111", -- 6372 - 0x18e4  :  255 - 0xff
    "11111111", -- 6373 - 0x18e5  :  255 - 0xff
    "11111111", -- 6374 - 0x18e6  :  255 - 0xff
    "11111111", -- 6375 - 0x18e7  :  255 - 0xff
    "11111111", -- 6376 - 0x18e8  :  255 - 0xff
    "11111111", -- 6377 - 0x18e9  :  255 - 0xff
    "11111111", -- 6378 - 0x18ea  :  255 - 0xff
    "11111111", -- 6379 - 0x18eb  :  255 - 0xff
    "11111111", -- 6380 - 0x18ec  :  255 - 0xff
    "11111111", -- 6381 - 0x18ed  :  255 - 0xff
    "11111111", -- 6382 - 0x18ee  :  255 - 0xff
    "11111111", -- 6383 - 0x18ef  :  255 - 0xff
    "11111111", -- 6384 - 0x18f0  :  255 - 0xff -- Background 0x8f
    "11111111", -- 6385 - 0x18f1  :  255 - 0xff
    "11111111", -- 6386 - 0x18f2  :  255 - 0xff
    "11111111", -- 6387 - 0x18f3  :  255 - 0xff
    "11111111", -- 6388 - 0x18f4  :  255 - 0xff
    "11111111", -- 6389 - 0x18f5  :  255 - 0xff
    "11111111", -- 6390 - 0x18f6  :  255 - 0xff
    "11111111", -- 6391 - 0x18f7  :  255 - 0xff
    "11111111", -- 6392 - 0x18f8  :  255 - 0xff
    "11111111", -- 6393 - 0x18f9  :  255 - 0xff
    "11111111", -- 6394 - 0x18fa  :  255 - 0xff
    "11111111", -- 6395 - 0x18fb  :  255 - 0xff
    "11111111", -- 6396 - 0x18fc  :  255 - 0xff
    "11111111", -- 6397 - 0x18fd  :  255 - 0xff
    "11111111", -- 6398 - 0x18fe  :  255 - 0xff
    "11111111", -- 6399 - 0x18ff  :  255 - 0xff
    "00000000", -- 6400 - 0x1900  :    0 - 0x0 -- Background 0x90
    "00000000", -- 6401 - 0x1901  :    0 - 0x0
    "00000000", -- 6402 - 0x1902  :    0 - 0x0
    "00000000", -- 6403 - 0x1903  :    0 - 0x0
    "00000000", -- 6404 - 0x1904  :    0 - 0x0
    "00000001", -- 6405 - 0x1905  :    1 - 0x1
    "00011110", -- 6406 - 0x1906  :   30 - 0x1e
    "00111011", -- 6407 - 0x1907  :   59 - 0x3b
    "00000000", -- 6408 - 0x1908  :    0 - 0x0
    "00000000", -- 6409 - 0x1909  :    0 - 0x0
    "00000000", -- 6410 - 0x190a  :    0 - 0x0
    "00000000", -- 6411 - 0x190b  :    0 - 0x0
    "00000000", -- 6412 - 0x190c  :    0 - 0x0
    "00000000", -- 6413 - 0x190d  :    0 - 0x0
    "00000000", -- 6414 - 0x190e  :    0 - 0x0
    "00000000", -- 6415 - 0x190f  :    0 - 0x0
    "00000000", -- 6416 - 0x1910  :    0 - 0x0 -- Background 0x91
    "00000000", -- 6417 - 0x1911  :    0 - 0x0
    "00001100", -- 6418 - 0x1912  :   12 - 0xc
    "00111100", -- 6419 - 0x1913  :   60 - 0x3c
    "11010000", -- 6420 - 0x1914  :  208 - 0xd0
    "00010000", -- 6421 - 0x1915  :   16 - 0x10
    "00100000", -- 6422 - 0x1916  :   32 - 0x20
    "01000000", -- 6423 - 0x1917  :   64 - 0x40
    "00000000", -- 6424 - 0x1918  :    0 - 0x0
    "00000000", -- 6425 - 0x1919  :    0 - 0x0
    "00000000", -- 6426 - 0x191a  :    0 - 0x0
    "00000000", -- 6427 - 0x191b  :    0 - 0x0
    "00000000", -- 6428 - 0x191c  :    0 - 0x0
    "00000000", -- 6429 - 0x191d  :    0 - 0x0
    "00000000", -- 6430 - 0x191e  :    0 - 0x0
    "00000000", -- 6431 - 0x191f  :    0 - 0x0
    "00111110", -- 6432 - 0x1920  :   62 - 0x3e -- Background 0x92
    "00101101", -- 6433 - 0x1921  :   45 - 0x2d
    "00110101", -- 6434 - 0x1922  :   53 - 0x35
    "00011101", -- 6435 - 0x1923  :   29 - 0x1d
    "00000001", -- 6436 - 0x1924  :    1 - 0x1
    "00000000", -- 6437 - 0x1925  :    0 - 0x0
    "00000000", -- 6438 - 0x1926  :    0 - 0x0
    "00000000", -- 6439 - 0x1927  :    0 - 0x0
    "00000000", -- 6440 - 0x1928  :    0 - 0x0
    "00000000", -- 6441 - 0x1929  :    0 - 0x0
    "00000000", -- 6442 - 0x192a  :    0 - 0x0
    "00000000", -- 6443 - 0x192b  :    0 - 0x0
    "00000000", -- 6444 - 0x192c  :    0 - 0x0
    "00000000", -- 6445 - 0x192d  :    0 - 0x0
    "00000000", -- 6446 - 0x192e  :    0 - 0x0
    "00000000", -- 6447 - 0x192f  :    0 - 0x0
    "10110000", -- 6448 - 0x1930  :  176 - 0xb0 -- Background 0x93
    "10111000", -- 6449 - 0x1931  :  184 - 0xb8
    "11111000", -- 6450 - 0x1932  :  248 - 0xf8
    "01111000", -- 6451 - 0x1933  :  120 - 0x78
    "10011000", -- 6452 - 0x1934  :  152 - 0x98
    "11110000", -- 6453 - 0x1935  :  240 - 0xf0
    "00000000", -- 6454 - 0x1936  :    0 - 0x0
    "00000000", -- 6455 - 0x1937  :    0 - 0x0
    "00000000", -- 6456 - 0x1938  :    0 - 0x0
    "00000000", -- 6457 - 0x1939  :    0 - 0x0
    "00000000", -- 6458 - 0x193a  :    0 - 0x0
    "00000000", -- 6459 - 0x193b  :    0 - 0x0
    "00000000", -- 6460 - 0x193c  :    0 - 0x0
    "00000000", -- 6461 - 0x193d  :    0 - 0x0
    "00000000", -- 6462 - 0x193e  :    0 - 0x0
    "00000000", -- 6463 - 0x193f  :    0 - 0x0
    "00000000", -- 6464 - 0x1940  :    0 - 0x0 -- Background 0x94
    "00000000", -- 6465 - 0x1941  :    0 - 0x0
    "00000111", -- 6466 - 0x1942  :    7 - 0x7
    "00000011", -- 6467 - 0x1943  :    3 - 0x3
    "00001101", -- 6468 - 0x1944  :   13 - 0xd
    "00011110", -- 6469 - 0x1945  :   30 - 0x1e
    "00010111", -- 6470 - 0x1946  :   23 - 0x17
    "00011101", -- 6471 - 0x1947  :   29 - 0x1d
    "00000000", -- 6472 - 0x1948  :    0 - 0x0
    "00000000", -- 6473 - 0x1949  :    0 - 0x0
    "00000000", -- 6474 - 0x194a  :    0 - 0x0
    "00000000", -- 6475 - 0x194b  :    0 - 0x0
    "00000000", -- 6476 - 0x194c  :    0 - 0x0
    "00000000", -- 6477 - 0x194d  :    0 - 0x0
    "00000000", -- 6478 - 0x194e  :    0 - 0x0
    "00000000", -- 6479 - 0x194f  :    0 - 0x0
    "00000000", -- 6480 - 0x1950  :    0 - 0x0 -- Background 0x95
    "10000000", -- 6481 - 0x1951  :  128 - 0x80
    "01110000", -- 6482 - 0x1952  :  112 - 0x70
    "11100000", -- 6483 - 0x1953  :  224 - 0xe0
    "11011000", -- 6484 - 0x1954  :  216 - 0xd8
    "10111100", -- 6485 - 0x1955  :  188 - 0xbc
    "01110100", -- 6486 - 0x1956  :  116 - 0x74
    "11011100", -- 6487 - 0x1957  :  220 - 0xdc
    "00000000", -- 6488 - 0x1958  :    0 - 0x0
    "00000000", -- 6489 - 0x1959  :    0 - 0x0
    "00000000", -- 6490 - 0x195a  :    0 - 0x0
    "00000000", -- 6491 - 0x195b  :    0 - 0x0
    "00000000", -- 6492 - 0x195c  :    0 - 0x0
    "00000000", -- 6493 - 0x195d  :    0 - 0x0
    "00000000", -- 6494 - 0x195e  :    0 - 0x0
    "00000000", -- 6495 - 0x195f  :    0 - 0x0
    "00011111", -- 6496 - 0x1960  :   31 - 0x1f -- Background 0x96
    "00001011", -- 6497 - 0x1961  :   11 - 0xb
    "00001111", -- 6498 - 0x1962  :   15 - 0xf
    "00000101", -- 6499 - 0x1963  :    5 - 0x5
    "00000011", -- 6500 - 0x1964  :    3 - 0x3
    "00000001", -- 6501 - 0x1965  :    1 - 0x1
    "00000000", -- 6502 - 0x1966  :    0 - 0x0
    "00000000", -- 6503 - 0x1967  :    0 - 0x0
    "00000000", -- 6504 - 0x1968  :    0 - 0x0
    "00000000", -- 6505 - 0x1969  :    0 - 0x0
    "00000000", -- 6506 - 0x196a  :    0 - 0x0
    "00000000", -- 6507 - 0x196b  :    0 - 0x0
    "00000000", -- 6508 - 0x196c  :    0 - 0x0
    "00000000", -- 6509 - 0x196d  :    0 - 0x0
    "00000000", -- 6510 - 0x196e  :    0 - 0x0
    "00000000", -- 6511 - 0x196f  :    0 - 0x0
    "11111100", -- 6512 - 0x1970  :  252 - 0xfc -- Background 0x97
    "01101000", -- 6513 - 0x1971  :  104 - 0x68
    "11111000", -- 6514 - 0x1972  :  248 - 0xf8
    "10110000", -- 6515 - 0x1973  :  176 - 0xb0
    "11100000", -- 6516 - 0x1974  :  224 - 0xe0
    "10000000", -- 6517 - 0x1975  :  128 - 0x80
    "00000000", -- 6518 - 0x1976  :    0 - 0x0
    "00000000", -- 6519 - 0x1977  :    0 - 0x0
    "00000000", -- 6520 - 0x1978  :    0 - 0x0
    "00000000", -- 6521 - 0x1979  :    0 - 0x0
    "00000000", -- 6522 - 0x197a  :    0 - 0x0
    "00000000", -- 6523 - 0x197b  :    0 - 0x0
    "00000000", -- 6524 - 0x197c  :    0 - 0x0
    "00000000", -- 6525 - 0x197d  :    0 - 0x0
    "00000000", -- 6526 - 0x197e  :    0 - 0x0
    "00000000", -- 6527 - 0x197f  :    0 - 0x0
    "00000000", -- 6528 - 0x1980  :    0 - 0x0 -- Background 0x98
    "00000000", -- 6529 - 0x1981  :    0 - 0x0
    "00000000", -- 6530 - 0x1982  :    0 - 0x0
    "00000001", -- 6531 - 0x1983  :    1 - 0x1
    "00000001", -- 6532 - 0x1984  :    1 - 0x1
    "00001011", -- 6533 - 0x1985  :   11 - 0xb
    "00011100", -- 6534 - 0x1986  :   28 - 0x1c
    "00111111", -- 6535 - 0x1987  :   63 - 0x3f
    "00000000", -- 6536 - 0x1988  :    0 - 0x0
    "00000000", -- 6537 - 0x1989  :    0 - 0x0
    "00000000", -- 6538 - 0x198a  :    0 - 0x0
    "00000000", -- 6539 - 0x198b  :    0 - 0x0
    "00000000", -- 6540 - 0x198c  :    0 - 0x0
    "00000000", -- 6541 - 0x198d  :    0 - 0x0
    "00000000", -- 6542 - 0x198e  :    0 - 0x0
    "00000000", -- 6543 - 0x198f  :    0 - 0x0
    "00000000", -- 6544 - 0x1990  :    0 - 0x0 -- Background 0x99
    "00000000", -- 6545 - 0x1991  :    0 - 0x0
    "00110000", -- 6546 - 0x1992  :   48 - 0x30
    "01111000", -- 6547 - 0x1993  :  120 - 0x78
    "10000000", -- 6548 - 0x1994  :  128 - 0x80
    "11110000", -- 6549 - 0x1995  :  240 - 0xf0
    "11111000", -- 6550 - 0x1996  :  248 - 0xf8
    "11111100", -- 6551 - 0x1997  :  252 - 0xfc
    "00000000", -- 6552 - 0x1998  :    0 - 0x0
    "00000000", -- 6553 - 0x1999  :    0 - 0x0
    "00000000", -- 6554 - 0x199a  :    0 - 0x0
    "00000000", -- 6555 - 0x199b  :    0 - 0x0
    "00000000", -- 6556 - 0x199c  :    0 - 0x0
    "00000000", -- 6557 - 0x199d  :    0 - 0x0
    "00000000", -- 6558 - 0x199e  :    0 - 0x0
    "00000000", -- 6559 - 0x199f  :    0 - 0x0
    "00111111", -- 6560 - 0x19a0  :   63 - 0x3f -- Background 0x9a
    "00111111", -- 6561 - 0x19a1  :   63 - 0x3f
    "00111111", -- 6562 - 0x19a2  :   63 - 0x3f
    "00011111", -- 6563 - 0x19a3  :   31 - 0x1f
    "00011111", -- 6564 - 0x19a4  :   31 - 0x1f
    "00000111", -- 6565 - 0x19a5  :    7 - 0x7
    "00000000", -- 6566 - 0x19a6  :    0 - 0x0
    "00000000", -- 6567 - 0x19a7  :    0 - 0x0
    "00000000", -- 6568 - 0x19a8  :    0 - 0x0
    "00000000", -- 6569 - 0x19a9  :    0 - 0x0
    "00000000", -- 6570 - 0x19aa  :    0 - 0x0
    "00000000", -- 6571 - 0x19ab  :    0 - 0x0
    "00000000", -- 6572 - 0x19ac  :    0 - 0x0
    "00000000", -- 6573 - 0x19ad  :    0 - 0x0
    "00000000", -- 6574 - 0x19ae  :    0 - 0x0
    "00000000", -- 6575 - 0x19af  :    0 - 0x0
    "11111100", -- 6576 - 0x19b0  :  252 - 0xfc -- Background 0x9b
    "11101100", -- 6577 - 0x19b1  :  236 - 0xec
    "11101100", -- 6578 - 0x19b2  :  236 - 0xec
    "11011000", -- 6579 - 0x19b3  :  216 - 0xd8
    "11111000", -- 6580 - 0x19b4  :  248 - 0xf8
    "11100000", -- 6581 - 0x19b5  :  224 - 0xe0
    "00000000", -- 6582 - 0x19b6  :    0 - 0x0
    "00000000", -- 6583 - 0x19b7  :    0 - 0x0
    "00000000", -- 6584 - 0x19b8  :    0 - 0x0
    "00000000", -- 6585 - 0x19b9  :    0 - 0x0
    "00000000", -- 6586 - 0x19ba  :    0 - 0x0
    "00000000", -- 6587 - 0x19bb  :    0 - 0x0
    "00000000", -- 6588 - 0x19bc  :    0 - 0x0
    "00000000", -- 6589 - 0x19bd  :    0 - 0x0
    "00000000", -- 6590 - 0x19be  :    0 - 0x0
    "00000000", -- 6591 - 0x19bf  :    0 - 0x0
    "00000000", -- 6592 - 0x19c0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 6593 - 0x19c1  :    0 - 0x0
    "00000001", -- 6594 - 0x19c2  :    1 - 0x1
    "00011101", -- 6595 - 0x19c3  :   29 - 0x1d
    "00111110", -- 6596 - 0x19c4  :   62 - 0x3e
    "00111111", -- 6597 - 0x19c5  :   63 - 0x3f
    "00111111", -- 6598 - 0x19c6  :   63 - 0x3f
    "00111111", -- 6599 - 0x19c7  :   63 - 0x3f
    "00000000", -- 6600 - 0x19c8  :    0 - 0x0
    "00000000", -- 6601 - 0x19c9  :    0 - 0x0
    "00000000", -- 6602 - 0x19ca  :    0 - 0x0
    "00000000", -- 6603 - 0x19cb  :    0 - 0x0
    "00000000", -- 6604 - 0x19cc  :    0 - 0x0
    "00000000", -- 6605 - 0x19cd  :    0 - 0x0
    "00000000", -- 6606 - 0x19ce  :    0 - 0x0
    "00000000", -- 6607 - 0x19cf  :    0 - 0x0
    "00000000", -- 6608 - 0x19d0  :    0 - 0x0 -- Background 0x9d
    "10000000", -- 6609 - 0x19d1  :  128 - 0x80
    "00000000", -- 6610 - 0x19d2  :    0 - 0x0
    "01110000", -- 6611 - 0x19d3  :  112 - 0x70
    "11111000", -- 6612 - 0x19d4  :  248 - 0xf8
    "11111100", -- 6613 - 0x19d5  :  252 - 0xfc
    "11111100", -- 6614 - 0x19d6  :  252 - 0xfc
    "11111100", -- 6615 - 0x19d7  :  252 - 0xfc
    "00000000", -- 6616 - 0x19d8  :    0 - 0x0
    "00000000", -- 6617 - 0x19d9  :    0 - 0x0
    "00000000", -- 6618 - 0x19da  :    0 - 0x0
    "00000000", -- 6619 - 0x19db  :    0 - 0x0
    "00000000", -- 6620 - 0x19dc  :    0 - 0x0
    "00000000", -- 6621 - 0x19dd  :    0 - 0x0
    "00000000", -- 6622 - 0x19de  :    0 - 0x0
    "00000000", -- 6623 - 0x19df  :    0 - 0x0
    "00111111", -- 6624 - 0x19e0  :   63 - 0x3f -- Background 0x9e
    "00111111", -- 6625 - 0x19e1  :   63 - 0x3f
    "00011111", -- 6626 - 0x19e2  :   31 - 0x1f
    "00011111", -- 6627 - 0x19e3  :   31 - 0x1f
    "00001111", -- 6628 - 0x19e4  :   15 - 0xf
    "00000110", -- 6629 - 0x19e5  :    6 - 0x6
    "00000000", -- 6630 - 0x19e6  :    0 - 0x0
    "00000000", -- 6631 - 0x19e7  :    0 - 0x0
    "00000000", -- 6632 - 0x19e8  :    0 - 0x0
    "00000000", -- 6633 - 0x19e9  :    0 - 0x0
    "00000000", -- 6634 - 0x19ea  :    0 - 0x0
    "00000000", -- 6635 - 0x19eb  :    0 - 0x0
    "00000000", -- 6636 - 0x19ec  :    0 - 0x0
    "00000000", -- 6637 - 0x19ed  :    0 - 0x0
    "00000000", -- 6638 - 0x19ee  :    0 - 0x0
    "00000000", -- 6639 - 0x19ef  :    0 - 0x0
    "11101100", -- 6640 - 0x19f0  :  236 - 0xec -- Background 0x9f
    "11101100", -- 6641 - 0x19f1  :  236 - 0xec
    "11011000", -- 6642 - 0x19f2  :  216 - 0xd8
    "11111000", -- 6643 - 0x19f3  :  248 - 0xf8
    "11110000", -- 6644 - 0x19f4  :  240 - 0xf0
    "11100000", -- 6645 - 0x19f5  :  224 - 0xe0
    "00000000", -- 6646 - 0x19f6  :    0 - 0x0
    "00000000", -- 6647 - 0x19f7  :    0 - 0x0
    "00000000", -- 6648 - 0x19f8  :    0 - 0x0
    "00000000", -- 6649 - 0x19f9  :    0 - 0x0
    "00000000", -- 6650 - 0x19fa  :    0 - 0x0
    "00000000", -- 6651 - 0x19fb  :    0 - 0x0
    "00000000", -- 6652 - 0x19fc  :    0 - 0x0
    "00000000", -- 6653 - 0x19fd  :    0 - 0x0
    "00000000", -- 6654 - 0x19fe  :    0 - 0x0
    "00000000", -- 6655 - 0x19ff  :    0 - 0x0
    "00000000", -- 6656 - 0x1a00  :    0 - 0x0 -- Background 0xa0
    "00000100", -- 6657 - 0x1a01  :    4 - 0x4
    "00000011", -- 6658 - 0x1a02  :    3 - 0x3
    "00000000", -- 6659 - 0x1a03  :    0 - 0x0
    "00000001", -- 6660 - 0x1a04  :    1 - 0x1
    "00000111", -- 6661 - 0x1a05  :    7 - 0x7
    "00001111", -- 6662 - 0x1a06  :   15 - 0xf
    "00001100", -- 6663 - 0x1a07  :   12 - 0xc
    "00000000", -- 6664 - 0x1a08  :    0 - 0x0
    "00000000", -- 6665 - 0x1a09  :    0 - 0x0
    "00000000", -- 6666 - 0x1a0a  :    0 - 0x0
    "00000000", -- 6667 - 0x1a0b  :    0 - 0x0
    "00000000", -- 6668 - 0x1a0c  :    0 - 0x0
    "00000000", -- 6669 - 0x1a0d  :    0 - 0x0
    "00000000", -- 6670 - 0x1a0e  :    0 - 0x0
    "00000000", -- 6671 - 0x1a0f  :    0 - 0x0
    "00000000", -- 6672 - 0x1a10  :    0 - 0x0 -- Background 0xa1
    "00000000", -- 6673 - 0x1a11  :    0 - 0x0
    "11100000", -- 6674 - 0x1a12  :  224 - 0xe0
    "10000000", -- 6675 - 0x1a13  :  128 - 0x80
    "01000000", -- 6676 - 0x1a14  :   64 - 0x40
    "11110000", -- 6677 - 0x1a15  :  240 - 0xf0
    "10011000", -- 6678 - 0x1a16  :  152 - 0x98
    "11111000", -- 6679 - 0x1a17  :  248 - 0xf8
    "00000000", -- 6680 - 0x1a18  :    0 - 0x0
    "00000000", -- 6681 - 0x1a19  :    0 - 0x0
    "00000000", -- 6682 - 0x1a1a  :    0 - 0x0
    "00000000", -- 6683 - 0x1a1b  :    0 - 0x0
    "00000000", -- 6684 - 0x1a1c  :    0 - 0x0
    "00000000", -- 6685 - 0x1a1d  :    0 - 0x0
    "00000000", -- 6686 - 0x1a1e  :    0 - 0x0
    "00000000", -- 6687 - 0x1a1f  :    0 - 0x0
    "00011111", -- 6688 - 0x1a20  :   31 - 0x1f -- Background 0xa2
    "00010011", -- 6689 - 0x1a21  :   19 - 0x13
    "00011111", -- 6690 - 0x1a22  :   31 - 0x1f
    "00001111", -- 6691 - 0x1a23  :   15 - 0xf
    "00001001", -- 6692 - 0x1a24  :    9 - 0x9
    "00000111", -- 6693 - 0x1a25  :    7 - 0x7
    "00000001", -- 6694 - 0x1a26  :    1 - 0x1
    "00000000", -- 6695 - 0x1a27  :    0 - 0x0
    "00000000", -- 6696 - 0x1a28  :    0 - 0x0
    "00000000", -- 6697 - 0x1a29  :    0 - 0x0
    "00000000", -- 6698 - 0x1a2a  :    0 - 0x0
    "00000000", -- 6699 - 0x1a2b  :    0 - 0x0
    "00000000", -- 6700 - 0x1a2c  :    0 - 0x0
    "00000000", -- 6701 - 0x1a2d  :    0 - 0x0
    "00000000", -- 6702 - 0x1a2e  :    0 - 0x0
    "00000000", -- 6703 - 0x1a2f  :    0 - 0x0
    "11100100", -- 6704 - 0x1a30  :  228 - 0xe4 -- Background 0xa3
    "00111100", -- 6705 - 0x1a31  :   60 - 0x3c
    "11100100", -- 6706 - 0x1a32  :  228 - 0xe4
    "00111000", -- 6707 - 0x1a33  :   56 - 0x38
    "11111000", -- 6708 - 0x1a34  :  248 - 0xf8
    "11110000", -- 6709 - 0x1a35  :  240 - 0xf0
    "11000000", -- 6710 - 0x1a36  :  192 - 0xc0
    "00000000", -- 6711 - 0x1a37  :    0 - 0x0
    "00000000", -- 6712 - 0x1a38  :    0 - 0x0
    "00000000", -- 6713 - 0x1a39  :    0 - 0x0
    "00000000", -- 6714 - 0x1a3a  :    0 - 0x0
    "00000000", -- 6715 - 0x1a3b  :    0 - 0x0
    "00000000", -- 6716 - 0x1a3c  :    0 - 0x0
    "00000000", -- 6717 - 0x1a3d  :    0 - 0x0
    "00000000", -- 6718 - 0x1a3e  :    0 - 0x0
    "00000000", -- 6719 - 0x1a3f  :    0 - 0x0
    "00000000", -- 6720 - 0x1a40  :    0 - 0x0 -- Background 0xa4
    "00000000", -- 6721 - 0x1a41  :    0 - 0x0
    "00000000", -- 6722 - 0x1a42  :    0 - 0x0
    "00000000", -- 6723 - 0x1a43  :    0 - 0x0
    "00010001", -- 6724 - 0x1a44  :   17 - 0x11
    "00010011", -- 6725 - 0x1a45  :   19 - 0x13
    "00011111", -- 6726 - 0x1a46  :   31 - 0x1f
    "00011111", -- 6727 - 0x1a47  :   31 - 0x1f
    "00000000", -- 6728 - 0x1a48  :    0 - 0x0
    "00000000", -- 6729 - 0x1a49  :    0 - 0x0
    "00000000", -- 6730 - 0x1a4a  :    0 - 0x0
    "00000000", -- 6731 - 0x1a4b  :    0 - 0x0
    "00000000", -- 6732 - 0x1a4c  :    0 - 0x0
    "00000000", -- 6733 - 0x1a4d  :    0 - 0x0
    "00000000", -- 6734 - 0x1a4e  :    0 - 0x0
    "00000000", -- 6735 - 0x1a4f  :    0 - 0x0
    "00000000", -- 6736 - 0x1a50  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 6737 - 0x1a51  :    0 - 0x0
    "00000000", -- 6738 - 0x1a52  :    0 - 0x0
    "10000000", -- 6739 - 0x1a53  :  128 - 0x80
    "11000100", -- 6740 - 0x1a54  :  196 - 0xc4
    "11100100", -- 6741 - 0x1a55  :  228 - 0xe4
    "11111100", -- 6742 - 0x1a56  :  252 - 0xfc
    "11111100", -- 6743 - 0x1a57  :  252 - 0xfc
    "00000000", -- 6744 - 0x1a58  :    0 - 0x0
    "00000000", -- 6745 - 0x1a59  :    0 - 0x0
    "00000000", -- 6746 - 0x1a5a  :    0 - 0x0
    "00000000", -- 6747 - 0x1a5b  :    0 - 0x0
    "00000000", -- 6748 - 0x1a5c  :    0 - 0x0
    "00000000", -- 6749 - 0x1a5d  :    0 - 0x0
    "00000000", -- 6750 - 0x1a5e  :    0 - 0x0
    "00000000", -- 6751 - 0x1a5f  :    0 - 0x0
    "00011111", -- 6752 - 0x1a60  :   31 - 0x1f -- Background 0xa6
    "00001110", -- 6753 - 0x1a61  :   14 - 0xe
    "00000110", -- 6754 - 0x1a62  :    6 - 0x6
    "00000010", -- 6755 - 0x1a63  :    2 - 0x2
    "00000000", -- 6756 - 0x1a64  :    0 - 0x0
    "00000000", -- 6757 - 0x1a65  :    0 - 0x0
    "00000000", -- 6758 - 0x1a66  :    0 - 0x0
    "00000000", -- 6759 - 0x1a67  :    0 - 0x0
    "00000000", -- 6760 - 0x1a68  :    0 - 0x0
    "00000000", -- 6761 - 0x1a69  :    0 - 0x0
    "00000000", -- 6762 - 0x1a6a  :    0 - 0x0
    "00000000", -- 6763 - 0x1a6b  :    0 - 0x0
    "00000000", -- 6764 - 0x1a6c  :    0 - 0x0
    "00000000", -- 6765 - 0x1a6d  :    0 - 0x0
    "00000000", -- 6766 - 0x1a6e  :    0 - 0x0
    "00000000", -- 6767 - 0x1a6f  :    0 - 0x0
    "11111100", -- 6768 - 0x1a70  :  252 - 0xfc -- Background 0xa7
    "10111000", -- 6769 - 0x1a71  :  184 - 0xb8
    "10110000", -- 6770 - 0x1a72  :  176 - 0xb0
    "10100000", -- 6771 - 0x1a73  :  160 - 0xa0
    "10000000", -- 6772 - 0x1a74  :  128 - 0x80
    "00000000", -- 6773 - 0x1a75  :    0 - 0x0
    "00000000", -- 6774 - 0x1a76  :    0 - 0x0
    "00000000", -- 6775 - 0x1a77  :    0 - 0x0
    "00000000", -- 6776 - 0x1a78  :    0 - 0x0
    "00000000", -- 6777 - 0x1a79  :    0 - 0x0
    "00000000", -- 6778 - 0x1a7a  :    0 - 0x0
    "00000000", -- 6779 - 0x1a7b  :    0 - 0x0
    "00000000", -- 6780 - 0x1a7c  :    0 - 0x0
    "00000000", -- 6781 - 0x1a7d  :    0 - 0x0
    "00000000", -- 6782 - 0x1a7e  :    0 - 0x0
    "00000000", -- 6783 - 0x1a7f  :    0 - 0x0
    "00000000", -- 6784 - 0x1a80  :    0 - 0x0 -- Background 0xa8
    "00000000", -- 6785 - 0x1a81  :    0 - 0x0
    "00000000", -- 6786 - 0x1a82  :    0 - 0x0
    "00000001", -- 6787 - 0x1a83  :    1 - 0x1
    "00000011", -- 6788 - 0x1a84  :    3 - 0x3
    "00000110", -- 6789 - 0x1a85  :    6 - 0x6
    "00000110", -- 6790 - 0x1a86  :    6 - 0x6
    "00001111", -- 6791 - 0x1a87  :   15 - 0xf
    "00000000", -- 6792 - 0x1a88  :    0 - 0x0
    "00000000", -- 6793 - 0x1a89  :    0 - 0x0
    "00000000", -- 6794 - 0x1a8a  :    0 - 0x0
    "00000000", -- 6795 - 0x1a8b  :    0 - 0x0
    "00000000", -- 6796 - 0x1a8c  :    0 - 0x0
    "00000000", -- 6797 - 0x1a8d  :    0 - 0x0
    "00000000", -- 6798 - 0x1a8e  :    0 - 0x0
    "00000000", -- 6799 - 0x1a8f  :    0 - 0x0
    "00000000", -- 6800 - 0x1a90  :    0 - 0x0 -- Background 0xa9
    "00011000", -- 6801 - 0x1a91  :   24 - 0x18
    "11110100", -- 6802 - 0x1a92  :  244 - 0xf4
    "11111000", -- 6803 - 0x1a93  :  248 - 0xf8
    "00111000", -- 6804 - 0x1a94  :   56 - 0x38
    "01111100", -- 6805 - 0x1a95  :  124 - 0x7c
    "11111100", -- 6806 - 0x1a96  :  252 - 0xfc
    "11111100", -- 6807 - 0x1a97  :  252 - 0xfc
    "00000000", -- 6808 - 0x1a98  :    0 - 0x0
    "00000000", -- 6809 - 0x1a99  :    0 - 0x0
    "00000000", -- 6810 - 0x1a9a  :    0 - 0x0
    "00000000", -- 6811 - 0x1a9b  :    0 - 0x0
    "00000000", -- 6812 - 0x1a9c  :    0 - 0x0
    "00000000", -- 6813 - 0x1a9d  :    0 - 0x0
    "00000000", -- 6814 - 0x1a9e  :    0 - 0x0
    "00000000", -- 6815 - 0x1a9f  :    0 - 0x0
    "00001111", -- 6816 - 0x1aa0  :   15 - 0xf -- Background 0xaa
    "00011111", -- 6817 - 0x1aa1  :   31 - 0x1f
    "00110000", -- 6818 - 0x1aa2  :   48 - 0x30
    "00111000", -- 6819 - 0x1aa3  :   56 - 0x38
    "00011101", -- 6820 - 0x1aa4  :   29 - 0x1d
    "00000011", -- 6821 - 0x1aa5  :    3 - 0x3
    "00000011", -- 6822 - 0x1aa6  :    3 - 0x3
    "00000000", -- 6823 - 0x1aa7  :    0 - 0x0
    "00000000", -- 6824 - 0x1aa8  :    0 - 0x0
    "00000000", -- 6825 - 0x1aa9  :    0 - 0x0
    "00000000", -- 6826 - 0x1aaa  :    0 - 0x0
    "00000000", -- 6827 - 0x1aab  :    0 - 0x0
    "00000000", -- 6828 - 0x1aac  :    0 - 0x0
    "00000000", -- 6829 - 0x1aad  :    0 - 0x0
    "00000000", -- 6830 - 0x1aae  :    0 - 0x0
    "00000000", -- 6831 - 0x1aaf  :    0 - 0x0
    "11111100", -- 6832 - 0x1ab0  :  252 - 0xfc -- Background 0xab
    "11111100", -- 6833 - 0x1ab1  :  252 - 0xfc
    "01111100", -- 6834 - 0x1ab2  :  124 - 0x7c
    "10001110", -- 6835 - 0x1ab3  :  142 - 0x8e
    "10000110", -- 6836 - 0x1ab4  :  134 - 0x86
    "10011100", -- 6837 - 0x1ab5  :  156 - 0x9c
    "01111000", -- 6838 - 0x1ab6  :  120 - 0x78
    "00000000", -- 6839 - 0x1ab7  :    0 - 0x0
    "00000000", -- 6840 - 0x1ab8  :    0 - 0x0
    "00000000", -- 6841 - 0x1ab9  :    0 - 0x0
    "00000000", -- 6842 - 0x1aba  :    0 - 0x0
    "00000000", -- 6843 - 0x1abb  :    0 - 0x0
    "00000000", -- 6844 - 0x1abc  :    0 - 0x0
    "00000000", -- 6845 - 0x1abd  :    0 - 0x0
    "00000000", -- 6846 - 0x1abe  :    0 - 0x0
    "00000000", -- 6847 - 0x1abf  :    0 - 0x0
    "00000000", -- 6848 - 0x1ac0  :    0 - 0x0 -- Background 0xac
    "00000001", -- 6849 - 0x1ac1  :    1 - 0x1
    "00000110", -- 6850 - 0x1ac2  :    6 - 0x6
    "00000111", -- 6851 - 0x1ac3  :    7 - 0x7
    "00000111", -- 6852 - 0x1ac4  :    7 - 0x7
    "00000111", -- 6853 - 0x1ac5  :    7 - 0x7
    "00000001", -- 6854 - 0x1ac6  :    1 - 0x1
    "00000011", -- 6855 - 0x1ac7  :    3 - 0x3
    "00000000", -- 6856 - 0x1ac8  :    0 - 0x0
    "00000000", -- 6857 - 0x1ac9  :    0 - 0x0
    "00000000", -- 6858 - 0x1aca  :    0 - 0x0
    "00000000", -- 6859 - 0x1acb  :    0 - 0x0
    "00000000", -- 6860 - 0x1acc  :    0 - 0x0
    "00000000", -- 6861 - 0x1acd  :    0 - 0x0
    "00000000", -- 6862 - 0x1ace  :    0 - 0x0
    "00000000", -- 6863 - 0x1acf  :    0 - 0x0
    "00000000", -- 6864 - 0x1ad0  :    0 - 0x0 -- Background 0xad
    "11000000", -- 6865 - 0x1ad1  :  192 - 0xc0
    "00110000", -- 6866 - 0x1ad2  :   48 - 0x30
    "11110000", -- 6867 - 0x1ad3  :  240 - 0xf0
    "11110000", -- 6868 - 0x1ad4  :  240 - 0xf0
    "11110000", -- 6869 - 0x1ad5  :  240 - 0xf0
    "01000000", -- 6870 - 0x1ad6  :   64 - 0x40
    "01000000", -- 6871 - 0x1ad7  :   64 - 0x40
    "00000000", -- 6872 - 0x1ad8  :    0 - 0x0
    "00000000", -- 6873 - 0x1ad9  :    0 - 0x0
    "00000000", -- 6874 - 0x1ada  :    0 - 0x0
    "00000000", -- 6875 - 0x1adb  :    0 - 0x0
    "00000000", -- 6876 - 0x1adc  :    0 - 0x0
    "00000000", -- 6877 - 0x1add  :    0 - 0x0
    "00000000", -- 6878 - 0x1ade  :    0 - 0x0
    "00000000", -- 6879 - 0x1adf  :    0 - 0x0
    "00000001", -- 6880 - 0x1ae0  :    1 - 0x1 -- Background 0xae
    "00000000", -- 6881 - 0x1ae1  :    0 - 0x0
    "00000001", -- 6882 - 0x1ae2  :    1 - 0x1
    "00000011", -- 6883 - 0x1ae3  :    3 - 0x3
    "00000001", -- 6884 - 0x1ae4  :    1 - 0x1
    "00000000", -- 6885 - 0x1ae5  :    0 - 0x0
    "00000000", -- 6886 - 0x1ae6  :    0 - 0x0
    "00000000", -- 6887 - 0x1ae7  :    0 - 0x0
    "00000000", -- 6888 - 0x1ae8  :    0 - 0x0
    "00000000", -- 6889 - 0x1ae9  :    0 - 0x0
    "00000000", -- 6890 - 0x1aea  :    0 - 0x0
    "00000000", -- 6891 - 0x1aeb  :    0 - 0x0
    "00000000", -- 6892 - 0x1aec  :    0 - 0x0
    "00000000", -- 6893 - 0x1aed  :    0 - 0x0
    "00000000", -- 6894 - 0x1aee  :    0 - 0x0
    "00000000", -- 6895 - 0x1aef  :    0 - 0x0
    "01000000", -- 6896 - 0x1af0  :   64 - 0x40 -- Background 0xaf
    "01000000", -- 6897 - 0x1af1  :   64 - 0x40
    "01000000", -- 6898 - 0x1af2  :   64 - 0x40
    "01000000", -- 6899 - 0x1af3  :   64 - 0x40
    "01000000", -- 6900 - 0x1af4  :   64 - 0x40
    "10000000", -- 6901 - 0x1af5  :  128 - 0x80
    "00000000", -- 6902 - 0x1af6  :    0 - 0x0
    "00000000", -- 6903 - 0x1af7  :    0 - 0x0
    "00000000", -- 6904 - 0x1af8  :    0 - 0x0
    "00000000", -- 6905 - 0x1af9  :    0 - 0x0
    "00000000", -- 6906 - 0x1afa  :    0 - 0x0
    "00000000", -- 6907 - 0x1afb  :    0 - 0x0
    "00000000", -- 6908 - 0x1afc  :    0 - 0x0
    "00000000", -- 6909 - 0x1afd  :    0 - 0x0
    "00000000", -- 6910 - 0x1afe  :    0 - 0x0
    "00000000", -- 6911 - 0x1aff  :    0 - 0x0
    "01111110", -- 6912 - 0x1b00  :  126 - 0x7e -- Background 0xb0
    "01100011", -- 6913 - 0x1b01  :   99 - 0x63
    "01100011", -- 6914 - 0x1b02  :   99 - 0x63
    "01100011", -- 6915 - 0x1b03  :   99 - 0x63
    "01111110", -- 6916 - 0x1b04  :  126 - 0x7e
    "01100000", -- 6917 - 0x1b05  :   96 - 0x60
    "01100000", -- 6918 - 0x1b06  :   96 - 0x60
    "00000000", -- 6919 - 0x1b07  :    0 - 0x0
    "01111110", -- 6920 - 0x1b08  :  126 - 0x7e
    "01100011", -- 6921 - 0x1b09  :   99 - 0x63
    "01100011", -- 6922 - 0x1b0a  :   99 - 0x63
    "01100011", -- 6923 - 0x1b0b  :   99 - 0x63
    "01111110", -- 6924 - 0x1b0c  :  126 - 0x7e
    "01100000", -- 6925 - 0x1b0d  :   96 - 0x60
    "01100000", -- 6926 - 0x1b0e  :   96 - 0x60
    "00000000", -- 6927 - 0x1b0f  :    0 - 0x0
    "01100000", -- 6928 - 0x1b10  :   96 - 0x60 -- Background 0xb1
    "01100000", -- 6929 - 0x1b11  :   96 - 0x60
    "01100000", -- 6930 - 0x1b12  :   96 - 0x60
    "01100000", -- 6931 - 0x1b13  :   96 - 0x60
    "01100000", -- 6932 - 0x1b14  :   96 - 0x60
    "01100000", -- 6933 - 0x1b15  :   96 - 0x60
    "01111111", -- 6934 - 0x1b16  :  127 - 0x7f
    "00000000", -- 6935 - 0x1b17  :    0 - 0x0
    "01100000", -- 6936 - 0x1b18  :   96 - 0x60
    "01100000", -- 6937 - 0x1b19  :   96 - 0x60
    "01100000", -- 6938 - 0x1b1a  :   96 - 0x60
    "01100000", -- 6939 - 0x1b1b  :   96 - 0x60
    "01100000", -- 6940 - 0x1b1c  :   96 - 0x60
    "01100000", -- 6941 - 0x1b1d  :   96 - 0x60
    "01111111", -- 6942 - 0x1b1e  :  127 - 0x7f
    "00000000", -- 6943 - 0x1b1f  :    0 - 0x0
    "00011100", -- 6944 - 0x1b20  :   28 - 0x1c -- Background 0xb2
    "00110110", -- 6945 - 0x1b21  :   54 - 0x36
    "01100011", -- 6946 - 0x1b22  :   99 - 0x63
    "01100011", -- 6947 - 0x1b23  :   99 - 0x63
    "01111111", -- 6948 - 0x1b24  :  127 - 0x7f
    "01100011", -- 6949 - 0x1b25  :   99 - 0x63
    "01100011", -- 6950 - 0x1b26  :   99 - 0x63
    "00000000", -- 6951 - 0x1b27  :    0 - 0x0
    "00011100", -- 6952 - 0x1b28  :   28 - 0x1c
    "00110110", -- 6953 - 0x1b29  :   54 - 0x36
    "01100011", -- 6954 - 0x1b2a  :   99 - 0x63
    "01100011", -- 6955 - 0x1b2b  :   99 - 0x63
    "01111111", -- 6956 - 0x1b2c  :  127 - 0x7f
    "01100011", -- 6957 - 0x1b2d  :   99 - 0x63
    "01100011", -- 6958 - 0x1b2e  :   99 - 0x63
    "00000000", -- 6959 - 0x1b2f  :    0 - 0x0
    "00110011", -- 6960 - 0x1b30  :   51 - 0x33 -- Background 0xb3
    "00110011", -- 6961 - 0x1b31  :   51 - 0x33
    "00110011", -- 6962 - 0x1b32  :   51 - 0x33
    "00011110", -- 6963 - 0x1b33  :   30 - 0x1e
    "00001100", -- 6964 - 0x1b34  :   12 - 0xc
    "00001100", -- 6965 - 0x1b35  :   12 - 0xc
    "00001100", -- 6966 - 0x1b36  :   12 - 0xc
    "00000000", -- 6967 - 0x1b37  :    0 - 0x0
    "00110011", -- 6968 - 0x1b38  :   51 - 0x33
    "00110011", -- 6969 - 0x1b39  :   51 - 0x33
    "00110011", -- 6970 - 0x1b3a  :   51 - 0x33
    "00011110", -- 6971 - 0x1b3b  :   30 - 0x1e
    "00001100", -- 6972 - 0x1b3c  :   12 - 0xc
    "00001100", -- 6973 - 0x1b3d  :   12 - 0xc
    "00001100", -- 6974 - 0x1b3e  :   12 - 0xc
    "00000000", -- 6975 - 0x1b3f  :    0 - 0x0
    "01111111", -- 6976 - 0x1b40  :  127 - 0x7f -- Background 0xb4
    "01100000", -- 6977 - 0x1b41  :   96 - 0x60
    "01100000", -- 6978 - 0x1b42  :   96 - 0x60
    "01111110", -- 6979 - 0x1b43  :  126 - 0x7e
    "01100000", -- 6980 - 0x1b44  :   96 - 0x60
    "01100000", -- 6981 - 0x1b45  :   96 - 0x60
    "01111111", -- 6982 - 0x1b46  :  127 - 0x7f
    "00000000", -- 6983 - 0x1b47  :    0 - 0x0
    "01111111", -- 6984 - 0x1b48  :  127 - 0x7f
    "01100000", -- 6985 - 0x1b49  :   96 - 0x60
    "01100000", -- 6986 - 0x1b4a  :   96 - 0x60
    "01111110", -- 6987 - 0x1b4b  :  126 - 0x7e
    "01100000", -- 6988 - 0x1b4c  :   96 - 0x60
    "01100000", -- 6989 - 0x1b4d  :   96 - 0x60
    "01111111", -- 6990 - 0x1b4e  :  127 - 0x7f
    "00000000", -- 6991 - 0x1b4f  :    0 - 0x0
    "01111110", -- 6992 - 0x1b50  :  126 - 0x7e -- Background 0xb5
    "01100011", -- 6993 - 0x1b51  :   99 - 0x63
    "01100011", -- 6994 - 0x1b52  :   99 - 0x63
    "01100111", -- 6995 - 0x1b53  :  103 - 0x67
    "01111100", -- 6996 - 0x1b54  :  124 - 0x7c
    "01101110", -- 6997 - 0x1b55  :  110 - 0x6e
    "01100111", -- 6998 - 0x1b56  :  103 - 0x67
    "00000000", -- 6999 - 0x1b57  :    0 - 0x0
    "01111110", -- 7000 - 0x1b58  :  126 - 0x7e
    "01100011", -- 7001 - 0x1b59  :   99 - 0x63
    "01100011", -- 7002 - 0x1b5a  :   99 - 0x63
    "01100111", -- 7003 - 0x1b5b  :  103 - 0x67
    "01111100", -- 7004 - 0x1b5c  :  124 - 0x7c
    "01101110", -- 7005 - 0x1b5d  :  110 - 0x6e
    "01100111", -- 7006 - 0x1b5e  :  103 - 0x67
    "00000000", -- 7007 - 0x1b5f  :    0 - 0x0
    "00111110", -- 7008 - 0x1b60  :   62 - 0x3e -- Background 0xb6
    "01100011", -- 7009 - 0x1b61  :   99 - 0x63
    "01100011", -- 7010 - 0x1b62  :   99 - 0x63
    "01100011", -- 7011 - 0x1b63  :   99 - 0x63
    "01100011", -- 7012 - 0x1b64  :   99 - 0x63
    "01100011", -- 7013 - 0x1b65  :   99 - 0x63
    "00111110", -- 7014 - 0x1b66  :   62 - 0x3e
    "00000000", -- 7015 - 0x1b67  :    0 - 0x0
    "00111110", -- 7016 - 0x1b68  :   62 - 0x3e
    "01100011", -- 7017 - 0x1b69  :   99 - 0x63
    "01100011", -- 7018 - 0x1b6a  :   99 - 0x63
    "01100011", -- 7019 - 0x1b6b  :   99 - 0x63
    "01100011", -- 7020 - 0x1b6c  :   99 - 0x63
    "01100011", -- 7021 - 0x1b6d  :   99 - 0x63
    "00111110", -- 7022 - 0x1b6e  :   62 - 0x3e
    "00000000", -- 7023 - 0x1b6f  :    0 - 0x0
    "01100011", -- 7024 - 0x1b70  :   99 - 0x63 -- Background 0xb7
    "01110011", -- 7025 - 0x1b71  :  115 - 0x73
    "01111011", -- 7026 - 0x1b72  :  123 - 0x7b
    "01111111", -- 7027 - 0x1b73  :  127 - 0x7f
    "01101111", -- 7028 - 0x1b74  :  111 - 0x6f
    "01100111", -- 7029 - 0x1b75  :  103 - 0x67
    "01100011", -- 7030 - 0x1b76  :   99 - 0x63
    "00000000", -- 7031 - 0x1b77  :    0 - 0x0
    "01100011", -- 7032 - 0x1b78  :   99 - 0x63
    "01110011", -- 7033 - 0x1b79  :  115 - 0x73
    "01111011", -- 7034 - 0x1b7a  :  123 - 0x7b
    "01111111", -- 7035 - 0x1b7b  :  127 - 0x7f
    "01101111", -- 7036 - 0x1b7c  :  111 - 0x6f
    "01100111", -- 7037 - 0x1b7d  :  103 - 0x67
    "01100011", -- 7038 - 0x1b7e  :   99 - 0x63
    "00000000", -- 7039 - 0x1b7f  :    0 - 0x0
    "00111111", -- 7040 - 0x1b80  :   63 - 0x3f -- Background 0xb8
    "00001100", -- 7041 - 0x1b81  :   12 - 0xc
    "00001100", -- 7042 - 0x1b82  :   12 - 0xc
    "00001100", -- 7043 - 0x1b83  :   12 - 0xc
    "00001100", -- 7044 - 0x1b84  :   12 - 0xc
    "00001100", -- 7045 - 0x1b85  :   12 - 0xc
    "00001100", -- 7046 - 0x1b86  :   12 - 0xc
    "00000000", -- 7047 - 0x1b87  :    0 - 0x0
    "00111111", -- 7048 - 0x1b88  :   63 - 0x3f
    "00001100", -- 7049 - 0x1b89  :   12 - 0xc
    "00001100", -- 7050 - 0x1b8a  :   12 - 0xc
    "00001100", -- 7051 - 0x1b8b  :   12 - 0xc
    "00001100", -- 7052 - 0x1b8c  :   12 - 0xc
    "00001100", -- 7053 - 0x1b8d  :   12 - 0xc
    "00001100", -- 7054 - 0x1b8e  :   12 - 0xc
    "00000000", -- 7055 - 0x1b8f  :    0 - 0x0
    "01100011", -- 7056 - 0x1b90  :   99 - 0x63 -- Background 0xb9
    "01100011", -- 7057 - 0x1b91  :   99 - 0x63
    "01101011", -- 7058 - 0x1b92  :  107 - 0x6b
    "01111111", -- 7059 - 0x1b93  :  127 - 0x7f
    "01111111", -- 7060 - 0x1b94  :  127 - 0x7f
    "01110111", -- 7061 - 0x1b95  :  119 - 0x77
    "01100011", -- 7062 - 0x1b96  :   99 - 0x63
    "00000000", -- 7063 - 0x1b97  :    0 - 0x0
    "01100011", -- 7064 - 0x1b98  :   99 - 0x63
    "01100011", -- 7065 - 0x1b99  :   99 - 0x63
    "01101011", -- 7066 - 0x1b9a  :  107 - 0x6b
    "01111111", -- 7067 - 0x1b9b  :  127 - 0x7f
    "01111111", -- 7068 - 0x1b9c  :  127 - 0x7f
    "01110111", -- 7069 - 0x1b9d  :  119 - 0x77
    "01100011", -- 7070 - 0x1b9e  :   99 - 0x63
    "00000000", -- 7071 - 0x1b9f  :    0 - 0x0
    "01111100", -- 7072 - 0x1ba0  :  124 - 0x7c -- Background 0xba
    "01100110", -- 7073 - 0x1ba1  :  102 - 0x66
    "01100011", -- 7074 - 0x1ba2  :   99 - 0x63
    "01100011", -- 7075 - 0x1ba3  :   99 - 0x63
    "01100011", -- 7076 - 0x1ba4  :   99 - 0x63
    "01100110", -- 7077 - 0x1ba5  :  102 - 0x66
    "01111100", -- 7078 - 0x1ba6  :  124 - 0x7c
    "00000000", -- 7079 - 0x1ba7  :    0 - 0x0
    "00000000", -- 7080 - 0x1ba8  :    0 - 0x0
    "00000000", -- 7081 - 0x1ba9  :    0 - 0x0
    "00000000", -- 7082 - 0x1baa  :    0 - 0x0
    "00000000", -- 7083 - 0x1bab  :    0 - 0x0
    "00000000", -- 7084 - 0x1bac  :    0 - 0x0
    "00000000", -- 7085 - 0x1bad  :    0 - 0x0
    "00000000", -- 7086 - 0x1bae  :    0 - 0x0
    "00000000", -- 7087 - 0x1baf  :    0 - 0x0
    "00011100", -- 7088 - 0x1bb0  :   28 - 0x1c -- Background 0xbb
    "00011100", -- 7089 - 0x1bb1  :   28 - 0x1c
    "00011100", -- 7090 - 0x1bb2  :   28 - 0x1c
    "00011000", -- 7091 - 0x1bb3  :   24 - 0x18
    "00011000", -- 7092 - 0x1bb4  :   24 - 0x18
    "00000000", -- 7093 - 0x1bb5  :    0 - 0x0
    "00011000", -- 7094 - 0x1bb6  :   24 - 0x18
    "00000000", -- 7095 - 0x1bb7  :    0 - 0x0
    "00000000", -- 7096 - 0x1bb8  :    0 - 0x0
    "00000000", -- 7097 - 0x1bb9  :    0 - 0x0
    "00000000", -- 7098 - 0x1bba  :    0 - 0x0
    "00000000", -- 7099 - 0x1bbb  :    0 - 0x0
    "00000000", -- 7100 - 0x1bbc  :    0 - 0x0
    "00000000", -- 7101 - 0x1bbd  :    0 - 0x0
    "00000000", -- 7102 - 0x1bbe  :    0 - 0x0
    "00000000", -- 7103 - 0x1bbf  :    0 - 0x0
    "00011111", -- 7104 - 0x1bc0  :   31 - 0x1f -- Background 0xbc
    "00110000", -- 7105 - 0x1bc1  :   48 - 0x30
    "01100000", -- 7106 - 0x1bc2  :   96 - 0x60
    "01100111", -- 7107 - 0x1bc3  :  103 - 0x67
    "01100011", -- 7108 - 0x1bc4  :   99 - 0x63
    "00110011", -- 7109 - 0x1bc5  :   51 - 0x33
    "00011111", -- 7110 - 0x1bc6  :   31 - 0x1f
    "00000000", -- 7111 - 0x1bc7  :    0 - 0x0
    "00011111", -- 7112 - 0x1bc8  :   31 - 0x1f
    "00110000", -- 7113 - 0x1bc9  :   48 - 0x30
    "01100000", -- 7114 - 0x1bca  :   96 - 0x60
    "01100111", -- 7115 - 0x1bcb  :  103 - 0x67
    "01100011", -- 7116 - 0x1bcc  :   99 - 0x63
    "00110011", -- 7117 - 0x1bcd  :   51 - 0x33
    "00011111", -- 7118 - 0x1bce  :   31 - 0x1f
    "00000000", -- 7119 - 0x1bcf  :    0 - 0x0
    "01100011", -- 7120 - 0x1bd0  :   99 - 0x63 -- Background 0xbd
    "01110111", -- 7121 - 0x1bd1  :  119 - 0x77
    "01111111", -- 7122 - 0x1bd2  :  127 - 0x7f
    "01111111", -- 7123 - 0x1bd3  :  127 - 0x7f
    "01101011", -- 7124 - 0x1bd4  :  107 - 0x6b
    "01100011", -- 7125 - 0x1bd5  :   99 - 0x63
    "01100011", -- 7126 - 0x1bd6  :   99 - 0x63
    "00000000", -- 7127 - 0x1bd7  :    0 - 0x0
    "01100011", -- 7128 - 0x1bd8  :   99 - 0x63
    "01110111", -- 7129 - 0x1bd9  :  119 - 0x77
    "01111111", -- 7130 - 0x1bda  :  127 - 0x7f
    "01111111", -- 7131 - 0x1bdb  :  127 - 0x7f
    "01101011", -- 7132 - 0x1bdc  :  107 - 0x6b
    "01100011", -- 7133 - 0x1bdd  :   99 - 0x63
    "01100011", -- 7134 - 0x1bde  :   99 - 0x63
    "00000000", -- 7135 - 0x1bdf  :    0 - 0x0
    "01100011", -- 7136 - 0x1be0  :   99 - 0x63 -- Background 0xbe
    "01100011", -- 7137 - 0x1be1  :   99 - 0x63
    "01100011", -- 7138 - 0x1be2  :   99 - 0x63
    "01110111", -- 7139 - 0x1be3  :  119 - 0x77
    "00111110", -- 7140 - 0x1be4  :   62 - 0x3e
    "00011100", -- 7141 - 0x1be5  :   28 - 0x1c
    "00001000", -- 7142 - 0x1be6  :    8 - 0x8
    "00000000", -- 7143 - 0x1be7  :    0 - 0x0
    "01100011", -- 7144 - 0x1be8  :   99 - 0x63
    "01100011", -- 7145 - 0x1be9  :   99 - 0x63
    "01100011", -- 7146 - 0x1bea  :   99 - 0x63
    "01110111", -- 7147 - 0x1beb  :  119 - 0x77
    "00111110", -- 7148 - 0x1bec  :   62 - 0x3e
    "00011100", -- 7149 - 0x1bed  :   28 - 0x1c
    "00001000", -- 7150 - 0x1bee  :    8 - 0x8
    "00000000", -- 7151 - 0x1bef  :    0 - 0x0
    "00000000", -- 7152 - 0x1bf0  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 7153 - 0x1bf1  :    0 - 0x0
    "00000000", -- 7154 - 0x1bf2  :    0 - 0x0
    "00000000", -- 7155 - 0x1bf3  :    0 - 0x0
    "00000000", -- 7156 - 0x1bf4  :    0 - 0x0
    "00000000", -- 7157 - 0x1bf5  :    0 - 0x0
    "00000000", -- 7158 - 0x1bf6  :    0 - 0x0
    "00000000", -- 7159 - 0x1bf7  :    0 - 0x0
    "00000000", -- 7160 - 0x1bf8  :    0 - 0x0
    "00000000", -- 7161 - 0x1bf9  :    0 - 0x0
    "00000000", -- 7162 - 0x1bfa  :    0 - 0x0
    "00000000", -- 7163 - 0x1bfb  :    0 - 0x0
    "00000000", -- 7164 - 0x1bfc  :    0 - 0x0
    "00000000", -- 7165 - 0x1bfd  :    0 - 0x0
    "00000000", -- 7166 - 0x1bfe  :    0 - 0x0
    "00000000", -- 7167 - 0x1bff  :    0 - 0x0
    "00011111", -- 7168 - 0x1c00  :   31 - 0x1f -- Background 0xc0
    "00110000", -- 7169 - 0x1c01  :   48 - 0x30
    "01100000", -- 7170 - 0x1c02  :   96 - 0x60
    "01100111", -- 7171 - 0x1c03  :  103 - 0x67
    "01100011", -- 7172 - 0x1c04  :   99 - 0x63
    "00110011", -- 7173 - 0x1c05  :   51 - 0x33
    "00011111", -- 7174 - 0x1c06  :   31 - 0x1f
    "00000000", -- 7175 - 0x1c07  :    0 - 0x0
    "00000000", -- 7176 - 0x1c08  :    0 - 0x0
    "00000000", -- 7177 - 0x1c09  :    0 - 0x0
    "00000000", -- 7178 - 0x1c0a  :    0 - 0x0
    "00000000", -- 7179 - 0x1c0b  :    0 - 0x0
    "00000000", -- 7180 - 0x1c0c  :    0 - 0x0
    "00000000", -- 7181 - 0x1c0d  :    0 - 0x0
    "00000000", -- 7182 - 0x1c0e  :    0 - 0x0
    "00000000", -- 7183 - 0x1c0f  :    0 - 0x0
    "00011100", -- 7184 - 0x1c10  :   28 - 0x1c -- Background 0xc1
    "00110110", -- 7185 - 0x1c11  :   54 - 0x36
    "01100011", -- 7186 - 0x1c12  :   99 - 0x63
    "01100011", -- 7187 - 0x1c13  :   99 - 0x63
    "01111111", -- 7188 - 0x1c14  :  127 - 0x7f
    "01100011", -- 7189 - 0x1c15  :   99 - 0x63
    "01100011", -- 7190 - 0x1c16  :   99 - 0x63
    "00000000", -- 7191 - 0x1c17  :    0 - 0x0
    "00000000", -- 7192 - 0x1c18  :    0 - 0x0
    "00000000", -- 7193 - 0x1c19  :    0 - 0x0
    "00000000", -- 7194 - 0x1c1a  :    0 - 0x0
    "00000000", -- 7195 - 0x1c1b  :    0 - 0x0
    "00000000", -- 7196 - 0x1c1c  :    0 - 0x0
    "00000000", -- 7197 - 0x1c1d  :    0 - 0x0
    "00000000", -- 7198 - 0x1c1e  :    0 - 0x0
    "00000000", -- 7199 - 0x1c1f  :    0 - 0x0
    "01100011", -- 7200 - 0x1c20  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 7201 - 0x1c21  :  119 - 0x77
    "01111111", -- 7202 - 0x1c22  :  127 - 0x7f
    "01111111", -- 7203 - 0x1c23  :  127 - 0x7f
    "01101011", -- 7204 - 0x1c24  :  107 - 0x6b
    "01100011", -- 7205 - 0x1c25  :   99 - 0x63
    "01100011", -- 7206 - 0x1c26  :   99 - 0x63
    "00000000", -- 7207 - 0x1c27  :    0 - 0x0
    "00000000", -- 7208 - 0x1c28  :    0 - 0x0
    "00000000", -- 7209 - 0x1c29  :    0 - 0x0
    "00000000", -- 7210 - 0x1c2a  :    0 - 0x0
    "00000000", -- 7211 - 0x1c2b  :    0 - 0x0
    "00000000", -- 7212 - 0x1c2c  :    0 - 0x0
    "00000000", -- 7213 - 0x1c2d  :    0 - 0x0
    "00000000", -- 7214 - 0x1c2e  :    0 - 0x0
    "00000000", -- 7215 - 0x1c2f  :    0 - 0x0
    "01111111", -- 7216 - 0x1c30  :  127 - 0x7f -- Background 0xc3
    "01100000", -- 7217 - 0x1c31  :   96 - 0x60
    "01100000", -- 7218 - 0x1c32  :   96 - 0x60
    "01111110", -- 7219 - 0x1c33  :  126 - 0x7e
    "01100000", -- 7220 - 0x1c34  :   96 - 0x60
    "01100000", -- 7221 - 0x1c35  :   96 - 0x60
    "01111111", -- 7222 - 0x1c36  :  127 - 0x7f
    "00000000", -- 7223 - 0x1c37  :    0 - 0x0
    "00000000", -- 7224 - 0x1c38  :    0 - 0x0
    "00000000", -- 7225 - 0x1c39  :    0 - 0x0
    "00000000", -- 7226 - 0x1c3a  :    0 - 0x0
    "00000000", -- 7227 - 0x1c3b  :    0 - 0x0
    "00000000", -- 7228 - 0x1c3c  :    0 - 0x0
    "00000000", -- 7229 - 0x1c3d  :    0 - 0x0
    "00000000", -- 7230 - 0x1c3e  :    0 - 0x0
    "00000000", -- 7231 - 0x1c3f  :    0 - 0x0
    "00111110", -- 7232 - 0x1c40  :   62 - 0x3e -- Background 0xc4
    "01100011", -- 7233 - 0x1c41  :   99 - 0x63
    "01100011", -- 7234 - 0x1c42  :   99 - 0x63
    "01100011", -- 7235 - 0x1c43  :   99 - 0x63
    "01100011", -- 7236 - 0x1c44  :   99 - 0x63
    "01100011", -- 7237 - 0x1c45  :   99 - 0x63
    "00111110", -- 7238 - 0x1c46  :   62 - 0x3e
    "00000000", -- 7239 - 0x1c47  :    0 - 0x0
    "00000000", -- 7240 - 0x1c48  :    0 - 0x0
    "00000000", -- 7241 - 0x1c49  :    0 - 0x0
    "00000000", -- 7242 - 0x1c4a  :    0 - 0x0
    "00000000", -- 7243 - 0x1c4b  :    0 - 0x0
    "00000000", -- 7244 - 0x1c4c  :    0 - 0x0
    "00000000", -- 7245 - 0x1c4d  :    0 - 0x0
    "00000000", -- 7246 - 0x1c4e  :    0 - 0x0
    "00000000", -- 7247 - 0x1c4f  :    0 - 0x0
    "01100011", -- 7248 - 0x1c50  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 7249 - 0x1c51  :   99 - 0x63
    "01100011", -- 7250 - 0x1c52  :   99 - 0x63
    "01110111", -- 7251 - 0x1c53  :  119 - 0x77
    "00111110", -- 7252 - 0x1c54  :   62 - 0x3e
    "00011100", -- 7253 - 0x1c55  :   28 - 0x1c
    "00001000", -- 7254 - 0x1c56  :    8 - 0x8
    "00000000", -- 7255 - 0x1c57  :    0 - 0x0
    "00000000", -- 7256 - 0x1c58  :    0 - 0x0
    "00000000", -- 7257 - 0x1c59  :    0 - 0x0
    "00000000", -- 7258 - 0x1c5a  :    0 - 0x0
    "00000000", -- 7259 - 0x1c5b  :    0 - 0x0
    "00000000", -- 7260 - 0x1c5c  :    0 - 0x0
    "00000000", -- 7261 - 0x1c5d  :    0 - 0x0
    "00000000", -- 7262 - 0x1c5e  :    0 - 0x0
    "00000000", -- 7263 - 0x1c5f  :    0 - 0x0
    "01111110", -- 7264 - 0x1c60  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 7265 - 0x1c61  :   99 - 0x63
    "01100011", -- 7266 - 0x1c62  :   99 - 0x63
    "01100111", -- 7267 - 0x1c63  :  103 - 0x67
    "01111100", -- 7268 - 0x1c64  :  124 - 0x7c
    "01101110", -- 7269 - 0x1c65  :  110 - 0x6e
    "01100111", -- 7270 - 0x1c66  :  103 - 0x67
    "00000000", -- 7271 - 0x1c67  :    0 - 0x0
    "00000000", -- 7272 - 0x1c68  :    0 - 0x0
    "00000000", -- 7273 - 0x1c69  :    0 - 0x0
    "00000000", -- 7274 - 0x1c6a  :    0 - 0x0
    "00000000", -- 7275 - 0x1c6b  :    0 - 0x0
    "00000000", -- 7276 - 0x1c6c  :    0 - 0x0
    "00000000", -- 7277 - 0x1c6d  :    0 - 0x0
    "00000000", -- 7278 - 0x1c6e  :    0 - 0x0
    "00000000", -- 7279 - 0x1c6f  :    0 - 0x0
    "00110011", -- 7280 - 0x1c70  :   51 - 0x33 -- Background 0xc7
    "00110011", -- 7281 - 0x1c71  :   51 - 0x33
    "00110011", -- 7282 - 0x1c72  :   51 - 0x33
    "00011110", -- 7283 - 0x1c73  :   30 - 0x1e
    "00001100", -- 7284 - 0x1c74  :   12 - 0xc
    "00001100", -- 7285 - 0x1c75  :   12 - 0xc
    "00001100", -- 7286 - 0x1c76  :   12 - 0xc
    "00000000", -- 7287 - 0x1c77  :    0 - 0x0
    "00000000", -- 7288 - 0x1c78  :    0 - 0x0
    "00000000", -- 7289 - 0x1c79  :    0 - 0x0
    "00000000", -- 7290 - 0x1c7a  :    0 - 0x0
    "00000000", -- 7291 - 0x1c7b  :    0 - 0x0
    "00000000", -- 7292 - 0x1c7c  :    0 - 0x0
    "00000000", -- 7293 - 0x1c7d  :    0 - 0x0
    "00000000", -- 7294 - 0x1c7e  :    0 - 0x0
    "00000000", -- 7295 - 0x1c7f  :    0 - 0x0
    "00000000", -- 7296 - 0x1c80  :    0 - 0x0 -- Background 0xc8
    "00000000", -- 7297 - 0x1c81  :    0 - 0x0
    "00000000", -- 7298 - 0x1c82  :    0 - 0x0
    "00000000", -- 7299 - 0x1c83  :    0 - 0x0
    "00000000", -- 7300 - 0x1c84  :    0 - 0x0
    "00000000", -- 7301 - 0x1c85  :    0 - 0x0
    "00000000", -- 7302 - 0x1c86  :    0 - 0x0
    "00000000", -- 7303 - 0x1c87  :    0 - 0x0
    "00000000", -- 7304 - 0x1c88  :    0 - 0x0
    "00000000", -- 7305 - 0x1c89  :    0 - 0x0
    "00000000", -- 7306 - 0x1c8a  :    0 - 0x0
    "00000000", -- 7307 - 0x1c8b  :    0 - 0x0
    "00000000", -- 7308 - 0x1c8c  :    0 - 0x0
    "00000000", -- 7309 - 0x1c8d  :    0 - 0x0
    "00000000", -- 7310 - 0x1c8e  :    0 - 0x0
    "00000000", -- 7311 - 0x1c8f  :    0 - 0x0
    "00000000", -- 7312 - 0x1c90  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 7313 - 0x1c91  :    0 - 0x0
    "00000000", -- 7314 - 0x1c92  :    0 - 0x0
    "00000000", -- 7315 - 0x1c93  :    0 - 0x0
    "00000000", -- 7316 - 0x1c94  :    0 - 0x0
    "00000000", -- 7317 - 0x1c95  :    0 - 0x0
    "00000000", -- 7318 - 0x1c96  :    0 - 0x0
    "00000000", -- 7319 - 0x1c97  :    0 - 0x0
    "00000000", -- 7320 - 0x1c98  :    0 - 0x0
    "00000000", -- 7321 - 0x1c99  :    0 - 0x0
    "00000000", -- 7322 - 0x1c9a  :    0 - 0x0
    "00000000", -- 7323 - 0x1c9b  :    0 - 0x0
    "00000000", -- 7324 - 0x1c9c  :    0 - 0x0
    "00000000", -- 7325 - 0x1c9d  :    0 - 0x0
    "00000000", -- 7326 - 0x1c9e  :    0 - 0x0
    "00000000", -- 7327 - 0x1c9f  :    0 - 0x0
    "00000000", -- 7328 - 0x1ca0  :    0 - 0x0 -- Background 0xca
    "00000000", -- 7329 - 0x1ca1  :    0 - 0x0
    "00000000", -- 7330 - 0x1ca2  :    0 - 0x0
    "00000000", -- 7331 - 0x1ca3  :    0 - 0x0
    "00000000", -- 7332 - 0x1ca4  :    0 - 0x0
    "00000000", -- 7333 - 0x1ca5  :    0 - 0x0
    "00000000", -- 7334 - 0x1ca6  :    0 - 0x0
    "00000000", -- 7335 - 0x1ca7  :    0 - 0x0
    "00000000", -- 7336 - 0x1ca8  :    0 - 0x0
    "00000000", -- 7337 - 0x1ca9  :    0 - 0x0
    "00000000", -- 7338 - 0x1caa  :    0 - 0x0
    "00000000", -- 7339 - 0x1cab  :    0 - 0x0
    "00000000", -- 7340 - 0x1cac  :    0 - 0x0
    "00000000", -- 7341 - 0x1cad  :    0 - 0x0
    "00000000", -- 7342 - 0x1cae  :    0 - 0x0
    "00000000", -- 7343 - 0x1caf  :    0 - 0x0
    "00000000", -- 7344 - 0x1cb0  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 7345 - 0x1cb1  :    0 - 0x0
    "00000000", -- 7346 - 0x1cb2  :    0 - 0x0
    "00000000", -- 7347 - 0x1cb3  :    0 - 0x0
    "00000000", -- 7348 - 0x1cb4  :    0 - 0x0
    "00000000", -- 7349 - 0x1cb5  :    0 - 0x0
    "00000000", -- 7350 - 0x1cb6  :    0 - 0x0
    "00000000", -- 7351 - 0x1cb7  :    0 - 0x0
    "00000000", -- 7352 - 0x1cb8  :    0 - 0x0
    "00000000", -- 7353 - 0x1cb9  :    0 - 0x0
    "00000000", -- 7354 - 0x1cba  :    0 - 0x0
    "00000000", -- 7355 - 0x1cbb  :    0 - 0x0
    "00000000", -- 7356 - 0x1cbc  :    0 - 0x0
    "00000000", -- 7357 - 0x1cbd  :    0 - 0x0
    "00000000", -- 7358 - 0x1cbe  :    0 - 0x0
    "00000000", -- 7359 - 0x1cbf  :    0 - 0x0
    "00000000", -- 7360 - 0x1cc0  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 7361 - 0x1cc1  :    0 - 0x0
    "00000000", -- 7362 - 0x1cc2  :    0 - 0x0
    "00000000", -- 7363 - 0x1cc3  :    0 - 0x0
    "00000000", -- 7364 - 0x1cc4  :    0 - 0x0
    "00000000", -- 7365 - 0x1cc5  :    0 - 0x0
    "00000000", -- 7366 - 0x1cc6  :    0 - 0x0
    "00000000", -- 7367 - 0x1cc7  :    0 - 0x0
    "00000000", -- 7368 - 0x1cc8  :    0 - 0x0
    "00000000", -- 7369 - 0x1cc9  :    0 - 0x0
    "00000000", -- 7370 - 0x1cca  :    0 - 0x0
    "00000000", -- 7371 - 0x1ccb  :    0 - 0x0
    "00000000", -- 7372 - 0x1ccc  :    0 - 0x0
    "00000000", -- 7373 - 0x1ccd  :    0 - 0x0
    "00000000", -- 7374 - 0x1cce  :    0 - 0x0
    "00000000", -- 7375 - 0x1ccf  :    0 - 0x0
    "00000000", -- 7376 - 0x1cd0  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 7377 - 0x1cd1  :    0 - 0x0
    "00000000", -- 7378 - 0x1cd2  :    0 - 0x0
    "00000000", -- 7379 - 0x1cd3  :    0 - 0x0
    "00000000", -- 7380 - 0x1cd4  :    0 - 0x0
    "00000000", -- 7381 - 0x1cd5  :    0 - 0x0
    "00000000", -- 7382 - 0x1cd6  :    0 - 0x0
    "00000000", -- 7383 - 0x1cd7  :    0 - 0x0
    "00000000", -- 7384 - 0x1cd8  :    0 - 0x0
    "00000000", -- 7385 - 0x1cd9  :    0 - 0x0
    "00000000", -- 7386 - 0x1cda  :    0 - 0x0
    "00000000", -- 7387 - 0x1cdb  :    0 - 0x0
    "00000000", -- 7388 - 0x1cdc  :    0 - 0x0
    "00000000", -- 7389 - 0x1cdd  :    0 - 0x0
    "00000000", -- 7390 - 0x1cde  :    0 - 0x0
    "00000000", -- 7391 - 0x1cdf  :    0 - 0x0
    "00000000", -- 7392 - 0x1ce0  :    0 - 0x0 -- Background 0xce
    "00000000", -- 7393 - 0x1ce1  :    0 - 0x0
    "00000000", -- 7394 - 0x1ce2  :    0 - 0x0
    "00000000", -- 7395 - 0x1ce3  :    0 - 0x0
    "00000000", -- 7396 - 0x1ce4  :    0 - 0x0
    "00000000", -- 7397 - 0x1ce5  :    0 - 0x0
    "00000000", -- 7398 - 0x1ce6  :    0 - 0x0
    "00000000", -- 7399 - 0x1ce7  :    0 - 0x0
    "00000000", -- 7400 - 0x1ce8  :    0 - 0x0
    "00000000", -- 7401 - 0x1ce9  :    0 - 0x0
    "00000000", -- 7402 - 0x1cea  :    0 - 0x0
    "00000000", -- 7403 - 0x1ceb  :    0 - 0x0
    "00000000", -- 7404 - 0x1cec  :    0 - 0x0
    "00000000", -- 7405 - 0x1ced  :    0 - 0x0
    "00000000", -- 7406 - 0x1cee  :    0 - 0x0
    "00000000", -- 7407 - 0x1cef  :    0 - 0x0
    "00000000", -- 7408 - 0x1cf0  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 7409 - 0x1cf1  :    0 - 0x0
    "00000000", -- 7410 - 0x1cf2  :    0 - 0x0
    "00000000", -- 7411 - 0x1cf3  :    0 - 0x0
    "00000000", -- 7412 - 0x1cf4  :    0 - 0x0
    "00000000", -- 7413 - 0x1cf5  :    0 - 0x0
    "00000000", -- 7414 - 0x1cf6  :    0 - 0x0
    "00000000", -- 7415 - 0x1cf7  :    0 - 0x0
    "00000000", -- 7416 - 0x1cf8  :    0 - 0x0
    "00000000", -- 7417 - 0x1cf9  :    0 - 0x0
    "00000000", -- 7418 - 0x1cfa  :    0 - 0x0
    "00000000", -- 7419 - 0x1cfb  :    0 - 0x0
    "00000000", -- 7420 - 0x1cfc  :    0 - 0x0
    "00000000", -- 7421 - 0x1cfd  :    0 - 0x0
    "00000000", -- 7422 - 0x1cfe  :    0 - 0x0
    "00000000", -- 7423 - 0x1cff  :    0 - 0x0
    "11111111", -- 7424 - 0x1d00  :  255 - 0xff -- Background 0xd0
    "11111111", -- 7425 - 0x1d01  :  255 - 0xff
    "11111111", -- 7426 - 0x1d02  :  255 - 0xff
    "11111111", -- 7427 - 0x1d03  :  255 - 0xff
    "11111111", -- 7428 - 0x1d04  :  255 - 0xff
    "11111111", -- 7429 - 0x1d05  :  255 - 0xff
    "11111111", -- 7430 - 0x1d06  :  255 - 0xff
    "11111111", -- 7431 - 0x1d07  :  255 - 0xff
    "11111111", -- 7432 - 0x1d08  :  255 - 0xff
    "11111111", -- 7433 - 0x1d09  :  255 - 0xff
    "11111111", -- 7434 - 0x1d0a  :  255 - 0xff
    "11111111", -- 7435 - 0x1d0b  :  255 - 0xff
    "11111111", -- 7436 - 0x1d0c  :  255 - 0xff
    "11111111", -- 7437 - 0x1d0d  :  255 - 0xff
    "11111111", -- 7438 - 0x1d0e  :  255 - 0xff
    "11111111", -- 7439 - 0x1d0f  :  255 - 0xff
    "11111111", -- 7440 - 0x1d10  :  255 - 0xff -- Background 0xd1
    "11111111", -- 7441 - 0x1d11  :  255 - 0xff
    "11111111", -- 7442 - 0x1d12  :  255 - 0xff
    "11111111", -- 7443 - 0x1d13  :  255 - 0xff
    "11111111", -- 7444 - 0x1d14  :  255 - 0xff
    "11111111", -- 7445 - 0x1d15  :  255 - 0xff
    "11111111", -- 7446 - 0x1d16  :  255 - 0xff
    "11111111", -- 7447 - 0x1d17  :  255 - 0xff
    "11111111", -- 7448 - 0x1d18  :  255 - 0xff
    "11111111", -- 7449 - 0x1d19  :  255 - 0xff
    "11111111", -- 7450 - 0x1d1a  :  255 - 0xff
    "11111111", -- 7451 - 0x1d1b  :  255 - 0xff
    "11111111", -- 7452 - 0x1d1c  :  255 - 0xff
    "11111111", -- 7453 - 0x1d1d  :  255 - 0xff
    "11111111", -- 7454 - 0x1d1e  :  255 - 0xff
    "11111111", -- 7455 - 0x1d1f  :  255 - 0xff
    "11111111", -- 7456 - 0x1d20  :  255 - 0xff -- Background 0xd2
    "11111111", -- 7457 - 0x1d21  :  255 - 0xff
    "11111111", -- 7458 - 0x1d22  :  255 - 0xff
    "11111111", -- 7459 - 0x1d23  :  255 - 0xff
    "11111111", -- 7460 - 0x1d24  :  255 - 0xff
    "11111111", -- 7461 - 0x1d25  :  255 - 0xff
    "11111111", -- 7462 - 0x1d26  :  255 - 0xff
    "11111111", -- 7463 - 0x1d27  :  255 - 0xff
    "11111111", -- 7464 - 0x1d28  :  255 - 0xff
    "11111111", -- 7465 - 0x1d29  :  255 - 0xff
    "11111111", -- 7466 - 0x1d2a  :  255 - 0xff
    "11111111", -- 7467 - 0x1d2b  :  255 - 0xff
    "11111111", -- 7468 - 0x1d2c  :  255 - 0xff
    "11111111", -- 7469 - 0x1d2d  :  255 - 0xff
    "11111111", -- 7470 - 0x1d2e  :  255 - 0xff
    "11111111", -- 7471 - 0x1d2f  :  255 - 0xff
    "11111111", -- 7472 - 0x1d30  :  255 - 0xff -- Background 0xd3
    "11111111", -- 7473 - 0x1d31  :  255 - 0xff
    "11111111", -- 7474 - 0x1d32  :  255 - 0xff
    "11111111", -- 7475 - 0x1d33  :  255 - 0xff
    "11111111", -- 7476 - 0x1d34  :  255 - 0xff
    "11111111", -- 7477 - 0x1d35  :  255 - 0xff
    "11111111", -- 7478 - 0x1d36  :  255 - 0xff
    "11111111", -- 7479 - 0x1d37  :  255 - 0xff
    "11111111", -- 7480 - 0x1d38  :  255 - 0xff
    "11111111", -- 7481 - 0x1d39  :  255 - 0xff
    "11111111", -- 7482 - 0x1d3a  :  255 - 0xff
    "11111111", -- 7483 - 0x1d3b  :  255 - 0xff
    "11111111", -- 7484 - 0x1d3c  :  255 - 0xff
    "11111111", -- 7485 - 0x1d3d  :  255 - 0xff
    "11111111", -- 7486 - 0x1d3e  :  255 - 0xff
    "11111111", -- 7487 - 0x1d3f  :  255 - 0xff
    "11111111", -- 7488 - 0x1d40  :  255 - 0xff -- Background 0xd4
    "11111111", -- 7489 - 0x1d41  :  255 - 0xff
    "11111111", -- 7490 - 0x1d42  :  255 - 0xff
    "11111111", -- 7491 - 0x1d43  :  255 - 0xff
    "11111111", -- 7492 - 0x1d44  :  255 - 0xff
    "11111111", -- 7493 - 0x1d45  :  255 - 0xff
    "11111111", -- 7494 - 0x1d46  :  255 - 0xff
    "11111111", -- 7495 - 0x1d47  :  255 - 0xff
    "11111111", -- 7496 - 0x1d48  :  255 - 0xff
    "11111111", -- 7497 - 0x1d49  :  255 - 0xff
    "11111111", -- 7498 - 0x1d4a  :  255 - 0xff
    "11111111", -- 7499 - 0x1d4b  :  255 - 0xff
    "11111111", -- 7500 - 0x1d4c  :  255 - 0xff
    "11111111", -- 7501 - 0x1d4d  :  255 - 0xff
    "11111111", -- 7502 - 0x1d4e  :  255 - 0xff
    "11111111", -- 7503 - 0x1d4f  :  255 - 0xff
    "11111111", -- 7504 - 0x1d50  :  255 - 0xff -- Background 0xd5
    "11111111", -- 7505 - 0x1d51  :  255 - 0xff
    "11111111", -- 7506 - 0x1d52  :  255 - 0xff
    "11111111", -- 7507 - 0x1d53  :  255 - 0xff
    "11111111", -- 7508 - 0x1d54  :  255 - 0xff
    "11111111", -- 7509 - 0x1d55  :  255 - 0xff
    "11111111", -- 7510 - 0x1d56  :  255 - 0xff
    "11111111", -- 7511 - 0x1d57  :  255 - 0xff
    "11111111", -- 7512 - 0x1d58  :  255 - 0xff
    "11111111", -- 7513 - 0x1d59  :  255 - 0xff
    "11111111", -- 7514 - 0x1d5a  :  255 - 0xff
    "11111111", -- 7515 - 0x1d5b  :  255 - 0xff
    "11111111", -- 7516 - 0x1d5c  :  255 - 0xff
    "11111111", -- 7517 - 0x1d5d  :  255 - 0xff
    "11111111", -- 7518 - 0x1d5e  :  255 - 0xff
    "11111111", -- 7519 - 0x1d5f  :  255 - 0xff
    "11111111", -- 7520 - 0x1d60  :  255 - 0xff -- Background 0xd6
    "11111111", -- 7521 - 0x1d61  :  255 - 0xff
    "11111111", -- 7522 - 0x1d62  :  255 - 0xff
    "11111111", -- 7523 - 0x1d63  :  255 - 0xff
    "11111111", -- 7524 - 0x1d64  :  255 - 0xff
    "11111111", -- 7525 - 0x1d65  :  255 - 0xff
    "11111111", -- 7526 - 0x1d66  :  255 - 0xff
    "11111111", -- 7527 - 0x1d67  :  255 - 0xff
    "11111111", -- 7528 - 0x1d68  :  255 - 0xff
    "11111111", -- 7529 - 0x1d69  :  255 - 0xff
    "11111111", -- 7530 - 0x1d6a  :  255 - 0xff
    "11111111", -- 7531 - 0x1d6b  :  255 - 0xff
    "11111111", -- 7532 - 0x1d6c  :  255 - 0xff
    "11111111", -- 7533 - 0x1d6d  :  255 - 0xff
    "11111111", -- 7534 - 0x1d6e  :  255 - 0xff
    "11111111", -- 7535 - 0x1d6f  :  255 - 0xff
    "11111111", -- 7536 - 0x1d70  :  255 - 0xff -- Background 0xd7
    "11111111", -- 7537 - 0x1d71  :  255 - 0xff
    "11111111", -- 7538 - 0x1d72  :  255 - 0xff
    "11111111", -- 7539 - 0x1d73  :  255 - 0xff
    "11111111", -- 7540 - 0x1d74  :  255 - 0xff
    "11111111", -- 7541 - 0x1d75  :  255 - 0xff
    "11111111", -- 7542 - 0x1d76  :  255 - 0xff
    "11111111", -- 7543 - 0x1d77  :  255 - 0xff
    "11111111", -- 7544 - 0x1d78  :  255 - 0xff
    "11111111", -- 7545 - 0x1d79  :  255 - 0xff
    "11111111", -- 7546 - 0x1d7a  :  255 - 0xff
    "11111111", -- 7547 - 0x1d7b  :  255 - 0xff
    "11111111", -- 7548 - 0x1d7c  :  255 - 0xff
    "11111111", -- 7549 - 0x1d7d  :  255 - 0xff
    "11111111", -- 7550 - 0x1d7e  :  255 - 0xff
    "11111111", -- 7551 - 0x1d7f  :  255 - 0xff
    "11111111", -- 7552 - 0x1d80  :  255 - 0xff -- Background 0xd8
    "11111111", -- 7553 - 0x1d81  :  255 - 0xff
    "11111111", -- 7554 - 0x1d82  :  255 - 0xff
    "11111111", -- 7555 - 0x1d83  :  255 - 0xff
    "11111111", -- 7556 - 0x1d84  :  255 - 0xff
    "11111111", -- 7557 - 0x1d85  :  255 - 0xff
    "11111111", -- 7558 - 0x1d86  :  255 - 0xff
    "11111111", -- 7559 - 0x1d87  :  255 - 0xff
    "11111111", -- 7560 - 0x1d88  :  255 - 0xff
    "11111111", -- 7561 - 0x1d89  :  255 - 0xff
    "11111111", -- 7562 - 0x1d8a  :  255 - 0xff
    "11111111", -- 7563 - 0x1d8b  :  255 - 0xff
    "11111111", -- 7564 - 0x1d8c  :  255 - 0xff
    "11111111", -- 7565 - 0x1d8d  :  255 - 0xff
    "11111111", -- 7566 - 0x1d8e  :  255 - 0xff
    "11111111", -- 7567 - 0x1d8f  :  255 - 0xff
    "11111111", -- 7568 - 0x1d90  :  255 - 0xff -- Background 0xd9
    "11111111", -- 7569 - 0x1d91  :  255 - 0xff
    "11111111", -- 7570 - 0x1d92  :  255 - 0xff
    "11111111", -- 7571 - 0x1d93  :  255 - 0xff
    "11111111", -- 7572 - 0x1d94  :  255 - 0xff
    "11111111", -- 7573 - 0x1d95  :  255 - 0xff
    "11111111", -- 7574 - 0x1d96  :  255 - 0xff
    "11111111", -- 7575 - 0x1d97  :  255 - 0xff
    "11111111", -- 7576 - 0x1d98  :  255 - 0xff
    "11111111", -- 7577 - 0x1d99  :  255 - 0xff
    "11111111", -- 7578 - 0x1d9a  :  255 - 0xff
    "11111111", -- 7579 - 0x1d9b  :  255 - 0xff
    "11111111", -- 7580 - 0x1d9c  :  255 - 0xff
    "11111111", -- 7581 - 0x1d9d  :  255 - 0xff
    "11111111", -- 7582 - 0x1d9e  :  255 - 0xff
    "11111111", -- 7583 - 0x1d9f  :  255 - 0xff
    "11111111", -- 7584 - 0x1da0  :  255 - 0xff -- Background 0xda
    "11111111", -- 7585 - 0x1da1  :  255 - 0xff
    "11111111", -- 7586 - 0x1da2  :  255 - 0xff
    "11111111", -- 7587 - 0x1da3  :  255 - 0xff
    "11111111", -- 7588 - 0x1da4  :  255 - 0xff
    "11111111", -- 7589 - 0x1da5  :  255 - 0xff
    "11111111", -- 7590 - 0x1da6  :  255 - 0xff
    "11111111", -- 7591 - 0x1da7  :  255 - 0xff
    "11111111", -- 7592 - 0x1da8  :  255 - 0xff
    "11111111", -- 7593 - 0x1da9  :  255 - 0xff
    "11111111", -- 7594 - 0x1daa  :  255 - 0xff
    "11111111", -- 7595 - 0x1dab  :  255 - 0xff
    "11111111", -- 7596 - 0x1dac  :  255 - 0xff
    "11111111", -- 7597 - 0x1dad  :  255 - 0xff
    "11111111", -- 7598 - 0x1dae  :  255 - 0xff
    "11111111", -- 7599 - 0x1daf  :  255 - 0xff
    "11111111", -- 7600 - 0x1db0  :  255 - 0xff -- Background 0xdb
    "11111111", -- 7601 - 0x1db1  :  255 - 0xff
    "11111111", -- 7602 - 0x1db2  :  255 - 0xff
    "11111111", -- 7603 - 0x1db3  :  255 - 0xff
    "11111111", -- 7604 - 0x1db4  :  255 - 0xff
    "11111111", -- 7605 - 0x1db5  :  255 - 0xff
    "11111111", -- 7606 - 0x1db6  :  255 - 0xff
    "11111111", -- 7607 - 0x1db7  :  255 - 0xff
    "11111111", -- 7608 - 0x1db8  :  255 - 0xff
    "11111111", -- 7609 - 0x1db9  :  255 - 0xff
    "11111111", -- 7610 - 0x1dba  :  255 - 0xff
    "11111111", -- 7611 - 0x1dbb  :  255 - 0xff
    "11111111", -- 7612 - 0x1dbc  :  255 - 0xff
    "11111111", -- 7613 - 0x1dbd  :  255 - 0xff
    "11111111", -- 7614 - 0x1dbe  :  255 - 0xff
    "11111111", -- 7615 - 0x1dbf  :  255 - 0xff
    "11111111", -- 7616 - 0x1dc0  :  255 - 0xff -- Background 0xdc
    "11111111", -- 7617 - 0x1dc1  :  255 - 0xff
    "11111111", -- 7618 - 0x1dc2  :  255 - 0xff
    "11111111", -- 7619 - 0x1dc3  :  255 - 0xff
    "11111111", -- 7620 - 0x1dc4  :  255 - 0xff
    "11111111", -- 7621 - 0x1dc5  :  255 - 0xff
    "11111111", -- 7622 - 0x1dc6  :  255 - 0xff
    "11111111", -- 7623 - 0x1dc7  :  255 - 0xff
    "11111111", -- 7624 - 0x1dc8  :  255 - 0xff
    "11111111", -- 7625 - 0x1dc9  :  255 - 0xff
    "11111111", -- 7626 - 0x1dca  :  255 - 0xff
    "11111111", -- 7627 - 0x1dcb  :  255 - 0xff
    "11111111", -- 7628 - 0x1dcc  :  255 - 0xff
    "11111111", -- 7629 - 0x1dcd  :  255 - 0xff
    "11111111", -- 7630 - 0x1dce  :  255 - 0xff
    "11111111", -- 7631 - 0x1dcf  :  255 - 0xff
    "11111111", -- 7632 - 0x1dd0  :  255 - 0xff -- Background 0xdd
    "11111111", -- 7633 - 0x1dd1  :  255 - 0xff
    "11111111", -- 7634 - 0x1dd2  :  255 - 0xff
    "11111111", -- 7635 - 0x1dd3  :  255 - 0xff
    "11111111", -- 7636 - 0x1dd4  :  255 - 0xff
    "11111111", -- 7637 - 0x1dd5  :  255 - 0xff
    "11111111", -- 7638 - 0x1dd6  :  255 - 0xff
    "11111111", -- 7639 - 0x1dd7  :  255 - 0xff
    "11111111", -- 7640 - 0x1dd8  :  255 - 0xff
    "11111111", -- 7641 - 0x1dd9  :  255 - 0xff
    "11111111", -- 7642 - 0x1dda  :  255 - 0xff
    "11111111", -- 7643 - 0x1ddb  :  255 - 0xff
    "11111111", -- 7644 - 0x1ddc  :  255 - 0xff
    "11111111", -- 7645 - 0x1ddd  :  255 - 0xff
    "11111111", -- 7646 - 0x1dde  :  255 - 0xff
    "11111111", -- 7647 - 0x1ddf  :  255 - 0xff
    "11111111", -- 7648 - 0x1de0  :  255 - 0xff -- Background 0xde
    "11111111", -- 7649 - 0x1de1  :  255 - 0xff
    "11111111", -- 7650 - 0x1de2  :  255 - 0xff
    "11111111", -- 7651 - 0x1de3  :  255 - 0xff
    "11111111", -- 7652 - 0x1de4  :  255 - 0xff
    "11111111", -- 7653 - 0x1de5  :  255 - 0xff
    "11111111", -- 7654 - 0x1de6  :  255 - 0xff
    "11111111", -- 7655 - 0x1de7  :  255 - 0xff
    "11111111", -- 7656 - 0x1de8  :  255 - 0xff
    "11111111", -- 7657 - 0x1de9  :  255 - 0xff
    "11111111", -- 7658 - 0x1dea  :  255 - 0xff
    "11111111", -- 7659 - 0x1deb  :  255 - 0xff
    "11111111", -- 7660 - 0x1dec  :  255 - 0xff
    "11111111", -- 7661 - 0x1ded  :  255 - 0xff
    "11111111", -- 7662 - 0x1dee  :  255 - 0xff
    "11111111", -- 7663 - 0x1def  :  255 - 0xff
    "11111111", -- 7664 - 0x1df0  :  255 - 0xff -- Background 0xdf
    "11111111", -- 7665 - 0x1df1  :  255 - 0xff
    "11111111", -- 7666 - 0x1df2  :  255 - 0xff
    "11111111", -- 7667 - 0x1df3  :  255 - 0xff
    "11111111", -- 7668 - 0x1df4  :  255 - 0xff
    "11111111", -- 7669 - 0x1df5  :  255 - 0xff
    "11111111", -- 7670 - 0x1df6  :  255 - 0xff
    "11111111", -- 7671 - 0x1df7  :  255 - 0xff
    "11111111", -- 7672 - 0x1df8  :  255 - 0xff
    "11111111", -- 7673 - 0x1df9  :  255 - 0xff
    "11111111", -- 7674 - 0x1dfa  :  255 - 0xff
    "11111111", -- 7675 - 0x1dfb  :  255 - 0xff
    "11111111", -- 7676 - 0x1dfc  :  255 - 0xff
    "11111111", -- 7677 - 0x1dfd  :  255 - 0xff
    "11111111", -- 7678 - 0x1dfe  :  255 - 0xff
    "11111111", -- 7679 - 0x1dff  :  255 - 0xff
    "11111111", -- 7680 - 0x1e00  :  255 - 0xff -- Background 0xe0
    "11111111", -- 7681 - 0x1e01  :  255 - 0xff
    "11111111", -- 7682 - 0x1e02  :  255 - 0xff
    "11111111", -- 7683 - 0x1e03  :  255 - 0xff
    "11111111", -- 7684 - 0x1e04  :  255 - 0xff
    "11111111", -- 7685 - 0x1e05  :  255 - 0xff
    "11111111", -- 7686 - 0x1e06  :  255 - 0xff
    "11111111", -- 7687 - 0x1e07  :  255 - 0xff
    "11111111", -- 7688 - 0x1e08  :  255 - 0xff
    "11111111", -- 7689 - 0x1e09  :  255 - 0xff
    "11111111", -- 7690 - 0x1e0a  :  255 - 0xff
    "11111111", -- 7691 - 0x1e0b  :  255 - 0xff
    "11111111", -- 7692 - 0x1e0c  :  255 - 0xff
    "11111111", -- 7693 - 0x1e0d  :  255 - 0xff
    "11111111", -- 7694 - 0x1e0e  :  255 - 0xff
    "11111111", -- 7695 - 0x1e0f  :  255 - 0xff
    "11111111", -- 7696 - 0x1e10  :  255 - 0xff -- Background 0xe1
    "11111111", -- 7697 - 0x1e11  :  255 - 0xff
    "11111111", -- 7698 - 0x1e12  :  255 - 0xff
    "11111111", -- 7699 - 0x1e13  :  255 - 0xff
    "11111111", -- 7700 - 0x1e14  :  255 - 0xff
    "11111111", -- 7701 - 0x1e15  :  255 - 0xff
    "11111111", -- 7702 - 0x1e16  :  255 - 0xff
    "11111111", -- 7703 - 0x1e17  :  255 - 0xff
    "11111111", -- 7704 - 0x1e18  :  255 - 0xff
    "11111111", -- 7705 - 0x1e19  :  255 - 0xff
    "11111111", -- 7706 - 0x1e1a  :  255 - 0xff
    "11111111", -- 7707 - 0x1e1b  :  255 - 0xff
    "11111111", -- 7708 - 0x1e1c  :  255 - 0xff
    "11111111", -- 7709 - 0x1e1d  :  255 - 0xff
    "11111111", -- 7710 - 0x1e1e  :  255 - 0xff
    "11111111", -- 7711 - 0x1e1f  :  255 - 0xff
    "11111111", -- 7712 - 0x1e20  :  255 - 0xff -- Background 0xe2
    "11111111", -- 7713 - 0x1e21  :  255 - 0xff
    "11111111", -- 7714 - 0x1e22  :  255 - 0xff
    "11111111", -- 7715 - 0x1e23  :  255 - 0xff
    "11111111", -- 7716 - 0x1e24  :  255 - 0xff
    "11111111", -- 7717 - 0x1e25  :  255 - 0xff
    "11111111", -- 7718 - 0x1e26  :  255 - 0xff
    "11111111", -- 7719 - 0x1e27  :  255 - 0xff
    "11111111", -- 7720 - 0x1e28  :  255 - 0xff
    "11111111", -- 7721 - 0x1e29  :  255 - 0xff
    "11111111", -- 7722 - 0x1e2a  :  255 - 0xff
    "11111111", -- 7723 - 0x1e2b  :  255 - 0xff
    "11111111", -- 7724 - 0x1e2c  :  255 - 0xff
    "11111111", -- 7725 - 0x1e2d  :  255 - 0xff
    "11111111", -- 7726 - 0x1e2e  :  255 - 0xff
    "11111111", -- 7727 - 0x1e2f  :  255 - 0xff
    "11111111", -- 7728 - 0x1e30  :  255 - 0xff -- Background 0xe3
    "11111111", -- 7729 - 0x1e31  :  255 - 0xff
    "11111111", -- 7730 - 0x1e32  :  255 - 0xff
    "11111111", -- 7731 - 0x1e33  :  255 - 0xff
    "11111111", -- 7732 - 0x1e34  :  255 - 0xff
    "11111111", -- 7733 - 0x1e35  :  255 - 0xff
    "11111111", -- 7734 - 0x1e36  :  255 - 0xff
    "11111111", -- 7735 - 0x1e37  :  255 - 0xff
    "11111111", -- 7736 - 0x1e38  :  255 - 0xff
    "11111111", -- 7737 - 0x1e39  :  255 - 0xff
    "11111111", -- 7738 - 0x1e3a  :  255 - 0xff
    "11111111", -- 7739 - 0x1e3b  :  255 - 0xff
    "11111111", -- 7740 - 0x1e3c  :  255 - 0xff
    "11111111", -- 7741 - 0x1e3d  :  255 - 0xff
    "11111111", -- 7742 - 0x1e3e  :  255 - 0xff
    "11111111", -- 7743 - 0x1e3f  :  255 - 0xff
    "11111111", -- 7744 - 0x1e40  :  255 - 0xff -- Background 0xe4
    "11111111", -- 7745 - 0x1e41  :  255 - 0xff
    "11111111", -- 7746 - 0x1e42  :  255 - 0xff
    "11111111", -- 7747 - 0x1e43  :  255 - 0xff
    "11111111", -- 7748 - 0x1e44  :  255 - 0xff
    "11111111", -- 7749 - 0x1e45  :  255 - 0xff
    "11111111", -- 7750 - 0x1e46  :  255 - 0xff
    "11111111", -- 7751 - 0x1e47  :  255 - 0xff
    "11111111", -- 7752 - 0x1e48  :  255 - 0xff
    "11111111", -- 7753 - 0x1e49  :  255 - 0xff
    "11111111", -- 7754 - 0x1e4a  :  255 - 0xff
    "11111111", -- 7755 - 0x1e4b  :  255 - 0xff
    "11111111", -- 7756 - 0x1e4c  :  255 - 0xff
    "11111111", -- 7757 - 0x1e4d  :  255 - 0xff
    "11111111", -- 7758 - 0x1e4e  :  255 - 0xff
    "11111111", -- 7759 - 0x1e4f  :  255 - 0xff
    "11111111", -- 7760 - 0x1e50  :  255 - 0xff -- Background 0xe5
    "11111111", -- 7761 - 0x1e51  :  255 - 0xff
    "11111111", -- 7762 - 0x1e52  :  255 - 0xff
    "11111111", -- 7763 - 0x1e53  :  255 - 0xff
    "11111111", -- 7764 - 0x1e54  :  255 - 0xff
    "11111111", -- 7765 - 0x1e55  :  255 - 0xff
    "11111111", -- 7766 - 0x1e56  :  255 - 0xff
    "11111111", -- 7767 - 0x1e57  :  255 - 0xff
    "11111111", -- 7768 - 0x1e58  :  255 - 0xff
    "11111111", -- 7769 - 0x1e59  :  255 - 0xff
    "11111111", -- 7770 - 0x1e5a  :  255 - 0xff
    "11111111", -- 7771 - 0x1e5b  :  255 - 0xff
    "11111111", -- 7772 - 0x1e5c  :  255 - 0xff
    "11111111", -- 7773 - 0x1e5d  :  255 - 0xff
    "11111111", -- 7774 - 0x1e5e  :  255 - 0xff
    "11111111", -- 7775 - 0x1e5f  :  255 - 0xff
    "11111111", -- 7776 - 0x1e60  :  255 - 0xff -- Background 0xe6
    "11111111", -- 7777 - 0x1e61  :  255 - 0xff
    "11111111", -- 7778 - 0x1e62  :  255 - 0xff
    "11111111", -- 7779 - 0x1e63  :  255 - 0xff
    "11111111", -- 7780 - 0x1e64  :  255 - 0xff
    "11111111", -- 7781 - 0x1e65  :  255 - 0xff
    "11111111", -- 7782 - 0x1e66  :  255 - 0xff
    "11111111", -- 7783 - 0x1e67  :  255 - 0xff
    "11111111", -- 7784 - 0x1e68  :  255 - 0xff
    "11111111", -- 7785 - 0x1e69  :  255 - 0xff
    "11111111", -- 7786 - 0x1e6a  :  255 - 0xff
    "11111111", -- 7787 - 0x1e6b  :  255 - 0xff
    "11111111", -- 7788 - 0x1e6c  :  255 - 0xff
    "11111111", -- 7789 - 0x1e6d  :  255 - 0xff
    "11111111", -- 7790 - 0x1e6e  :  255 - 0xff
    "11111111", -- 7791 - 0x1e6f  :  255 - 0xff
    "11111111", -- 7792 - 0x1e70  :  255 - 0xff -- Background 0xe7
    "11111111", -- 7793 - 0x1e71  :  255 - 0xff
    "11111111", -- 7794 - 0x1e72  :  255 - 0xff
    "11111111", -- 7795 - 0x1e73  :  255 - 0xff
    "11111111", -- 7796 - 0x1e74  :  255 - 0xff
    "11111111", -- 7797 - 0x1e75  :  255 - 0xff
    "11111111", -- 7798 - 0x1e76  :  255 - 0xff
    "11111111", -- 7799 - 0x1e77  :  255 - 0xff
    "11111111", -- 7800 - 0x1e78  :  255 - 0xff
    "11111111", -- 7801 - 0x1e79  :  255 - 0xff
    "11111111", -- 7802 - 0x1e7a  :  255 - 0xff
    "11111111", -- 7803 - 0x1e7b  :  255 - 0xff
    "11111111", -- 7804 - 0x1e7c  :  255 - 0xff
    "11111111", -- 7805 - 0x1e7d  :  255 - 0xff
    "11111111", -- 7806 - 0x1e7e  :  255 - 0xff
    "11111111", -- 7807 - 0x1e7f  :  255 - 0xff
    "11111111", -- 7808 - 0x1e80  :  255 - 0xff -- Background 0xe8
    "11111111", -- 7809 - 0x1e81  :  255 - 0xff
    "11111111", -- 7810 - 0x1e82  :  255 - 0xff
    "11111111", -- 7811 - 0x1e83  :  255 - 0xff
    "11111111", -- 7812 - 0x1e84  :  255 - 0xff
    "11111111", -- 7813 - 0x1e85  :  255 - 0xff
    "11111111", -- 7814 - 0x1e86  :  255 - 0xff
    "11111111", -- 7815 - 0x1e87  :  255 - 0xff
    "11111111", -- 7816 - 0x1e88  :  255 - 0xff
    "11111111", -- 7817 - 0x1e89  :  255 - 0xff
    "11111111", -- 7818 - 0x1e8a  :  255 - 0xff
    "11111111", -- 7819 - 0x1e8b  :  255 - 0xff
    "11111111", -- 7820 - 0x1e8c  :  255 - 0xff
    "11111111", -- 7821 - 0x1e8d  :  255 - 0xff
    "11111111", -- 7822 - 0x1e8e  :  255 - 0xff
    "11111111", -- 7823 - 0x1e8f  :  255 - 0xff
    "11111111", -- 7824 - 0x1e90  :  255 - 0xff -- Background 0xe9
    "11111111", -- 7825 - 0x1e91  :  255 - 0xff
    "11111111", -- 7826 - 0x1e92  :  255 - 0xff
    "11111111", -- 7827 - 0x1e93  :  255 - 0xff
    "11111111", -- 7828 - 0x1e94  :  255 - 0xff
    "11111111", -- 7829 - 0x1e95  :  255 - 0xff
    "11111111", -- 7830 - 0x1e96  :  255 - 0xff
    "11111111", -- 7831 - 0x1e97  :  255 - 0xff
    "11111111", -- 7832 - 0x1e98  :  255 - 0xff
    "11111111", -- 7833 - 0x1e99  :  255 - 0xff
    "11111111", -- 7834 - 0x1e9a  :  255 - 0xff
    "11111111", -- 7835 - 0x1e9b  :  255 - 0xff
    "11111111", -- 7836 - 0x1e9c  :  255 - 0xff
    "11111111", -- 7837 - 0x1e9d  :  255 - 0xff
    "11111111", -- 7838 - 0x1e9e  :  255 - 0xff
    "11111111", -- 7839 - 0x1e9f  :  255 - 0xff
    "11111111", -- 7840 - 0x1ea0  :  255 - 0xff -- Background 0xea
    "11111111", -- 7841 - 0x1ea1  :  255 - 0xff
    "11111111", -- 7842 - 0x1ea2  :  255 - 0xff
    "11111111", -- 7843 - 0x1ea3  :  255 - 0xff
    "11111111", -- 7844 - 0x1ea4  :  255 - 0xff
    "11111111", -- 7845 - 0x1ea5  :  255 - 0xff
    "11111111", -- 7846 - 0x1ea6  :  255 - 0xff
    "11111111", -- 7847 - 0x1ea7  :  255 - 0xff
    "11111111", -- 7848 - 0x1ea8  :  255 - 0xff
    "11111111", -- 7849 - 0x1ea9  :  255 - 0xff
    "11111111", -- 7850 - 0x1eaa  :  255 - 0xff
    "11111111", -- 7851 - 0x1eab  :  255 - 0xff
    "11111111", -- 7852 - 0x1eac  :  255 - 0xff
    "11111111", -- 7853 - 0x1ead  :  255 - 0xff
    "11111111", -- 7854 - 0x1eae  :  255 - 0xff
    "11111111", -- 7855 - 0x1eaf  :  255 - 0xff
    "11111111", -- 7856 - 0x1eb0  :  255 - 0xff -- Background 0xeb
    "11111111", -- 7857 - 0x1eb1  :  255 - 0xff
    "11111111", -- 7858 - 0x1eb2  :  255 - 0xff
    "11111111", -- 7859 - 0x1eb3  :  255 - 0xff
    "11111111", -- 7860 - 0x1eb4  :  255 - 0xff
    "11111111", -- 7861 - 0x1eb5  :  255 - 0xff
    "11111111", -- 7862 - 0x1eb6  :  255 - 0xff
    "11111111", -- 7863 - 0x1eb7  :  255 - 0xff
    "11111111", -- 7864 - 0x1eb8  :  255 - 0xff
    "11111111", -- 7865 - 0x1eb9  :  255 - 0xff
    "11111111", -- 7866 - 0x1eba  :  255 - 0xff
    "11111111", -- 7867 - 0x1ebb  :  255 - 0xff
    "11111111", -- 7868 - 0x1ebc  :  255 - 0xff
    "11111111", -- 7869 - 0x1ebd  :  255 - 0xff
    "11111111", -- 7870 - 0x1ebe  :  255 - 0xff
    "11111111", -- 7871 - 0x1ebf  :  255 - 0xff
    "11111111", -- 7872 - 0x1ec0  :  255 - 0xff -- Background 0xec
    "11111111", -- 7873 - 0x1ec1  :  255 - 0xff
    "11111111", -- 7874 - 0x1ec2  :  255 - 0xff
    "11111111", -- 7875 - 0x1ec3  :  255 - 0xff
    "11111111", -- 7876 - 0x1ec4  :  255 - 0xff
    "11111111", -- 7877 - 0x1ec5  :  255 - 0xff
    "11111111", -- 7878 - 0x1ec6  :  255 - 0xff
    "11111111", -- 7879 - 0x1ec7  :  255 - 0xff
    "11111111", -- 7880 - 0x1ec8  :  255 - 0xff
    "11111111", -- 7881 - 0x1ec9  :  255 - 0xff
    "11111111", -- 7882 - 0x1eca  :  255 - 0xff
    "11111111", -- 7883 - 0x1ecb  :  255 - 0xff
    "11111111", -- 7884 - 0x1ecc  :  255 - 0xff
    "11111111", -- 7885 - 0x1ecd  :  255 - 0xff
    "11111111", -- 7886 - 0x1ece  :  255 - 0xff
    "11111111", -- 7887 - 0x1ecf  :  255 - 0xff
    "11111111", -- 7888 - 0x1ed0  :  255 - 0xff -- Background 0xed
    "11111111", -- 7889 - 0x1ed1  :  255 - 0xff
    "11111111", -- 7890 - 0x1ed2  :  255 - 0xff
    "11111111", -- 7891 - 0x1ed3  :  255 - 0xff
    "11111111", -- 7892 - 0x1ed4  :  255 - 0xff
    "11111111", -- 7893 - 0x1ed5  :  255 - 0xff
    "11111111", -- 7894 - 0x1ed6  :  255 - 0xff
    "11111111", -- 7895 - 0x1ed7  :  255 - 0xff
    "11111111", -- 7896 - 0x1ed8  :  255 - 0xff
    "11111111", -- 7897 - 0x1ed9  :  255 - 0xff
    "11111111", -- 7898 - 0x1eda  :  255 - 0xff
    "11111111", -- 7899 - 0x1edb  :  255 - 0xff
    "11111111", -- 7900 - 0x1edc  :  255 - 0xff
    "11111111", -- 7901 - 0x1edd  :  255 - 0xff
    "11111111", -- 7902 - 0x1ede  :  255 - 0xff
    "11111111", -- 7903 - 0x1edf  :  255 - 0xff
    "11111111", -- 7904 - 0x1ee0  :  255 - 0xff -- Background 0xee
    "11111111", -- 7905 - 0x1ee1  :  255 - 0xff
    "11111111", -- 7906 - 0x1ee2  :  255 - 0xff
    "11111111", -- 7907 - 0x1ee3  :  255 - 0xff
    "11111111", -- 7908 - 0x1ee4  :  255 - 0xff
    "11111111", -- 7909 - 0x1ee5  :  255 - 0xff
    "11111111", -- 7910 - 0x1ee6  :  255 - 0xff
    "11111111", -- 7911 - 0x1ee7  :  255 - 0xff
    "11111111", -- 7912 - 0x1ee8  :  255 - 0xff
    "11111111", -- 7913 - 0x1ee9  :  255 - 0xff
    "11111111", -- 7914 - 0x1eea  :  255 - 0xff
    "11111111", -- 7915 - 0x1eeb  :  255 - 0xff
    "11111111", -- 7916 - 0x1eec  :  255 - 0xff
    "11111111", -- 7917 - 0x1eed  :  255 - 0xff
    "11111111", -- 7918 - 0x1eee  :  255 - 0xff
    "11111111", -- 7919 - 0x1eef  :  255 - 0xff
    "11111111", -- 7920 - 0x1ef0  :  255 - 0xff -- Background 0xef
    "11111111", -- 7921 - 0x1ef1  :  255 - 0xff
    "11111111", -- 7922 - 0x1ef2  :  255 - 0xff
    "11111111", -- 7923 - 0x1ef3  :  255 - 0xff
    "11111111", -- 7924 - 0x1ef4  :  255 - 0xff
    "11111111", -- 7925 - 0x1ef5  :  255 - 0xff
    "11111111", -- 7926 - 0x1ef6  :  255 - 0xff
    "11111111", -- 7927 - 0x1ef7  :  255 - 0xff
    "11111111", -- 7928 - 0x1ef8  :  255 - 0xff
    "11111111", -- 7929 - 0x1ef9  :  255 - 0xff
    "11111111", -- 7930 - 0x1efa  :  255 - 0xff
    "11111111", -- 7931 - 0x1efb  :  255 - 0xff
    "11111111", -- 7932 - 0x1efc  :  255 - 0xff
    "11111111", -- 7933 - 0x1efd  :  255 - 0xff
    "11111111", -- 7934 - 0x1efe  :  255 - 0xff
    "11111111", -- 7935 - 0x1eff  :  255 - 0xff
    "11111111", -- 7936 - 0x1f00  :  255 - 0xff -- Background 0xf0
    "11111111", -- 7937 - 0x1f01  :  255 - 0xff
    "11111111", -- 7938 - 0x1f02  :  255 - 0xff
    "11111111", -- 7939 - 0x1f03  :  255 - 0xff
    "11111111", -- 7940 - 0x1f04  :  255 - 0xff
    "11111111", -- 7941 - 0x1f05  :  255 - 0xff
    "11111111", -- 7942 - 0x1f06  :  255 - 0xff
    "11111111", -- 7943 - 0x1f07  :  255 - 0xff
    "11111111", -- 7944 - 0x1f08  :  255 - 0xff
    "11111111", -- 7945 - 0x1f09  :  255 - 0xff
    "11111111", -- 7946 - 0x1f0a  :  255 - 0xff
    "11111111", -- 7947 - 0x1f0b  :  255 - 0xff
    "11111111", -- 7948 - 0x1f0c  :  255 - 0xff
    "11111111", -- 7949 - 0x1f0d  :  255 - 0xff
    "11111111", -- 7950 - 0x1f0e  :  255 - 0xff
    "11111111", -- 7951 - 0x1f0f  :  255 - 0xff
    "11111111", -- 7952 - 0x1f10  :  255 - 0xff -- Background 0xf1
    "11111111", -- 7953 - 0x1f11  :  255 - 0xff
    "11111111", -- 7954 - 0x1f12  :  255 - 0xff
    "11111111", -- 7955 - 0x1f13  :  255 - 0xff
    "11111111", -- 7956 - 0x1f14  :  255 - 0xff
    "11111111", -- 7957 - 0x1f15  :  255 - 0xff
    "11111111", -- 7958 - 0x1f16  :  255 - 0xff
    "11111111", -- 7959 - 0x1f17  :  255 - 0xff
    "11111111", -- 7960 - 0x1f18  :  255 - 0xff
    "11111111", -- 7961 - 0x1f19  :  255 - 0xff
    "11111111", -- 7962 - 0x1f1a  :  255 - 0xff
    "11111111", -- 7963 - 0x1f1b  :  255 - 0xff
    "11111111", -- 7964 - 0x1f1c  :  255 - 0xff
    "11111111", -- 7965 - 0x1f1d  :  255 - 0xff
    "11111111", -- 7966 - 0x1f1e  :  255 - 0xff
    "11111111", -- 7967 - 0x1f1f  :  255 - 0xff
    "11111111", -- 7968 - 0x1f20  :  255 - 0xff -- Background 0xf2
    "11111111", -- 7969 - 0x1f21  :  255 - 0xff
    "11111111", -- 7970 - 0x1f22  :  255 - 0xff
    "11111111", -- 7971 - 0x1f23  :  255 - 0xff
    "11111111", -- 7972 - 0x1f24  :  255 - 0xff
    "11111111", -- 7973 - 0x1f25  :  255 - 0xff
    "11111111", -- 7974 - 0x1f26  :  255 - 0xff
    "11111111", -- 7975 - 0x1f27  :  255 - 0xff
    "11111111", -- 7976 - 0x1f28  :  255 - 0xff
    "11111111", -- 7977 - 0x1f29  :  255 - 0xff
    "11111111", -- 7978 - 0x1f2a  :  255 - 0xff
    "11111111", -- 7979 - 0x1f2b  :  255 - 0xff
    "11111111", -- 7980 - 0x1f2c  :  255 - 0xff
    "11111111", -- 7981 - 0x1f2d  :  255 - 0xff
    "11111111", -- 7982 - 0x1f2e  :  255 - 0xff
    "11111111", -- 7983 - 0x1f2f  :  255 - 0xff
    "11111111", -- 7984 - 0x1f30  :  255 - 0xff -- Background 0xf3
    "11111111", -- 7985 - 0x1f31  :  255 - 0xff
    "11111111", -- 7986 - 0x1f32  :  255 - 0xff
    "11111111", -- 7987 - 0x1f33  :  255 - 0xff
    "11111111", -- 7988 - 0x1f34  :  255 - 0xff
    "11111111", -- 7989 - 0x1f35  :  255 - 0xff
    "11111111", -- 7990 - 0x1f36  :  255 - 0xff
    "11111111", -- 7991 - 0x1f37  :  255 - 0xff
    "11111111", -- 7992 - 0x1f38  :  255 - 0xff
    "11111111", -- 7993 - 0x1f39  :  255 - 0xff
    "11111111", -- 7994 - 0x1f3a  :  255 - 0xff
    "11111111", -- 7995 - 0x1f3b  :  255 - 0xff
    "11111111", -- 7996 - 0x1f3c  :  255 - 0xff
    "11111111", -- 7997 - 0x1f3d  :  255 - 0xff
    "11111111", -- 7998 - 0x1f3e  :  255 - 0xff
    "11111111", -- 7999 - 0x1f3f  :  255 - 0xff
    "11111111", -- 8000 - 0x1f40  :  255 - 0xff -- Background 0xf4
    "11111111", -- 8001 - 0x1f41  :  255 - 0xff
    "11111111", -- 8002 - 0x1f42  :  255 - 0xff
    "11111111", -- 8003 - 0x1f43  :  255 - 0xff
    "11111111", -- 8004 - 0x1f44  :  255 - 0xff
    "11111111", -- 8005 - 0x1f45  :  255 - 0xff
    "11111111", -- 8006 - 0x1f46  :  255 - 0xff
    "11111111", -- 8007 - 0x1f47  :  255 - 0xff
    "11111111", -- 8008 - 0x1f48  :  255 - 0xff
    "11111111", -- 8009 - 0x1f49  :  255 - 0xff
    "11111111", -- 8010 - 0x1f4a  :  255 - 0xff
    "11111111", -- 8011 - 0x1f4b  :  255 - 0xff
    "11111111", -- 8012 - 0x1f4c  :  255 - 0xff
    "11111111", -- 8013 - 0x1f4d  :  255 - 0xff
    "11111111", -- 8014 - 0x1f4e  :  255 - 0xff
    "11111111", -- 8015 - 0x1f4f  :  255 - 0xff
    "11111111", -- 8016 - 0x1f50  :  255 - 0xff -- Background 0xf5
    "11111111", -- 8017 - 0x1f51  :  255 - 0xff
    "11111111", -- 8018 - 0x1f52  :  255 - 0xff
    "11111111", -- 8019 - 0x1f53  :  255 - 0xff
    "11111111", -- 8020 - 0x1f54  :  255 - 0xff
    "11111111", -- 8021 - 0x1f55  :  255 - 0xff
    "11111111", -- 8022 - 0x1f56  :  255 - 0xff
    "11111111", -- 8023 - 0x1f57  :  255 - 0xff
    "11111111", -- 8024 - 0x1f58  :  255 - 0xff
    "11111111", -- 8025 - 0x1f59  :  255 - 0xff
    "11111111", -- 8026 - 0x1f5a  :  255 - 0xff
    "11111111", -- 8027 - 0x1f5b  :  255 - 0xff
    "11111111", -- 8028 - 0x1f5c  :  255 - 0xff
    "11111111", -- 8029 - 0x1f5d  :  255 - 0xff
    "11111111", -- 8030 - 0x1f5e  :  255 - 0xff
    "11111111", -- 8031 - 0x1f5f  :  255 - 0xff
    "11111111", -- 8032 - 0x1f60  :  255 - 0xff -- Background 0xf6
    "11111111", -- 8033 - 0x1f61  :  255 - 0xff
    "11111111", -- 8034 - 0x1f62  :  255 - 0xff
    "11111111", -- 8035 - 0x1f63  :  255 - 0xff
    "11111111", -- 8036 - 0x1f64  :  255 - 0xff
    "11111111", -- 8037 - 0x1f65  :  255 - 0xff
    "11111111", -- 8038 - 0x1f66  :  255 - 0xff
    "11111111", -- 8039 - 0x1f67  :  255 - 0xff
    "11111111", -- 8040 - 0x1f68  :  255 - 0xff
    "11111111", -- 8041 - 0x1f69  :  255 - 0xff
    "11111111", -- 8042 - 0x1f6a  :  255 - 0xff
    "11111111", -- 8043 - 0x1f6b  :  255 - 0xff
    "11111111", -- 8044 - 0x1f6c  :  255 - 0xff
    "11111111", -- 8045 - 0x1f6d  :  255 - 0xff
    "11111111", -- 8046 - 0x1f6e  :  255 - 0xff
    "11111111", -- 8047 - 0x1f6f  :  255 - 0xff
    "11111111", -- 8048 - 0x1f70  :  255 - 0xff -- Background 0xf7
    "11111111", -- 8049 - 0x1f71  :  255 - 0xff
    "11111111", -- 8050 - 0x1f72  :  255 - 0xff
    "11111111", -- 8051 - 0x1f73  :  255 - 0xff
    "11111111", -- 8052 - 0x1f74  :  255 - 0xff
    "11111111", -- 8053 - 0x1f75  :  255 - 0xff
    "11111111", -- 8054 - 0x1f76  :  255 - 0xff
    "11111111", -- 8055 - 0x1f77  :  255 - 0xff
    "11111111", -- 8056 - 0x1f78  :  255 - 0xff
    "11111111", -- 8057 - 0x1f79  :  255 - 0xff
    "11111111", -- 8058 - 0x1f7a  :  255 - 0xff
    "11111111", -- 8059 - 0x1f7b  :  255 - 0xff
    "11111111", -- 8060 - 0x1f7c  :  255 - 0xff
    "11111111", -- 8061 - 0x1f7d  :  255 - 0xff
    "11111111", -- 8062 - 0x1f7e  :  255 - 0xff
    "11111111", -- 8063 - 0x1f7f  :  255 - 0xff
    "11111111", -- 8064 - 0x1f80  :  255 - 0xff -- Background 0xf8
    "11111111", -- 8065 - 0x1f81  :  255 - 0xff
    "11111111", -- 8066 - 0x1f82  :  255 - 0xff
    "11111111", -- 8067 - 0x1f83  :  255 - 0xff
    "11111111", -- 8068 - 0x1f84  :  255 - 0xff
    "11111111", -- 8069 - 0x1f85  :  255 - 0xff
    "11111111", -- 8070 - 0x1f86  :  255 - 0xff
    "11111111", -- 8071 - 0x1f87  :  255 - 0xff
    "11111111", -- 8072 - 0x1f88  :  255 - 0xff
    "11111111", -- 8073 - 0x1f89  :  255 - 0xff
    "11111111", -- 8074 - 0x1f8a  :  255 - 0xff
    "11111111", -- 8075 - 0x1f8b  :  255 - 0xff
    "11111111", -- 8076 - 0x1f8c  :  255 - 0xff
    "11111111", -- 8077 - 0x1f8d  :  255 - 0xff
    "11111111", -- 8078 - 0x1f8e  :  255 - 0xff
    "11111111", -- 8079 - 0x1f8f  :  255 - 0xff
    "11111111", -- 8080 - 0x1f90  :  255 - 0xff -- Background 0xf9
    "11111111", -- 8081 - 0x1f91  :  255 - 0xff
    "11111111", -- 8082 - 0x1f92  :  255 - 0xff
    "11111111", -- 8083 - 0x1f93  :  255 - 0xff
    "11111111", -- 8084 - 0x1f94  :  255 - 0xff
    "11111111", -- 8085 - 0x1f95  :  255 - 0xff
    "11111111", -- 8086 - 0x1f96  :  255 - 0xff
    "11111111", -- 8087 - 0x1f97  :  255 - 0xff
    "11111111", -- 8088 - 0x1f98  :  255 - 0xff
    "11111111", -- 8089 - 0x1f99  :  255 - 0xff
    "11111111", -- 8090 - 0x1f9a  :  255 - 0xff
    "11111111", -- 8091 - 0x1f9b  :  255 - 0xff
    "11111111", -- 8092 - 0x1f9c  :  255 - 0xff
    "11111111", -- 8093 - 0x1f9d  :  255 - 0xff
    "11111111", -- 8094 - 0x1f9e  :  255 - 0xff
    "11111111", -- 8095 - 0x1f9f  :  255 - 0xff
    "11111111", -- 8096 - 0x1fa0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 8097 - 0x1fa1  :  255 - 0xff
    "11111111", -- 8098 - 0x1fa2  :  255 - 0xff
    "11111111", -- 8099 - 0x1fa3  :  255 - 0xff
    "11111111", -- 8100 - 0x1fa4  :  255 - 0xff
    "11111111", -- 8101 - 0x1fa5  :  255 - 0xff
    "11111111", -- 8102 - 0x1fa6  :  255 - 0xff
    "11111111", -- 8103 - 0x1fa7  :  255 - 0xff
    "11111111", -- 8104 - 0x1fa8  :  255 - 0xff
    "11111111", -- 8105 - 0x1fa9  :  255 - 0xff
    "11111111", -- 8106 - 0x1faa  :  255 - 0xff
    "11111111", -- 8107 - 0x1fab  :  255 - 0xff
    "11111111", -- 8108 - 0x1fac  :  255 - 0xff
    "11111111", -- 8109 - 0x1fad  :  255 - 0xff
    "11111111", -- 8110 - 0x1fae  :  255 - 0xff
    "11111111", -- 8111 - 0x1faf  :  255 - 0xff
    "11111111", -- 8112 - 0x1fb0  :  255 - 0xff -- Background 0xfb
    "11111111", -- 8113 - 0x1fb1  :  255 - 0xff
    "11111111", -- 8114 - 0x1fb2  :  255 - 0xff
    "11111111", -- 8115 - 0x1fb3  :  255 - 0xff
    "11111111", -- 8116 - 0x1fb4  :  255 - 0xff
    "11111111", -- 8117 - 0x1fb5  :  255 - 0xff
    "11111111", -- 8118 - 0x1fb6  :  255 - 0xff
    "11111111", -- 8119 - 0x1fb7  :  255 - 0xff
    "11111111", -- 8120 - 0x1fb8  :  255 - 0xff
    "11111111", -- 8121 - 0x1fb9  :  255 - 0xff
    "11111111", -- 8122 - 0x1fba  :  255 - 0xff
    "11111111", -- 8123 - 0x1fbb  :  255 - 0xff
    "11111111", -- 8124 - 0x1fbc  :  255 - 0xff
    "11111111", -- 8125 - 0x1fbd  :  255 - 0xff
    "11111111", -- 8126 - 0x1fbe  :  255 - 0xff
    "11111111", -- 8127 - 0x1fbf  :  255 - 0xff
    "11111111", -- 8128 - 0x1fc0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 8129 - 0x1fc1  :  255 - 0xff
    "11111111", -- 8130 - 0x1fc2  :  255 - 0xff
    "11111111", -- 8131 - 0x1fc3  :  255 - 0xff
    "11111111", -- 8132 - 0x1fc4  :  255 - 0xff
    "11111111", -- 8133 - 0x1fc5  :  255 - 0xff
    "11111111", -- 8134 - 0x1fc6  :  255 - 0xff
    "11111111", -- 8135 - 0x1fc7  :  255 - 0xff
    "11111111", -- 8136 - 0x1fc8  :  255 - 0xff
    "11111111", -- 8137 - 0x1fc9  :  255 - 0xff
    "11111111", -- 8138 - 0x1fca  :  255 - 0xff
    "11111111", -- 8139 - 0x1fcb  :  255 - 0xff
    "11111111", -- 8140 - 0x1fcc  :  255 - 0xff
    "11111111", -- 8141 - 0x1fcd  :  255 - 0xff
    "11111111", -- 8142 - 0x1fce  :  255 - 0xff
    "11111111", -- 8143 - 0x1fcf  :  255 - 0xff
    "11111111", -- 8144 - 0x1fd0  :  255 - 0xff -- Background 0xfd
    "11111111", -- 8145 - 0x1fd1  :  255 - 0xff
    "11111111", -- 8146 - 0x1fd2  :  255 - 0xff
    "11111111", -- 8147 - 0x1fd3  :  255 - 0xff
    "11111111", -- 8148 - 0x1fd4  :  255 - 0xff
    "11111111", -- 8149 - 0x1fd5  :  255 - 0xff
    "11111111", -- 8150 - 0x1fd6  :  255 - 0xff
    "11111111", -- 8151 - 0x1fd7  :  255 - 0xff
    "11111111", -- 8152 - 0x1fd8  :  255 - 0xff
    "11111111", -- 8153 - 0x1fd9  :  255 - 0xff
    "11111111", -- 8154 - 0x1fda  :  255 - 0xff
    "11111111", -- 8155 - 0x1fdb  :  255 - 0xff
    "11111111", -- 8156 - 0x1fdc  :  255 - 0xff
    "11111111", -- 8157 - 0x1fdd  :  255 - 0xff
    "11111111", -- 8158 - 0x1fde  :  255 - 0xff
    "11111111", -- 8159 - 0x1fdf  :  255 - 0xff
    "11111111", -- 8160 - 0x1fe0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 8161 - 0x1fe1  :  255 - 0xff
    "11111111", -- 8162 - 0x1fe2  :  255 - 0xff
    "11111111", -- 8163 - 0x1fe3  :  255 - 0xff
    "11111111", -- 8164 - 0x1fe4  :  255 - 0xff
    "11111111", -- 8165 - 0x1fe5  :  255 - 0xff
    "11111111", -- 8166 - 0x1fe6  :  255 - 0xff
    "11111111", -- 8167 - 0x1fe7  :  255 - 0xff
    "11111111", -- 8168 - 0x1fe8  :  255 - 0xff
    "11111111", -- 8169 - 0x1fe9  :  255 - 0xff
    "11111111", -- 8170 - 0x1fea  :  255 - 0xff
    "11111111", -- 8171 - 0x1feb  :  255 - 0xff
    "11111111", -- 8172 - 0x1fec  :  255 - 0xff
    "11111111", -- 8173 - 0x1fed  :  255 - 0xff
    "11111111", -- 8174 - 0x1fee  :  255 - 0xff
    "11111111", -- 8175 - 0x1fef  :  255 - 0xff
    "11111111", -- 8176 - 0x1ff0  :  255 - 0xff -- Background 0xff
    "11111111", -- 8177 - 0x1ff1  :  255 - 0xff
    "11111111", -- 8178 - 0x1ff2  :  255 - 0xff
    "11111111", -- 8179 - 0x1ff3  :  255 - 0xff
    "11111111", -- 8180 - 0x1ff4  :  255 - 0xff
    "11111111", -- 8181 - 0x1ff5  :  255 - 0xff
    "11111111", -- 8182 - 0x1ff6  :  255 - 0xff
    "11111111", -- 8183 - 0x1ff7  :  255 - 0xff
    "11111111", -- 8184 - 0x1ff8  :  255 - 0xff
    "11111111", -- 8185 - 0x1ff9  :  255 - 0xff
    "11111111", -- 8186 - 0x1ffa  :  255 - 0xff
    "11111111", -- 8187 - 0x1ffb  :  255 - 0xff
    "11111111", -- 8188 - 0x1ffc  :  255 - 0xff
    "11111111", -- 8189 - 0x1ffd  :  255 - 0xff
    "11111111", -- 8190 - 0x1ffe  :  255 - 0xff
    "11111111"  -- 8191 - 0x1fff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
