//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: nova_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE_NOVA_00
  (
     //input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout  = 8'b00110000; //    0 :  48 - 0x30 -- line 0x0
      10'h1: dout  = 8'b00111111; //    1 :  63 - 0x3f
      10'h2: dout  = 8'b00110000; //    2 :  48 - 0x30
      10'h3: dout  = 8'b00111111; //    3 :  63 - 0x3f
      10'h4: dout  = 8'b00110000; //    4 :  48 - 0x30
      10'h5: dout  = 8'b00111111; //    5 :  63 - 0x3f
      10'h6: dout  = 8'b00110000; //    6 :  48 - 0x30
      10'h7: dout  = 8'b00111111; //    7 :  63 - 0x3f
      10'h8: dout  = 8'b00110000; //    8 :  48 - 0x30
      10'h9: dout  = 8'b00111111; //    9 :  63 - 0x3f
      10'hA: dout  = 8'b00110000; //   10 :  48 - 0x30
      10'hB: dout  = 8'b00111111; //   11 :  63 - 0x3f
      10'hC: dout  = 8'b00110000; //   12 :  48 - 0x30
      10'hD: dout  = 8'b00111111; //   13 :  63 - 0x3f
      10'hE: dout  = 8'b00110000; //   14 :  48 - 0x30
      10'hF: dout  = 8'b00111111; //   15 :  63 - 0x3f
      10'h10: dout  = 8'b00110000; //   16 :  48 - 0x30
      10'h11: dout  = 8'b00111111; //   17 :  63 - 0x3f
      10'h12: dout  = 8'b00110000; //   18 :  48 - 0x30
      10'h13: dout  = 8'b00111111; //   19 :  63 - 0x3f
      10'h14: dout  = 8'b01110000; //   20 : 112 - 0x70
      10'h15: dout  = 8'b01110001; //   21 : 113 - 0x71
      10'h16: dout  = 8'b01110001; //   22 : 113 - 0x71
      10'h17: dout  = 8'b01110001; //   23 : 113 - 0x71
      10'h18: dout  = 8'b01110001; //   24 : 113 - 0x71
      10'h19: dout  = 8'b01110001; //   25 : 113 - 0x71
      10'h1A: dout  = 8'b01110001; //   26 : 113 - 0x71
      10'h1B: dout  = 8'b01110001; //   27 : 113 - 0x71
      10'h1C: dout  = 8'b01110001; //   28 : 113 - 0x71
      10'h1D: dout  = 8'b01110001; //   29 : 113 - 0x71
      10'h1E: dout  = 8'b01110001; //   30 : 113 - 0x71
      10'h1F: dout  = 8'b01110001; //   31 : 113 - 0x71
      10'h20: dout  = 8'b00111111; //   32 :  63 - 0x3f -- line 0x1
      10'h21: dout  = 8'b00110000; //   33 :  48 - 0x30
      10'h22: dout  = 8'b00111111; //   34 :  63 - 0x3f
      10'h23: dout  = 8'b00110000; //   35 :  48 - 0x30
      10'h24: dout  = 8'b00111111; //   36 :  63 - 0x3f
      10'h25: dout  = 8'b00110000; //   37 :  48 - 0x30
      10'h26: dout  = 8'b00111111; //   38 :  63 - 0x3f
      10'h27: dout  = 8'b00110000; //   39 :  48 - 0x30
      10'h28: dout  = 8'b00111111; //   40 :  63 - 0x3f
      10'h29: dout  = 8'b00110000; //   41 :  48 - 0x30
      10'h2A: dout  = 8'b00111111; //   42 :  63 - 0x3f
      10'h2B: dout  = 8'b00110000; //   43 :  48 - 0x30
      10'h2C: dout  = 8'b00111111; //   44 :  63 - 0x3f
      10'h2D: dout  = 8'b00110000; //   45 :  48 - 0x30
      10'h2E: dout  = 8'b00111111; //   46 :  63 - 0x3f
      10'h2F: dout  = 8'b00110000; //   47 :  48 - 0x30
      10'h30: dout  = 8'b00111111; //   48 :  63 - 0x3f
      10'h31: dout  = 8'b00110000; //   49 :  48 - 0x30
      10'h32: dout  = 8'b00111111; //   50 :  63 - 0x3f
      10'h33: dout  = 8'b00110000; //   51 :  48 - 0x30
      10'h34: dout  = 8'b01100000; //   52 :  96 - 0x60
      10'h35: dout  = 8'b01110111; //   53 : 119 - 0x77
      10'h36: dout  = 8'b01110111; //   54 : 119 - 0x77
      10'h37: dout  = 8'b01110111; //   55 : 119 - 0x77
      10'h38: dout  = 8'b01110111; //   56 : 119 - 0x77
      10'h39: dout  = 8'b01110111; //   57 : 119 - 0x77
      10'h3A: dout  = 8'b01110111; //   58 : 119 - 0x77
      10'h3B: dout  = 8'b01110111; //   59 : 119 - 0x77
      10'h3C: dout  = 8'b01110111; //   60 : 119 - 0x77
      10'h3D: dout  = 8'b01110111; //   61 : 119 - 0x77
      10'h3E: dout  = 8'b01110111; //   62 : 119 - 0x77
      10'h3F: dout  = 8'b01110111; //   63 : 119 - 0x77
      10'h40: dout  = 8'b00110000; //   64 :  48 - 0x30 -- line 0x2
      10'h41: dout  = 8'b00111111; //   65 :  63 - 0x3f
      10'h42: dout  = 8'b00110000; //   66 :  48 - 0x30
      10'h43: dout  = 8'b00111111; //   67 :  63 - 0x3f
      10'h44: dout  = 8'b00110000; //   68 :  48 - 0x30
      10'h45: dout  = 8'b00111111; //   69 :  63 - 0x3f
      10'h46: dout  = 8'b00110000; //   70 :  48 - 0x30
      10'h47: dout  = 8'b00111111; //   71 :  63 - 0x3f
      10'h48: dout  = 8'b00110000; //   72 :  48 - 0x30
      10'h49: dout  = 8'b00111111; //   73 :  63 - 0x3f
      10'h4A: dout  = 8'b00110000; //   74 :  48 - 0x30
      10'h4B: dout  = 8'b00111111; //   75 :  63 - 0x3f
      10'h4C: dout  = 8'b00110000; //   76 :  48 - 0x30
      10'h4D: dout  = 8'b00111111; //   77 :  63 - 0x3f
      10'h4E: dout  = 8'b00110000; //   78 :  48 - 0x30
      10'h4F: dout  = 8'b00111111; //   79 :  63 - 0x3f
      10'h50: dout  = 8'b00110000; //   80 :  48 - 0x30
      10'h51: dout  = 8'b00111111; //   81 :  63 - 0x3f
      10'h52: dout  = 8'b00110000; //   82 :  48 - 0x30
      10'h53: dout  = 8'b00111111; //   83 :  63 - 0x3f
      10'h54: dout  = 8'b00111001; //   84 :  57 - 0x39
      10'h55: dout  = 8'b00111001; //   85 :  57 - 0x39
      10'h56: dout  = 8'b00111001; //   86 :  57 - 0x39
      10'h57: dout  = 8'b00111001; //   87 :  57 - 0x39
      10'h58: dout  = 8'b00111001; //   88 :  57 - 0x39
      10'h59: dout  = 8'b00111001; //   89 :  57 - 0x39
      10'h5A: dout  = 8'b00111001; //   90 :  57 - 0x39
      10'h5B: dout  = 8'b00111001; //   91 :  57 - 0x39
      10'h5C: dout  = 8'b00111001; //   92 :  57 - 0x39
      10'h5D: dout  = 8'b00111001; //   93 :  57 - 0x39
      10'h5E: dout  = 8'b00111001; //   94 :  57 - 0x39
      10'h5F: dout  = 8'b00111001; //   95 :  57 - 0x39
      10'h60: dout  = 8'b00111111; //   96 :  63 - 0x3f -- line 0x3
      10'h61: dout  = 8'b00110000; //   97 :  48 - 0x30
      10'h62: dout  = 8'b00111111; //   98 :  63 - 0x3f
      10'h63: dout  = 8'b00110000; //   99 :  48 - 0x30
      10'h64: dout  = 8'b00111111; //  100 :  63 - 0x3f
      10'h65: dout  = 8'b00110000; //  101 :  48 - 0x30
      10'h66: dout  = 8'b00111111; //  102 :  63 - 0x3f
      10'h67: dout  = 8'b00110000; //  103 :  48 - 0x30
      10'h68: dout  = 8'b00111111; //  104 :  63 - 0x3f
      10'h69: dout  = 8'b00110000; //  105 :  48 - 0x30
      10'h6A: dout  = 8'b00111111; //  106 :  63 - 0x3f
      10'h6B: dout  = 8'b00110000; //  107 :  48 - 0x30
      10'h6C: dout  = 8'b00111111; //  108 :  63 - 0x3f
      10'h6D: dout  = 8'b00110000; //  109 :  48 - 0x30
      10'h6E: dout  = 8'b00111111; //  110 :  63 - 0x3f
      10'h6F: dout  = 8'b00110000; //  111 :  48 - 0x30
      10'h70: dout  = 8'b00111111; //  112 :  63 - 0x3f
      10'h71: dout  = 8'b00110000; //  113 :  48 - 0x30
      10'h72: dout  = 8'b00111111; //  114 :  63 - 0x3f
      10'h73: dout  = 8'b00110000; //  115 :  48 - 0x30
      10'h74: dout  = 8'b00111111; //  116 :  63 - 0x3f
      10'h75: dout  = 8'b00111111; //  117 :  63 - 0x3f
      10'h76: dout  = 8'b00111111; //  118 :  63 - 0x3f
      10'h77: dout  = 8'b00111111; //  119 :  63 - 0x3f
      10'h78: dout  = 8'b00111111; //  120 :  63 - 0x3f
      10'h79: dout  = 8'b00111111; //  121 :  63 - 0x3f
      10'h7A: dout  = 8'b00111111; //  122 :  63 - 0x3f
      10'h7B: dout  = 8'b00111111; //  123 :  63 - 0x3f
      10'h7C: dout  = 8'b00111111; //  124 :  63 - 0x3f
      10'h7D: dout  = 8'b00111111; //  125 :  63 - 0x3f
      10'h7E: dout  = 8'b00111111; //  126 :  63 - 0x3f
      10'h7F: dout  = 8'b00111111; //  127 :  63 - 0x3f
      10'h80: dout  = 8'b00111111; //  128 :  63 - 0x3f -- line 0x4
      10'h81: dout  = 8'b00111111; //  129 :  63 - 0x3f
      10'h82: dout  = 8'b00111111; //  130 :  63 - 0x3f
      10'h83: dout  = 8'b00111111; //  131 :  63 - 0x3f
      10'h84: dout  = 8'b00111111; //  132 :  63 - 0x3f
      10'h85: dout  = 8'b00111111; //  133 :  63 - 0x3f
      10'h86: dout  = 8'b00111111; //  134 :  63 - 0x3f
      10'h87: dout  = 8'b00111111; //  135 :  63 - 0x3f
      10'h88: dout  = 8'b00111111; //  136 :  63 - 0x3f
      10'h89: dout  = 8'b00111111; //  137 :  63 - 0x3f
      10'h8A: dout  = 8'b00111111; //  138 :  63 - 0x3f
      10'h8B: dout  = 8'b00111111; //  139 :  63 - 0x3f
      10'h8C: dout  = 8'b00111111; //  140 :  63 - 0x3f
      10'h8D: dout  = 8'b00111111; //  141 :  63 - 0x3f
      10'h8E: dout  = 8'b00111111; //  142 :  63 - 0x3f
      10'h8F: dout  = 8'b00111111; //  143 :  63 - 0x3f
      10'h90: dout  = 8'b00111111; //  144 :  63 - 0x3f
      10'h91: dout  = 8'b00111111; //  145 :  63 - 0x3f
      10'h92: dout  = 8'b00111111; //  146 :  63 - 0x3f
      10'h93: dout  = 8'b00111111; //  147 :  63 - 0x3f
      10'h94: dout  = 8'b00111111; //  148 :  63 - 0x3f
      10'h95: dout  = 8'b00111111; //  149 :  63 - 0x3f
      10'h96: dout  = 8'b00111111; //  150 :  63 - 0x3f
      10'h97: dout  = 8'b00111111; //  151 :  63 - 0x3f
      10'h98: dout  = 8'b00111111; //  152 :  63 - 0x3f
      10'h99: dout  = 8'b00111111; //  153 :  63 - 0x3f
      10'h9A: dout  = 8'b00000100; //  154 :   4 - 0x4
      10'h9B: dout  = 8'b00000110; //  155 :   6 - 0x6
      10'h9C: dout  = 8'b00111111; //  156 :  63 - 0x3f
      10'h9D: dout  = 8'b00111111; //  157 :  63 - 0x3f
      10'h9E: dout  = 8'b00010100; //  158 :  20 - 0x14
      10'h9F: dout  = 8'b00010110; //  159 :  22 - 0x16
      10'hA0: dout  = 8'b00111111; //  160 :  63 - 0x3f -- line 0x5
      10'hA1: dout  = 8'b00111111; //  161 :  63 - 0x3f
      10'hA2: dout  = 8'b00111111; //  162 :  63 - 0x3f
      10'hA3: dout  = 8'b00111111; //  163 :  63 - 0x3f
      10'hA4: dout  = 8'b00111111; //  164 :  63 - 0x3f
      10'hA5: dout  = 8'b00111111; //  165 :  63 - 0x3f
      10'hA6: dout  = 8'b00111111; //  166 :  63 - 0x3f
      10'hA7: dout  = 8'b00111111; //  167 :  63 - 0x3f
      10'hA8: dout  = 8'b00111111; //  168 :  63 - 0x3f
      10'hA9: dout  = 8'b00111111; //  169 :  63 - 0x3f
      10'hAA: dout  = 8'b00111111; //  170 :  63 - 0x3f
      10'hAB: dout  = 8'b00111111; //  171 :  63 - 0x3f
      10'hAC: dout  = 8'b00111111; //  172 :  63 - 0x3f
      10'hAD: dout  = 8'b00111111; //  173 :  63 - 0x3f
      10'hAE: dout  = 8'b00111111; //  174 :  63 - 0x3f
      10'hAF: dout  = 8'b00111111; //  175 :  63 - 0x3f
      10'hB0: dout  = 8'b00111111; //  176 :  63 - 0x3f
      10'hB1: dout  = 8'b00111111; //  177 :  63 - 0x3f
      10'hB2: dout  = 8'b00111111; //  178 :  63 - 0x3f
      10'hB3: dout  = 8'b00111111; //  179 :  63 - 0x3f
      10'hB4: dout  = 8'b00111111; //  180 :  63 - 0x3f
      10'hB5: dout  = 8'b00111111; //  181 :  63 - 0x3f
      10'hB6: dout  = 8'b00111111; //  182 :  63 - 0x3f
      10'hB7: dout  = 8'b00111111; //  183 :  63 - 0x3f
      10'hB8: dout  = 8'b00111111; //  184 :  63 - 0x3f
      10'hB9: dout  = 8'b00111111; //  185 :  63 - 0x3f
      10'hBA: dout  = 8'b00000101; //  186 :   5 - 0x5
      10'hBB: dout  = 8'b00000111; //  187 :   7 - 0x7
      10'hBC: dout  = 8'b00111111; //  188 :  63 - 0x3f
      10'hBD: dout  = 8'b00111111; //  189 :  63 - 0x3f
      10'hBE: dout  = 8'b00010101; //  190 :  21 - 0x15
      10'hBF: dout  = 8'b00010111; //  191 :  23 - 0x17
      10'hC0: dout  = 8'b00111111; //  192 :  63 - 0x3f -- line 0x6
      10'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      10'hC2: dout  = 8'b00111111; //  194 :  63 - 0x3f
      10'hC3: dout  = 8'b00111111; //  195 :  63 - 0x3f
      10'hC4: dout  = 8'b00111111; //  196 :  63 - 0x3f
      10'hC5: dout  = 8'b00111111; //  197 :  63 - 0x3f
      10'hC6: dout  = 8'b00111111; //  198 :  63 - 0x3f
      10'hC7: dout  = 8'b00111111; //  199 :  63 - 0x3f
      10'hC8: dout  = 8'b00111111; //  200 :  63 - 0x3f
      10'hC9: dout  = 8'b00111111; //  201 :  63 - 0x3f
      10'hCA: dout  = 8'b00111111; //  202 :  63 - 0x3f
      10'hCB: dout  = 8'b00111111; //  203 :  63 - 0x3f
      10'hCC: dout  = 8'b00111111; //  204 :  63 - 0x3f
      10'hCD: dout  = 8'b00111111; //  205 :  63 - 0x3f
      10'hCE: dout  = 8'b00111111; //  206 :  63 - 0x3f
      10'hCF: dout  = 8'b00111111; //  207 :  63 - 0x3f
      10'hD0: dout  = 8'b00111111; //  208 :  63 - 0x3f
      10'hD1: dout  = 8'b00111111; //  209 :  63 - 0x3f
      10'hD2: dout  = 8'b00111111; //  210 :  63 - 0x3f
      10'hD3: dout  = 8'b00111111; //  211 :  63 - 0x3f
      10'hD4: dout  = 8'b00111111; //  212 :  63 - 0x3f
      10'hD5: dout  = 8'b00111111; //  213 :  63 - 0x3f
      10'hD6: dout  = 8'b00111111; //  214 :  63 - 0x3f
      10'hD7: dout  = 8'b00111111; //  215 :  63 - 0x3f
      10'hD8: dout  = 8'b00111111; //  216 :  63 - 0x3f
      10'hD9: dout  = 8'b00111111; //  217 :  63 - 0x3f
      10'hDA: dout  = 8'b00111111; //  218 :  63 - 0x3f
      10'hDB: dout  = 8'b00111111; //  219 :  63 - 0x3f
      10'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      10'hDD: dout  = 8'b00111111; //  221 :  63 - 0x3f
      10'hDE: dout  = 8'b00111111; //  222 :  63 - 0x3f
      10'hDF: dout  = 8'b00111111; //  223 :  63 - 0x3f
      10'hE0: dout  = 8'b00111111; //  224 :  63 - 0x3f -- line 0x7
      10'hE1: dout  = 8'b00111111; //  225 :  63 - 0x3f
      10'hE2: dout  = 8'b00111111; //  226 :  63 - 0x3f
      10'hE3: dout  = 8'b00111111; //  227 :  63 - 0x3f
      10'hE4: dout  = 8'b00111111; //  228 :  63 - 0x3f
      10'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      10'hE6: dout  = 8'b00111111; //  230 :  63 - 0x3f
      10'hE7: dout  = 8'b00111111; //  231 :  63 - 0x3f
      10'hE8: dout  = 8'b00111111; //  232 :  63 - 0x3f
      10'hE9: dout  = 8'b00111111; //  233 :  63 - 0x3f
      10'hEA: dout  = 8'b00111111; //  234 :  63 - 0x3f
      10'hEB: dout  = 8'b00111111; //  235 :  63 - 0x3f
      10'hEC: dout  = 8'b00111111; //  236 :  63 - 0x3f
      10'hED: dout  = 8'b00111111; //  237 :  63 - 0x3f
      10'hEE: dout  = 8'b00111111; //  238 :  63 - 0x3f
      10'hEF: dout  = 8'b00111111; //  239 :  63 - 0x3f
      10'hF0: dout  = 8'b00111111; //  240 :  63 - 0x3f
      10'hF1: dout  = 8'b00111111; //  241 :  63 - 0x3f
      10'hF2: dout  = 8'b00111111; //  242 :  63 - 0x3f
      10'hF3: dout  = 8'b00111111; //  243 :  63 - 0x3f
      10'hF4: dout  = 8'b00111111; //  244 :  63 - 0x3f
      10'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      10'hF6: dout  = 8'b00111111; //  246 :  63 - 0x3f
      10'hF7: dout  = 8'b00111111; //  247 :  63 - 0x3f
      10'hF8: dout  = 8'b00111111; //  248 :  63 - 0x3f
      10'hF9: dout  = 8'b00111111; //  249 :  63 - 0x3f
      10'hFA: dout  = 8'b00111111; //  250 :  63 - 0x3f
      10'hFB: dout  = 8'b00111111; //  251 :  63 - 0x3f
      10'hFC: dout  = 8'b00111111; //  252 :  63 - 0x3f
      10'hFD: dout  = 8'b00111111; //  253 :  63 - 0x3f
      10'hFE: dout  = 8'b00111111; //  254 :  63 - 0x3f
      10'hFF: dout  = 8'b00111111; //  255 :  63 - 0x3f
      10'h100: dout  = 8'b00111111; //  256 :  63 - 0x3f -- line 0x8
      10'h101: dout  = 8'b00111111; //  257 :  63 - 0x3f
      10'h102: dout  = 8'b00111111; //  258 :  63 - 0x3f
      10'h103: dout  = 8'b00111111; //  259 :  63 - 0x3f
      10'h104: dout  = 8'b00111111; //  260 :  63 - 0x3f
      10'h105: dout  = 8'b00111111; //  261 :  63 - 0x3f
      10'h106: dout  = 8'b00111111; //  262 :  63 - 0x3f
      10'h107: dout  = 8'b00111111; //  263 :  63 - 0x3f
      10'h108: dout  = 8'b00111111; //  264 :  63 - 0x3f
      10'h109: dout  = 8'b00111111; //  265 :  63 - 0x3f
      10'h10A: dout  = 8'b00111111; //  266 :  63 - 0x3f
      10'h10B: dout  = 8'b00111111; //  267 :  63 - 0x3f
      10'h10C: dout  = 8'b00111111; //  268 :  63 - 0x3f
      10'h10D: dout  = 8'b00111111; //  269 :  63 - 0x3f
      10'h10E: dout  = 8'b00111111; //  270 :  63 - 0x3f
      10'h10F: dout  = 8'b00111111; //  271 :  63 - 0x3f
      10'h110: dout  = 8'b00111111; //  272 :  63 - 0x3f
      10'h111: dout  = 8'b00111111; //  273 :  63 - 0x3f
      10'h112: dout  = 8'b00111111; //  274 :  63 - 0x3f
      10'h113: dout  = 8'b00111111; //  275 :  63 - 0x3f
      10'h114: dout  = 8'b00001100; //  276 :  12 - 0xc
      10'h115: dout  = 8'b00001110; //  277 :  14 - 0xe
      10'h116: dout  = 8'b00111111; //  278 :  63 - 0x3f
      10'h117: dout  = 8'b00111111; //  279 :  63 - 0x3f
      10'h118: dout  = 8'b00111111; //  280 :  63 - 0x3f
      10'h119: dout  = 8'b00111111; //  281 :  63 - 0x3f
      10'h11A: dout  = 8'b00111111; //  282 :  63 - 0x3f
      10'h11B: dout  = 8'b00111111; //  283 :  63 - 0x3f
      10'h11C: dout  = 8'b00111111; //  284 :  63 - 0x3f
      10'h11D: dout  = 8'b00111111; //  285 :  63 - 0x3f
      10'h11E: dout  = 8'b00111111; //  286 :  63 - 0x3f
      10'h11F: dout  = 8'b00111111; //  287 :  63 - 0x3f
      10'h120: dout  = 8'b00111111; //  288 :  63 - 0x3f -- line 0x9
      10'h121: dout  = 8'b00111111; //  289 :  63 - 0x3f
      10'h122: dout  = 8'b00111111; //  290 :  63 - 0x3f
      10'h123: dout  = 8'b00111111; //  291 :  63 - 0x3f
      10'h124: dout  = 8'b00111111; //  292 :  63 - 0x3f
      10'h125: dout  = 8'b00111111; //  293 :  63 - 0x3f
      10'h126: dout  = 8'b00111111; //  294 :  63 - 0x3f
      10'h127: dout  = 8'b00111111; //  295 :  63 - 0x3f
      10'h128: dout  = 8'b00111111; //  296 :  63 - 0x3f
      10'h129: dout  = 8'b00111111; //  297 :  63 - 0x3f
      10'h12A: dout  = 8'b00111111; //  298 :  63 - 0x3f
      10'h12B: dout  = 8'b00111111; //  299 :  63 - 0x3f
      10'h12C: dout  = 8'b00111111; //  300 :  63 - 0x3f
      10'h12D: dout  = 8'b00111111; //  301 :  63 - 0x3f
      10'h12E: dout  = 8'b00111111; //  302 :  63 - 0x3f
      10'h12F: dout  = 8'b00111111; //  303 :  63 - 0x3f
      10'h130: dout  = 8'b00111111; //  304 :  63 - 0x3f
      10'h131: dout  = 8'b00111111; //  305 :  63 - 0x3f
      10'h132: dout  = 8'b00111111; //  306 :  63 - 0x3f
      10'h133: dout  = 8'b00111111; //  307 :  63 - 0x3f
      10'h134: dout  = 8'b00001101; //  308 :  13 - 0xd
      10'h135: dout  = 8'b00001111; //  309 :  15 - 0xf
      10'h136: dout  = 8'b00111111; //  310 :  63 - 0x3f
      10'h137: dout  = 8'b00111111; //  311 :  63 - 0x3f
      10'h138: dout  = 8'b00111111; //  312 :  63 - 0x3f
      10'h139: dout  = 8'b00111111; //  313 :  63 - 0x3f
      10'h13A: dout  = 8'b00111111; //  314 :  63 - 0x3f
      10'h13B: dout  = 8'b00111111; //  315 :  63 - 0x3f
      10'h13C: dout  = 8'b00111111; //  316 :  63 - 0x3f
      10'h13D: dout  = 8'b00111111; //  317 :  63 - 0x3f
      10'h13E: dout  = 8'b00111111; //  318 :  63 - 0x3f
      10'h13F: dout  = 8'b00111111; //  319 :  63 - 0x3f
      10'h140: dout  = 8'b00111111; //  320 :  63 - 0x3f -- line 0xa
      10'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      10'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      10'h143: dout  = 8'b00111111; //  323 :  63 - 0x3f
      10'h144: dout  = 8'b00111111; //  324 :  63 - 0x3f
      10'h145: dout  = 8'b00111111; //  325 :  63 - 0x3f
      10'h146: dout  = 8'b00111111; //  326 :  63 - 0x3f
      10'h147: dout  = 8'b00111111; //  327 :  63 - 0x3f
      10'h148: dout  = 8'b00111111; //  328 :  63 - 0x3f
      10'h149: dout  = 8'b00111111; //  329 :  63 - 0x3f
      10'h14A: dout  = 8'b00111111; //  330 :  63 - 0x3f
      10'h14B: dout  = 8'b00111111; //  331 :  63 - 0x3f
      10'h14C: dout  = 8'b00111111; //  332 :  63 - 0x3f
      10'h14D: dout  = 8'b00111111; //  333 :  63 - 0x3f
      10'h14E: dout  = 8'b00111111; //  334 :  63 - 0x3f
      10'h14F: dout  = 8'b00111111; //  335 :  63 - 0x3f
      10'h150: dout  = 8'b00111111; //  336 :  63 - 0x3f
      10'h151: dout  = 8'b00111111; //  337 :  63 - 0x3f
      10'h152: dout  = 8'b00111111; //  338 :  63 - 0x3f
      10'h153: dout  = 8'b00111111; //  339 :  63 - 0x3f
      10'h154: dout  = 8'b01010111; //  340 :  87 - 0x57
      10'h155: dout  = 8'b01011000; //  341 :  88 - 0x58
      10'h156: dout  = 8'b01011000; //  342 :  88 - 0x58
      10'h157: dout  = 8'b01011000; //  343 :  88 - 0x58
      10'h158: dout  = 8'b01011000; //  344 :  88 - 0x58
      10'h159: dout  = 8'b01011000; //  345 :  88 - 0x58
      10'h15A: dout  = 8'b01011000; //  346 :  88 - 0x58
      10'h15B: dout  = 8'b01011000; //  347 :  88 - 0x58
      10'h15C: dout  = 8'b01011000; //  348 :  88 - 0x58
      10'h15D: dout  = 8'b01011000; //  349 :  88 - 0x58
      10'h15E: dout  = 8'b01011000; //  350 :  88 - 0x58
      10'h15F: dout  = 8'b01011000; //  351 :  88 - 0x58
      10'h160: dout  = 8'b00111111; //  352 :  63 - 0x3f -- line 0xb
      10'h161: dout  = 8'b00111111; //  353 :  63 - 0x3f
      10'h162: dout  = 8'b00111111; //  354 :  63 - 0x3f
      10'h163: dout  = 8'b00111111; //  355 :  63 - 0x3f
      10'h164: dout  = 8'b00111111; //  356 :  63 - 0x3f
      10'h165: dout  = 8'b00111111; //  357 :  63 - 0x3f
      10'h166: dout  = 8'b00111111; //  358 :  63 - 0x3f
      10'h167: dout  = 8'b00111111; //  359 :  63 - 0x3f
      10'h168: dout  = 8'b00111111; //  360 :  63 - 0x3f
      10'h169: dout  = 8'b00111111; //  361 :  63 - 0x3f
      10'h16A: dout  = 8'b00111111; //  362 :  63 - 0x3f
      10'h16B: dout  = 8'b00111111; //  363 :  63 - 0x3f
      10'h16C: dout  = 8'b00111111; //  364 :  63 - 0x3f
      10'h16D: dout  = 8'b00111111; //  365 :  63 - 0x3f
      10'h16E: dout  = 8'b00111111; //  366 :  63 - 0x3f
      10'h16F: dout  = 8'b00111111; //  367 :  63 - 0x3f
      10'h170: dout  = 8'b00111111; //  368 :  63 - 0x3f
      10'h171: dout  = 8'b00111111; //  369 :  63 - 0x3f
      10'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      10'h173: dout  = 8'b00111111; //  371 :  63 - 0x3f
      10'h174: dout  = 8'b00111111; //  372 :  63 - 0x3f
      10'h175: dout  = 8'b00111111; //  373 :  63 - 0x3f
      10'h176: dout  = 8'b00111111; //  374 :  63 - 0x3f
      10'h177: dout  = 8'b00111111; //  375 :  63 - 0x3f
      10'h178: dout  = 8'b00111111; //  376 :  63 - 0x3f
      10'h179: dout  = 8'b00111111; //  377 :  63 - 0x3f
      10'h17A: dout  = 8'b00111111; //  378 :  63 - 0x3f
      10'h17B: dout  = 8'b00111111; //  379 :  63 - 0x3f
      10'h17C: dout  = 8'b00111111; //  380 :  63 - 0x3f
      10'h17D: dout  = 8'b00111111; //  381 :  63 - 0x3f
      10'h17E: dout  = 8'b00111111; //  382 :  63 - 0x3f
      10'h17F: dout  = 8'b00111111; //  383 :  63 - 0x3f
      10'h180: dout  = 8'b00111111; //  384 :  63 - 0x3f -- line 0xc
      10'h181: dout  = 8'b00111111; //  385 :  63 - 0x3f
      10'h182: dout  = 8'b00111111; //  386 :  63 - 0x3f
      10'h183: dout  = 8'b00111111; //  387 :  63 - 0x3f
      10'h184: dout  = 8'b00111111; //  388 :  63 - 0x3f
      10'h185: dout  = 8'b00111111; //  389 :  63 - 0x3f
      10'h186: dout  = 8'b00111111; //  390 :  63 - 0x3f
      10'h187: dout  = 8'b00111111; //  391 :  63 - 0x3f
      10'h188: dout  = 8'b00111111; //  392 :  63 - 0x3f
      10'h189: dout  = 8'b00111111; //  393 :  63 - 0x3f
      10'h18A: dout  = 8'b00111111; //  394 :  63 - 0x3f
      10'h18B: dout  = 8'b00111111; //  395 :  63 - 0x3f
      10'h18C: dout  = 8'b00111111; //  396 :  63 - 0x3f
      10'h18D: dout  = 8'b00111111; //  397 :  63 - 0x3f
      10'h18E: dout  = 8'b00111111; //  398 :  63 - 0x3f
      10'h18F: dout  = 8'b00111111; //  399 :  63 - 0x3f
      10'h190: dout  = 8'b00111111; //  400 :  63 - 0x3f
      10'h191: dout  = 8'b00111111; //  401 :  63 - 0x3f
      10'h192: dout  = 8'b00111111; //  402 :  63 - 0x3f
      10'h193: dout  = 8'b00111111; //  403 :  63 - 0x3f
      10'h194: dout  = 8'b00111111; //  404 :  63 - 0x3f
      10'h195: dout  = 8'b00111111; //  405 :  63 - 0x3f
      10'h196: dout  = 8'b00111111; //  406 :  63 - 0x3f
      10'h197: dout  = 8'b00111111; //  407 :  63 - 0x3f
      10'h198: dout  = 8'b00111111; //  408 :  63 - 0x3f
      10'h199: dout  = 8'b00111111; //  409 :  63 - 0x3f
      10'h19A: dout  = 8'b00111111; //  410 :  63 - 0x3f
      10'h19B: dout  = 8'b00111111; //  411 :  63 - 0x3f
      10'h19C: dout  = 8'b00111111; //  412 :  63 - 0x3f
      10'h19D: dout  = 8'b00111111; //  413 :  63 - 0x3f
      10'h19E: dout  = 8'b00111111; //  414 :  63 - 0x3f
      10'h19F: dout  = 8'b00111111; //  415 :  63 - 0x3f
      10'h1A0: dout  = 8'b00111111; //  416 :  63 - 0x3f -- line 0xd
      10'h1A1: dout  = 8'b00111111; //  417 :  63 - 0x3f
      10'h1A2: dout  = 8'b00111111; //  418 :  63 - 0x3f
      10'h1A3: dout  = 8'b00111111; //  419 :  63 - 0x3f
      10'h1A4: dout  = 8'b00111111; //  420 :  63 - 0x3f
      10'h1A5: dout  = 8'b00111111; //  421 :  63 - 0x3f
      10'h1A6: dout  = 8'b00111111; //  422 :  63 - 0x3f
      10'h1A7: dout  = 8'b00111111; //  423 :  63 - 0x3f
      10'h1A8: dout  = 8'b00111111; //  424 :  63 - 0x3f
      10'h1A9: dout  = 8'b00111111; //  425 :  63 - 0x3f
      10'h1AA: dout  = 8'b00111111; //  426 :  63 - 0x3f
      10'h1AB: dout  = 8'b00111111; //  427 :  63 - 0x3f
      10'h1AC: dout  = 8'b00111111; //  428 :  63 - 0x3f
      10'h1AD: dout  = 8'b00111111; //  429 :  63 - 0x3f
      10'h1AE: dout  = 8'b00111111; //  430 :  63 - 0x3f
      10'h1AF: dout  = 8'b00111111; //  431 :  63 - 0x3f
      10'h1B0: dout  = 8'b00111111; //  432 :  63 - 0x3f
      10'h1B1: dout  = 8'b00111111; //  433 :  63 - 0x3f
      10'h1B2: dout  = 8'b00111111; //  434 :  63 - 0x3f
      10'h1B3: dout  = 8'b00111111; //  435 :  63 - 0x3f
      10'h1B4: dout  = 8'b00111111; //  436 :  63 - 0x3f
      10'h1B5: dout  = 8'b00111111; //  437 :  63 - 0x3f
      10'h1B6: dout  = 8'b00111111; //  438 :  63 - 0x3f
      10'h1B7: dout  = 8'b00111111; //  439 :  63 - 0x3f
      10'h1B8: dout  = 8'b00111111; //  440 :  63 - 0x3f
      10'h1B9: dout  = 8'b00111111; //  441 :  63 - 0x3f
      10'h1BA: dout  = 8'b00111111; //  442 :  63 - 0x3f
      10'h1BB: dout  = 8'b00111111; //  443 :  63 - 0x3f
      10'h1BC: dout  = 8'b00111111; //  444 :  63 - 0x3f
      10'h1BD: dout  = 8'b00111111; //  445 :  63 - 0x3f
      10'h1BE: dout  = 8'b00111111; //  446 :  63 - 0x3f
      10'h1BF: dout  = 8'b00111111; //  447 :  63 - 0x3f
      10'h1C0: dout  = 8'b00111111; //  448 :  63 - 0x3f -- line 0xe
      10'h1C1: dout  = 8'b00111111; //  449 :  63 - 0x3f
      10'h1C2: dout  = 8'b00111111; //  450 :  63 - 0x3f
      10'h1C3: dout  = 8'b00111111; //  451 :  63 - 0x3f
      10'h1C4: dout  = 8'b00111111; //  452 :  63 - 0x3f
      10'h1C5: dout  = 8'b00111111; //  453 :  63 - 0x3f
      10'h1C6: dout  = 8'b00111111; //  454 :  63 - 0x3f
      10'h1C7: dout  = 8'b00111111; //  455 :  63 - 0x3f
      10'h1C8: dout  = 8'b00111111; //  456 :  63 - 0x3f
      10'h1C9: dout  = 8'b00111111; //  457 :  63 - 0x3f
      10'h1CA: dout  = 8'b00111111; //  458 :  63 - 0x3f
      10'h1CB: dout  = 8'b00111111; //  459 :  63 - 0x3f
      10'h1CC: dout  = 8'b00111111; //  460 :  63 - 0x3f
      10'h1CD: dout  = 8'b00111111; //  461 :  63 - 0x3f
      10'h1CE: dout  = 8'b00111111; //  462 :  63 - 0x3f
      10'h1CF: dout  = 8'b00111111; //  463 :  63 - 0x3f
      10'h1D0: dout  = 8'b00111111; //  464 :  63 - 0x3f
      10'h1D1: dout  = 8'b00111111; //  465 :  63 - 0x3f
      10'h1D2: dout  = 8'b00111111; //  466 :  63 - 0x3f
      10'h1D3: dout  = 8'b00111111; //  467 :  63 - 0x3f
      10'h1D4: dout  = 8'b00111111; //  468 :  63 - 0x3f
      10'h1D5: dout  = 8'b00111111; //  469 :  63 - 0x3f
      10'h1D6: dout  = 8'b00111111; //  470 :  63 - 0x3f
      10'h1D7: dout  = 8'b00111111; //  471 :  63 - 0x3f
      10'h1D8: dout  = 8'b00111111; //  472 :  63 - 0x3f
      10'h1D9: dout  = 8'b00111111; //  473 :  63 - 0x3f
      10'h1DA: dout  = 8'b00111111; //  474 :  63 - 0x3f
      10'h1DB: dout  = 8'b00111111; //  475 :  63 - 0x3f
      10'h1DC: dout  = 8'b00111111; //  476 :  63 - 0x3f
      10'h1DD: dout  = 8'b00111111; //  477 :  63 - 0x3f
      10'h1DE: dout  = 8'b00111111; //  478 :  63 - 0x3f
      10'h1DF: dout  = 8'b00111111; //  479 :  63 - 0x3f
      10'h1E0: dout  = 8'b00111111; //  480 :  63 - 0x3f -- line 0xf
      10'h1E1: dout  = 8'b00111111; //  481 :  63 - 0x3f
      10'h1E2: dout  = 8'b00111111; //  482 :  63 - 0x3f
      10'h1E3: dout  = 8'b00111111; //  483 :  63 - 0x3f
      10'h1E4: dout  = 8'b00111111; //  484 :  63 - 0x3f
      10'h1E5: dout  = 8'b00111111; //  485 :  63 - 0x3f
      10'h1E6: dout  = 8'b00111111; //  486 :  63 - 0x3f
      10'h1E7: dout  = 8'b00111111; //  487 :  63 - 0x3f
      10'h1E8: dout  = 8'b00111111; //  488 :  63 - 0x3f
      10'h1E9: dout  = 8'b00111111; //  489 :  63 - 0x3f
      10'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      10'h1EB: dout  = 8'b00111111; //  491 :  63 - 0x3f
      10'h1EC: dout  = 8'b00111111; //  492 :  63 - 0x3f
      10'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      10'h1EE: dout  = 8'b00111111; //  494 :  63 - 0x3f
      10'h1EF: dout  = 8'b00111111; //  495 :  63 - 0x3f
      10'h1F0: dout  = 8'b00111111; //  496 :  63 - 0x3f
      10'h1F1: dout  = 8'b00111111; //  497 :  63 - 0x3f
      10'h1F2: dout  = 8'b00111111; //  498 :  63 - 0x3f
      10'h1F3: dout  = 8'b00111111; //  499 :  63 - 0x3f
      10'h1F4: dout  = 8'b00111111; //  500 :  63 - 0x3f
      10'h1F5: dout  = 8'b00111111; //  501 :  63 - 0x3f
      10'h1F6: dout  = 8'b00111111; //  502 :  63 - 0x3f
      10'h1F7: dout  = 8'b00111111; //  503 :  63 - 0x3f
      10'h1F8: dout  = 8'b00111111; //  504 :  63 - 0x3f
      10'h1F9: dout  = 8'b00111111; //  505 :  63 - 0x3f
      10'h1FA: dout  = 8'b00111111; //  506 :  63 - 0x3f
      10'h1FB: dout  = 8'b00111111; //  507 :  63 - 0x3f
      10'h1FC: dout  = 8'b00111111; //  508 :  63 - 0x3f
      10'h1FD: dout  = 8'b00111111; //  509 :  63 - 0x3f
      10'h1FE: dout  = 8'b00111111; //  510 :  63 - 0x3f
      10'h1FF: dout  = 8'b00111111; //  511 :  63 - 0x3f
      10'h200: dout  = 8'b00111111; //  512 :  63 - 0x3f -- line 0x10
      10'h201: dout  = 8'b00111111; //  513 :  63 - 0x3f
      10'h202: dout  = 8'b00111111; //  514 :  63 - 0x3f
      10'h203: dout  = 8'b00111111; //  515 :  63 - 0x3f
      10'h204: dout  = 8'b00111111; //  516 :  63 - 0x3f
      10'h205: dout  = 8'b00111111; //  517 :  63 - 0x3f
      10'h206: dout  = 8'b00111111; //  518 :  63 - 0x3f
      10'h207: dout  = 8'b00111111; //  519 :  63 - 0x3f
      10'h208: dout  = 8'b00111111; //  520 :  63 - 0x3f
      10'h209: dout  = 8'b00111111; //  521 :  63 - 0x3f
      10'h20A: dout  = 8'b00111111; //  522 :  63 - 0x3f
      10'h20B: dout  = 8'b00111111; //  523 :  63 - 0x3f
      10'h20C: dout  = 8'b00111111; //  524 :  63 - 0x3f
      10'h20D: dout  = 8'b00111111; //  525 :  63 - 0x3f
      10'h20E: dout  = 8'b00111111; //  526 :  63 - 0x3f
      10'h20F: dout  = 8'b00111111; //  527 :  63 - 0x3f
      10'h210: dout  = 8'b00111111; //  528 :  63 - 0x3f
      10'h211: dout  = 8'b00111111; //  529 :  63 - 0x3f
      10'h212: dout  = 8'b00111111; //  530 :  63 - 0x3f
      10'h213: dout  = 8'b00111111; //  531 :  63 - 0x3f
      10'h214: dout  = 8'b00111111; //  532 :  63 - 0x3f
      10'h215: dout  = 8'b00111111; //  533 :  63 - 0x3f
      10'h216: dout  = 8'b00111111; //  534 :  63 - 0x3f
      10'h217: dout  = 8'b00111111; //  535 :  63 - 0x3f
      10'h218: dout  = 8'b00111111; //  536 :  63 - 0x3f
      10'h219: dout  = 8'b00111111; //  537 :  63 - 0x3f
      10'h21A: dout  = 8'b00111111; //  538 :  63 - 0x3f
      10'h21B: dout  = 8'b00111111; //  539 :  63 - 0x3f
      10'h21C: dout  = 8'b00111111; //  540 :  63 - 0x3f
      10'h21D: dout  = 8'b00111111; //  541 :  63 - 0x3f
      10'h21E: dout  = 8'b00111111; //  542 :  63 - 0x3f
      10'h21F: dout  = 8'b00111111; //  543 :  63 - 0x3f
      10'h220: dout  = 8'b00111111; //  544 :  63 - 0x3f -- line 0x11
      10'h221: dout  = 8'b00111111; //  545 :  63 - 0x3f
      10'h222: dout  = 8'b00111111; //  546 :  63 - 0x3f
      10'h223: dout  = 8'b00111111; //  547 :  63 - 0x3f
      10'h224: dout  = 8'b00111111; //  548 :  63 - 0x3f
      10'h225: dout  = 8'b00111111; //  549 :  63 - 0x3f
      10'h226: dout  = 8'b00111111; //  550 :  63 - 0x3f
      10'h227: dout  = 8'b00111111; //  551 :  63 - 0x3f
      10'h228: dout  = 8'b00111111; //  552 :  63 - 0x3f
      10'h229: dout  = 8'b00111111; //  553 :  63 - 0x3f
      10'h22A: dout  = 8'b00111111; //  554 :  63 - 0x3f
      10'h22B: dout  = 8'b00111111; //  555 :  63 - 0x3f
      10'h22C: dout  = 8'b00111111; //  556 :  63 - 0x3f
      10'h22D: dout  = 8'b00111111; //  557 :  63 - 0x3f
      10'h22E: dout  = 8'b00111111; //  558 :  63 - 0x3f
      10'h22F: dout  = 8'b00111111; //  559 :  63 - 0x3f
      10'h230: dout  = 8'b00111111; //  560 :  63 - 0x3f
      10'h231: dout  = 8'b00111111; //  561 :  63 - 0x3f
      10'h232: dout  = 8'b00111111; //  562 :  63 - 0x3f
      10'h233: dout  = 8'b00111111; //  563 :  63 - 0x3f
      10'h234: dout  = 8'b00111111; //  564 :  63 - 0x3f
      10'h235: dout  = 8'b00111111; //  565 :  63 - 0x3f
      10'h236: dout  = 8'b00111111; //  566 :  63 - 0x3f
      10'h237: dout  = 8'b00111111; //  567 :  63 - 0x3f
      10'h238: dout  = 8'b00111111; //  568 :  63 - 0x3f
      10'h239: dout  = 8'b00111111; //  569 :  63 - 0x3f
      10'h23A: dout  = 8'b00111111; //  570 :  63 - 0x3f
      10'h23B: dout  = 8'b00111111; //  571 :  63 - 0x3f
      10'h23C: dout  = 8'b00111111; //  572 :  63 - 0x3f
      10'h23D: dout  = 8'b00111111; //  573 :  63 - 0x3f
      10'h23E: dout  = 8'b00111111; //  574 :  63 - 0x3f
      10'h23F: dout  = 8'b00111111; //  575 :  63 - 0x3f
      10'h240: dout  = 8'b00111111; //  576 :  63 - 0x3f -- line 0x12
      10'h241: dout  = 8'b00111111; //  577 :  63 - 0x3f
      10'h242: dout  = 8'b00111111; //  578 :  63 - 0x3f
      10'h243: dout  = 8'b00111111; //  579 :  63 - 0x3f
      10'h244: dout  = 8'b00111111; //  580 :  63 - 0x3f
      10'h245: dout  = 8'b00111111; //  581 :  63 - 0x3f
      10'h246: dout  = 8'b00111111; //  582 :  63 - 0x3f
      10'h247: dout  = 8'b00111111; //  583 :  63 - 0x3f
      10'h248: dout  = 8'b00111111; //  584 :  63 - 0x3f
      10'h249: dout  = 8'b00111111; //  585 :  63 - 0x3f
      10'h24A: dout  = 8'b00111111; //  586 :  63 - 0x3f
      10'h24B: dout  = 8'b00111111; //  587 :  63 - 0x3f
      10'h24C: dout  = 8'b00111111; //  588 :  63 - 0x3f
      10'h24D: dout  = 8'b00111111; //  589 :  63 - 0x3f
      10'h24E: dout  = 8'b00111111; //  590 :  63 - 0x3f
      10'h24F: dout  = 8'b00111111; //  591 :  63 - 0x3f
      10'h250: dout  = 8'b00000000; //  592 :   0 - 0x0
      10'h251: dout  = 8'b00000010; //  593 :   2 - 0x2
      10'h252: dout  = 8'b00000000; //  594 :   0 - 0x0
      10'h253: dout  = 8'b00000010; //  595 :   2 - 0x2
      10'h254: dout  = 8'b00000000; //  596 :   0 - 0x0
      10'h255: dout  = 8'b00000010; //  597 :   2 - 0x2
      10'h256: dout  = 8'b00000100; //  598 :   4 - 0x4
      10'h257: dout  = 8'b00000110; //  599 :   6 - 0x6
      10'h258: dout  = 8'b00000000; //  600 :   0 - 0x0
      10'h259: dout  = 8'b00000010; //  601 :   2 - 0x2
      10'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      10'h25B: dout  = 8'b00000010; //  603 :   2 - 0x2
      10'h25C: dout  = 8'b00000100; //  604 :   4 - 0x4
      10'h25D: dout  = 8'b00000110; //  605 :   6 - 0x6
      10'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      10'h25F: dout  = 8'b00000010; //  607 :   2 - 0x2
      10'h260: dout  = 8'b00111111; //  608 :  63 - 0x3f -- line 0x13
      10'h261: dout  = 8'b00111111; //  609 :  63 - 0x3f
      10'h262: dout  = 8'b00111111; //  610 :  63 - 0x3f
      10'h263: dout  = 8'b00111111; //  611 :  63 - 0x3f
      10'h264: dout  = 8'b00111111; //  612 :  63 - 0x3f
      10'h265: dout  = 8'b00111111; //  613 :  63 - 0x3f
      10'h266: dout  = 8'b00111111; //  614 :  63 - 0x3f
      10'h267: dout  = 8'b00111111; //  615 :  63 - 0x3f
      10'h268: dout  = 8'b00111111; //  616 :  63 - 0x3f
      10'h269: dout  = 8'b00111111; //  617 :  63 - 0x3f
      10'h26A: dout  = 8'b00111111; //  618 :  63 - 0x3f
      10'h26B: dout  = 8'b00111111; //  619 :  63 - 0x3f
      10'h26C: dout  = 8'b00111111; //  620 :  63 - 0x3f
      10'h26D: dout  = 8'b00111111; //  621 :  63 - 0x3f
      10'h26E: dout  = 8'b00111111; //  622 :  63 - 0x3f
      10'h26F: dout  = 8'b00111111; //  623 :  63 - 0x3f
      10'h270: dout  = 8'b00000001; //  624 :   1 - 0x1
      10'h271: dout  = 8'b00000011; //  625 :   3 - 0x3
      10'h272: dout  = 8'b00000001; //  626 :   1 - 0x1
      10'h273: dout  = 8'b00000011; //  627 :   3 - 0x3
      10'h274: dout  = 8'b00000001; //  628 :   1 - 0x1
      10'h275: dout  = 8'b00000011; //  629 :   3 - 0x3
      10'h276: dout  = 8'b00000101; //  630 :   5 - 0x5
      10'h277: dout  = 8'b00000111; //  631 :   7 - 0x7
      10'h278: dout  = 8'b00000001; //  632 :   1 - 0x1
      10'h279: dout  = 8'b00000011; //  633 :   3 - 0x3
      10'h27A: dout  = 8'b00000001; //  634 :   1 - 0x1
      10'h27B: dout  = 8'b00000011; //  635 :   3 - 0x3
      10'h27C: dout  = 8'b00000101; //  636 :   5 - 0x5
      10'h27D: dout  = 8'b00000111; //  637 :   7 - 0x7
      10'h27E: dout  = 8'b00000001; //  638 :   1 - 0x1
      10'h27F: dout  = 8'b00000011; //  639 :   3 - 0x3
      10'h280: dout  = 8'b00111111; //  640 :  63 - 0x3f -- line 0x14
      10'h281: dout  = 8'b00111111; //  641 :  63 - 0x3f
      10'h282: dout  = 8'b00111111; //  642 :  63 - 0x3f
      10'h283: dout  = 8'b00111111; //  643 :  63 - 0x3f
      10'h284: dout  = 8'b00111111; //  644 :  63 - 0x3f
      10'h285: dout  = 8'b00111111; //  645 :  63 - 0x3f
      10'h286: dout  = 8'b00111111; //  646 :  63 - 0x3f
      10'h287: dout  = 8'b00111111; //  647 :  63 - 0x3f
      10'h288: dout  = 8'b00111111; //  648 :  63 - 0x3f
      10'h289: dout  = 8'b00111111; //  649 :  63 - 0x3f
      10'h28A: dout  = 8'b00111111; //  650 :  63 - 0x3f
      10'h28B: dout  = 8'b00111111; //  651 :  63 - 0x3f
      10'h28C: dout  = 8'b00111111; //  652 :  63 - 0x3f
      10'h28D: dout  = 8'b00111111; //  653 :  63 - 0x3f
      10'h28E: dout  = 8'b00111111; //  654 :  63 - 0x3f
      10'h28F: dout  = 8'b00111111; //  655 :  63 - 0x3f
      10'h290: dout  = 8'b00111111; //  656 :  63 - 0x3f
      10'h291: dout  = 8'b00111111; //  657 :  63 - 0x3f
      10'h292: dout  = 8'b00111111; //  658 :  63 - 0x3f
      10'h293: dout  = 8'b00111111; //  659 :  63 - 0x3f
      10'h294: dout  = 8'b00111111; //  660 :  63 - 0x3f
      10'h295: dout  = 8'b00111111; //  661 :  63 - 0x3f
      10'h296: dout  = 8'b00111111; //  662 :  63 - 0x3f
      10'h297: dout  = 8'b00111111; //  663 :  63 - 0x3f
      10'h298: dout  = 8'b00111111; //  664 :  63 - 0x3f
      10'h299: dout  = 8'b00111111; //  665 :  63 - 0x3f
      10'h29A: dout  = 8'b00111111; //  666 :  63 - 0x3f
      10'h29B: dout  = 8'b00111111; //  667 :  63 - 0x3f
      10'h29C: dout  = 8'b00111111; //  668 :  63 - 0x3f
      10'h29D: dout  = 8'b00111111; //  669 :  63 - 0x3f
      10'h29E: dout  = 8'b00111111; //  670 :  63 - 0x3f
      10'h29F: dout  = 8'b00111111; //  671 :  63 - 0x3f
      10'h2A0: dout  = 8'b00111111; //  672 :  63 - 0x3f -- line 0x15
      10'h2A1: dout  = 8'b00111111; //  673 :  63 - 0x3f
      10'h2A2: dout  = 8'b00111111; //  674 :  63 - 0x3f
      10'h2A3: dout  = 8'b00111111; //  675 :  63 - 0x3f
      10'h2A4: dout  = 8'b00111111; //  676 :  63 - 0x3f
      10'h2A5: dout  = 8'b00111111; //  677 :  63 - 0x3f
      10'h2A6: dout  = 8'b00111111; //  678 :  63 - 0x3f
      10'h2A7: dout  = 8'b00111111; //  679 :  63 - 0x3f
      10'h2A8: dout  = 8'b00111111; //  680 :  63 - 0x3f
      10'h2A9: dout  = 8'b00111111; //  681 :  63 - 0x3f
      10'h2AA: dout  = 8'b00111111; //  682 :  63 - 0x3f
      10'h2AB: dout  = 8'b00111111; //  683 :  63 - 0x3f
      10'h2AC: dout  = 8'b00111111; //  684 :  63 - 0x3f
      10'h2AD: dout  = 8'b00111111; //  685 :  63 - 0x3f
      10'h2AE: dout  = 8'b00111111; //  686 :  63 - 0x3f
      10'h2AF: dout  = 8'b00111111; //  687 :  63 - 0x3f
      10'h2B0: dout  = 8'b00111111; //  688 :  63 - 0x3f
      10'h2B1: dout  = 8'b00111111; //  689 :  63 - 0x3f
      10'h2B2: dout  = 8'b00111111; //  690 :  63 - 0x3f
      10'h2B3: dout  = 8'b00111111; //  691 :  63 - 0x3f
      10'h2B4: dout  = 8'b00111111; //  692 :  63 - 0x3f
      10'h2B5: dout  = 8'b00111111; //  693 :  63 - 0x3f
      10'h2B6: dout  = 8'b00111111; //  694 :  63 - 0x3f
      10'h2B7: dout  = 8'b00111111; //  695 :  63 - 0x3f
      10'h2B8: dout  = 8'b00111111; //  696 :  63 - 0x3f
      10'h2B9: dout  = 8'b00111111; //  697 :  63 - 0x3f
      10'h2BA: dout  = 8'b00111111; //  698 :  63 - 0x3f
      10'h2BB: dout  = 8'b00111111; //  699 :  63 - 0x3f
      10'h2BC: dout  = 8'b00111111; //  700 :  63 - 0x3f
      10'h2BD: dout  = 8'b00111111; //  701 :  63 - 0x3f
      10'h2BE: dout  = 8'b00111111; //  702 :  63 - 0x3f
      10'h2BF: dout  = 8'b00111111; //  703 :  63 - 0x3f
      10'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- line 0x16
      10'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      10'h2C2: dout  = 8'b00111111; //  706 :  63 - 0x3f
      10'h2C3: dout  = 8'b00111111; //  707 :  63 - 0x3f
      10'h2C4: dout  = 8'b00111111; //  708 :  63 - 0x3f
      10'h2C5: dout  = 8'b00111111; //  709 :  63 - 0x3f
      10'h2C6: dout  = 8'b00111111; //  710 :  63 - 0x3f
      10'h2C7: dout  = 8'b00111111; //  711 :  63 - 0x3f
      10'h2C8: dout  = 8'b00111111; //  712 :  63 - 0x3f
      10'h2C9: dout  = 8'b00111111; //  713 :  63 - 0x3f
      10'h2CA: dout  = 8'b00111111; //  714 :  63 - 0x3f
      10'h2CB: dout  = 8'b00111111; //  715 :  63 - 0x3f
      10'h2CC: dout  = 8'b00111111; //  716 :  63 - 0x3f
      10'h2CD: dout  = 8'b00111111; //  717 :  63 - 0x3f
      10'h2CE: dout  = 8'b00111111; //  718 :  63 - 0x3f
      10'h2CF: dout  = 8'b00111111; //  719 :  63 - 0x3f
      10'h2D0: dout  = 8'b00111111; //  720 :  63 - 0x3f
      10'h2D1: dout  = 8'b00111111; //  721 :  63 - 0x3f
      10'h2D2: dout  = 8'b00111111; //  722 :  63 - 0x3f
      10'h2D3: dout  = 8'b00111111; //  723 :  63 - 0x3f
      10'h2D4: dout  = 8'b00111111; //  724 :  63 - 0x3f
      10'h2D5: dout  = 8'b00111111; //  725 :  63 - 0x3f
      10'h2D6: dout  = 8'b00111111; //  726 :  63 - 0x3f
      10'h2D7: dout  = 8'b00111111; //  727 :  63 - 0x3f
      10'h2D8: dout  = 8'b00111111; //  728 :  63 - 0x3f
      10'h2D9: dout  = 8'b00111111; //  729 :  63 - 0x3f
      10'h2DA: dout  = 8'b00111111; //  730 :  63 - 0x3f
      10'h2DB: dout  = 8'b00111111; //  731 :  63 - 0x3f
      10'h2DC: dout  = 8'b00111111; //  732 :  63 - 0x3f
      10'h2DD: dout  = 8'b00111111; //  733 :  63 - 0x3f
      10'h2DE: dout  = 8'b00111111; //  734 :  63 - 0x3f
      10'h2DF: dout  = 8'b00111111; //  735 :  63 - 0x3f
      10'h2E0: dout  = 8'b00111111; //  736 :  63 - 0x3f -- line 0x17
      10'h2E1: dout  = 8'b00111111; //  737 :  63 - 0x3f
      10'h2E2: dout  = 8'b00111111; //  738 :  63 - 0x3f
      10'h2E3: dout  = 8'b00111111; //  739 :  63 - 0x3f
      10'h2E4: dout  = 8'b00111111; //  740 :  63 - 0x3f
      10'h2E5: dout  = 8'b00111111; //  741 :  63 - 0x3f
      10'h2E6: dout  = 8'b00111111; //  742 :  63 - 0x3f
      10'h2E7: dout  = 8'b00111111; //  743 :  63 - 0x3f
      10'h2E8: dout  = 8'b00111111; //  744 :  63 - 0x3f
      10'h2E9: dout  = 8'b00111111; //  745 :  63 - 0x3f
      10'h2EA: dout  = 8'b00111111; //  746 :  63 - 0x3f
      10'h2EB: dout  = 8'b00111111; //  747 :  63 - 0x3f
      10'h2EC: dout  = 8'b00111111; //  748 :  63 - 0x3f
      10'h2ED: dout  = 8'b00111111; //  749 :  63 - 0x3f
      10'h2EE: dout  = 8'b00111111; //  750 :  63 - 0x3f
      10'h2EF: dout  = 8'b00111111; //  751 :  63 - 0x3f
      10'h2F0: dout  = 8'b11000101; //  752 : 197 - 0xc5
      10'h2F1: dout  = 8'b11010110; //  753 : 214 - 0xd6
      10'h2F2: dout  = 8'b11000101; //  754 : 197 - 0xc5
      10'h2F3: dout  = 8'b11010110; //  755 : 214 - 0xd6
      10'h2F4: dout  = 8'b11000101; //  756 : 197 - 0xc5
      10'h2F5: dout  = 8'b11010110; //  757 : 214 - 0xd6
      10'h2F6: dout  = 8'b11000101; //  758 : 197 - 0xc5
      10'h2F7: dout  = 8'b11010110; //  759 : 214 - 0xd6
      10'h2F8: dout  = 8'b11000101; //  760 : 197 - 0xc5
      10'h2F9: dout  = 8'b11010110; //  761 : 214 - 0xd6
      10'h2FA: dout  = 8'b11000101; //  762 : 197 - 0xc5
      10'h2FB: dout  = 8'b11010110; //  763 : 214 - 0xd6
      10'h2FC: dout  = 8'b11000101; //  764 : 197 - 0xc5
      10'h2FD: dout  = 8'b11010110; //  765 : 214 - 0xd6
      10'h2FE: dout  = 8'b11000101; //  766 : 197 - 0xc5
      10'h2FF: dout  = 8'b11010110; //  767 : 214 - 0xd6
      10'h300: dout  = 8'b00111111; //  768 :  63 - 0x3f -- line 0x18
      10'h301: dout  = 8'b00111111; //  769 :  63 - 0x3f
      10'h302: dout  = 8'b00111111; //  770 :  63 - 0x3f
      10'h303: dout  = 8'b00111111; //  771 :  63 - 0x3f
      10'h304: dout  = 8'b00011100; //  772 :  28 - 0x1c
      10'h305: dout  = 8'b00011110; //  773 :  30 - 0x1e
      10'h306: dout  = 8'b00111111; //  774 :  63 - 0x3f
      10'h307: dout  = 8'b00111111; //  775 :  63 - 0x3f
      10'h308: dout  = 8'b00111111; //  776 :  63 - 0x3f
      10'h309: dout  = 8'b00111111; //  777 :  63 - 0x3f
      10'h30A: dout  = 8'b00111111; //  778 :  63 - 0x3f
      10'h30B: dout  = 8'b00111111; //  779 :  63 - 0x3f
      10'h30C: dout  = 8'b00111111; //  780 :  63 - 0x3f
      10'h30D: dout  = 8'b00111111; //  781 :  63 - 0x3f
      10'h30E: dout  = 8'b00111111; //  782 :  63 - 0x3f
      10'h30F: dout  = 8'b00111111; //  783 :  63 - 0x3f
      10'h310: dout  = 8'b11000111; //  784 : 199 - 0xc7
      10'h311: dout  = 8'b11001001; //  785 : 201 - 0xc9
      10'h312: dout  = 8'b11000111; //  786 : 199 - 0xc7
      10'h313: dout  = 8'b11001001; //  787 : 201 - 0xc9
      10'h314: dout  = 8'b11000111; //  788 : 199 - 0xc7
      10'h315: dout  = 8'b11001001; //  789 : 201 - 0xc9
      10'h316: dout  = 8'b11000111; //  790 : 199 - 0xc7
      10'h317: dout  = 8'b11001001; //  791 : 201 - 0xc9
      10'h318: dout  = 8'b11000111; //  792 : 199 - 0xc7
      10'h319: dout  = 8'b11001001; //  793 : 201 - 0xc9
      10'h31A: dout  = 8'b11000111; //  794 : 199 - 0xc7
      10'h31B: dout  = 8'b11001001; //  795 : 201 - 0xc9
      10'h31C: dout  = 8'b11000111; //  796 : 199 - 0xc7
      10'h31D: dout  = 8'b11001001; //  797 : 201 - 0xc9
      10'h31E: dout  = 8'b11000111; //  798 : 199 - 0xc7
      10'h31F: dout  = 8'b11001001; //  799 : 201 - 0xc9
      10'h320: dout  = 8'b00111111; //  800 :  63 - 0x3f -- line 0x19
      10'h321: dout  = 8'b00111111; //  801 :  63 - 0x3f
      10'h322: dout  = 8'b00111111; //  802 :  63 - 0x3f
      10'h323: dout  = 8'b00111111; //  803 :  63 - 0x3f
      10'h324: dout  = 8'b00011101; //  804 :  29 - 0x1d
      10'h325: dout  = 8'b00011111; //  805 :  31 - 0x1f
      10'h326: dout  = 8'b00111111; //  806 :  63 - 0x3f
      10'h327: dout  = 8'b00111111; //  807 :  63 - 0x3f
      10'h328: dout  = 8'b00111111; //  808 :  63 - 0x3f
      10'h329: dout  = 8'b00111111; //  809 :  63 - 0x3f
      10'h32A: dout  = 8'b00111111; //  810 :  63 - 0x3f
      10'h32B: dout  = 8'b00111111; //  811 :  63 - 0x3f
      10'h32C: dout  = 8'b00111111; //  812 :  63 - 0x3f
      10'h32D: dout  = 8'b00111111; //  813 :  63 - 0x3f
      10'h32E: dout  = 8'b00111111; //  814 :  63 - 0x3f
      10'h32F: dout  = 8'b00111111; //  815 :  63 - 0x3f
      10'h330: dout  = 8'b11010111; //  816 : 215 - 0xd7
      10'h331: dout  = 8'b11011001; //  817 : 217 - 0xd9
      10'h332: dout  = 8'b11010111; //  818 : 215 - 0xd7
      10'h333: dout  = 8'b11011001; //  819 : 217 - 0xd9
      10'h334: dout  = 8'b11010111; //  820 : 215 - 0xd7
      10'h335: dout  = 8'b11011001; //  821 : 217 - 0xd9
      10'h336: dout  = 8'b11010111; //  822 : 215 - 0xd7
      10'h337: dout  = 8'b11011001; //  823 : 217 - 0xd9
      10'h338: dout  = 8'b11010111; //  824 : 215 - 0xd7
      10'h339: dout  = 8'b11011001; //  825 : 217 - 0xd9
      10'h33A: dout  = 8'b11010111; //  826 : 215 - 0xd7
      10'h33B: dout  = 8'b11011001; //  827 : 217 - 0xd9
      10'h33C: dout  = 8'b11010111; //  828 : 215 - 0xd7
      10'h33D: dout  = 8'b11011001; //  829 : 217 - 0xd9
      10'h33E: dout  = 8'b11010111; //  830 : 215 - 0xd7
      10'h33F: dout  = 8'b11011001; //  831 : 217 - 0xd9
      10'h340: dout  = 8'b01110000; //  832 : 112 - 0x70 -- line 0x1a
      10'h341: dout  = 8'b01110001; //  833 : 113 - 0x71
      10'h342: dout  = 8'b01110001; //  834 : 113 - 0x71
      10'h343: dout  = 8'b01110001; //  835 : 113 - 0x71
      10'h344: dout  = 8'b01110001; //  836 : 113 - 0x71
      10'h345: dout  = 8'b01110001; //  837 : 113 - 0x71
      10'h346: dout  = 8'b01110001; //  838 : 113 - 0x71
      10'h347: dout  = 8'b01110001; //  839 : 113 - 0x71
      10'h348: dout  = 8'b01110001; //  840 : 113 - 0x71
      10'h349: dout  = 8'b01110001; //  841 : 113 - 0x71
      10'h34A: dout  = 8'b01110001; //  842 : 113 - 0x71
      10'h34B: dout  = 8'b01110001; //  843 : 113 - 0x71
      10'h34C: dout  = 8'b01110001; //  844 : 113 - 0x71
      10'h34D: dout  = 8'b01110001; //  845 : 113 - 0x71
      10'h34E: dout  = 8'b01110001; //  846 : 113 - 0x71
      10'h34F: dout  = 8'b01110001; //  847 : 113 - 0x71
      10'h350: dout  = 8'b01110001; //  848 : 113 - 0x71
      10'h351: dout  = 8'b01110001; //  849 : 113 - 0x71
      10'h352: dout  = 8'b01110001; //  850 : 113 - 0x71
      10'h353: dout  = 8'b01110001; //  851 : 113 - 0x71
      10'h354: dout  = 8'b01110001; //  852 : 113 - 0x71
      10'h355: dout  = 8'b01110001; //  853 : 113 - 0x71
      10'h356: dout  = 8'b01110001; //  854 : 113 - 0x71
      10'h357: dout  = 8'b01110001; //  855 : 113 - 0x71
      10'h358: dout  = 8'b01110001; //  856 : 113 - 0x71
      10'h359: dout  = 8'b01110001; //  857 : 113 - 0x71
      10'h35A: dout  = 8'b01110001; //  858 : 113 - 0x71
      10'h35B: dout  = 8'b01110001; //  859 : 113 - 0x71
      10'h35C: dout  = 8'b01110001; //  860 : 113 - 0x71
      10'h35D: dout  = 8'b01110001; //  861 : 113 - 0x71
      10'h35E: dout  = 8'b01110001; //  862 : 113 - 0x71
      10'h35F: dout  = 8'b01110001; //  863 : 113 - 0x71
      10'h360: dout  = 8'b01100000; //  864 :  96 - 0x60 -- line 0x1b
      10'h361: dout  = 8'b01110111; //  865 : 119 - 0x77
      10'h362: dout  = 8'b01110111; //  866 : 119 - 0x77
      10'h363: dout  = 8'b01110111; //  867 : 119 - 0x77
      10'h364: dout  = 8'b01110111; //  868 : 119 - 0x77
      10'h365: dout  = 8'b01110111; //  869 : 119 - 0x77
      10'h366: dout  = 8'b01110111; //  870 : 119 - 0x77
      10'h367: dout  = 8'b01110111; //  871 : 119 - 0x77
      10'h368: dout  = 8'b01110111; //  872 : 119 - 0x77
      10'h369: dout  = 8'b01110111; //  873 : 119 - 0x77
      10'h36A: dout  = 8'b01110111; //  874 : 119 - 0x77
      10'h36B: dout  = 8'b01110111; //  875 : 119 - 0x77
      10'h36C: dout  = 8'b01110111; //  876 : 119 - 0x77
      10'h36D: dout  = 8'b01110111; //  877 : 119 - 0x77
      10'h36E: dout  = 8'b01110111; //  878 : 119 - 0x77
      10'h36F: dout  = 8'b01110111; //  879 : 119 - 0x77
      10'h370: dout  = 8'b01110111; //  880 : 119 - 0x77
      10'h371: dout  = 8'b01110111; //  881 : 119 - 0x77
      10'h372: dout  = 8'b01110111; //  882 : 119 - 0x77
      10'h373: dout  = 8'b01110111; //  883 : 119 - 0x77
      10'h374: dout  = 8'b01110111; //  884 : 119 - 0x77
      10'h375: dout  = 8'b01110111; //  885 : 119 - 0x77
      10'h376: dout  = 8'b01110111; //  886 : 119 - 0x77
      10'h377: dout  = 8'b01110111; //  887 : 119 - 0x77
      10'h378: dout  = 8'b01110111; //  888 : 119 - 0x77
      10'h379: dout  = 8'b01110111; //  889 : 119 - 0x77
      10'h37A: dout  = 8'b01110111; //  890 : 119 - 0x77
      10'h37B: dout  = 8'b01110111; //  891 : 119 - 0x77
      10'h37C: dout  = 8'b01110111; //  892 : 119 - 0x77
      10'h37D: dout  = 8'b01110111; //  893 : 119 - 0x77
      10'h37E: dout  = 8'b01110111; //  894 : 119 - 0x77
      10'h37F: dout  = 8'b01110111; //  895 : 119 - 0x77
      10'h380: dout  = 8'b01100000; //  896 :  96 - 0x60 -- line 0x1c
      10'h381: dout  = 8'b01110011; //  897 : 115 - 0x73
      10'h382: dout  = 8'b01110011; //  898 : 115 - 0x73
      10'h383: dout  = 8'b01110011; //  899 : 115 - 0x73
      10'h384: dout  = 8'b01110011; //  900 : 115 - 0x73
      10'h385: dout  = 8'b01110011; //  901 : 115 - 0x73
      10'h386: dout  = 8'b01110011; //  902 : 115 - 0x73
      10'h387: dout  = 8'b01110011; //  903 : 115 - 0x73
      10'h388: dout  = 8'b01110011; //  904 : 115 - 0x73
      10'h389: dout  = 8'b01110011; //  905 : 115 - 0x73
      10'h38A: dout  = 8'b01110011; //  906 : 115 - 0x73
      10'h38B: dout  = 8'b01110011; //  907 : 115 - 0x73
      10'h38C: dout  = 8'b01110011; //  908 : 115 - 0x73
      10'h38D: dout  = 8'b01110011; //  909 : 115 - 0x73
      10'h38E: dout  = 8'b01110011; //  910 : 115 - 0x73
      10'h38F: dout  = 8'b01110011; //  911 : 115 - 0x73
      10'h390: dout  = 8'b01110011; //  912 : 115 - 0x73
      10'h391: dout  = 8'b01110011; //  913 : 115 - 0x73
      10'h392: dout  = 8'b01110011; //  914 : 115 - 0x73
      10'h393: dout  = 8'b01110011; //  915 : 115 - 0x73
      10'h394: dout  = 8'b01110011; //  916 : 115 - 0x73
      10'h395: dout  = 8'b01110011; //  917 : 115 - 0x73
      10'h396: dout  = 8'b01110011; //  918 : 115 - 0x73
      10'h397: dout  = 8'b01110011; //  919 : 115 - 0x73
      10'h398: dout  = 8'b01110011; //  920 : 115 - 0x73
      10'h399: dout  = 8'b01110011; //  921 : 115 - 0x73
      10'h39A: dout  = 8'b01110011; //  922 : 115 - 0x73
      10'h39B: dout  = 8'b01110011; //  923 : 115 - 0x73
      10'h39C: dout  = 8'b01110011; //  924 : 115 - 0x73
      10'h39D: dout  = 8'b01110011; //  925 : 115 - 0x73
      10'h39E: dout  = 8'b01110011; //  926 : 115 - 0x73
      10'h39F: dout  = 8'b01110011; //  927 : 115 - 0x73
      10'h3A0: dout  = 8'b01100000; //  928 :  96 - 0x60 -- line 0x1d
      10'h3A1: dout  = 8'b01110011; //  929 : 115 - 0x73
      10'h3A2: dout  = 8'b01110011; //  930 : 115 - 0x73
      10'h3A3: dout  = 8'b01110011; //  931 : 115 - 0x73
      10'h3A4: dout  = 8'b01110011; //  932 : 115 - 0x73
      10'h3A5: dout  = 8'b01110011; //  933 : 115 - 0x73
      10'h3A6: dout  = 8'b01110011; //  934 : 115 - 0x73
      10'h3A7: dout  = 8'b01110011; //  935 : 115 - 0x73
      10'h3A8: dout  = 8'b01110011; //  936 : 115 - 0x73
      10'h3A9: dout  = 8'b01110011; //  937 : 115 - 0x73
      10'h3AA: dout  = 8'b01110011; //  938 : 115 - 0x73
      10'h3AB: dout  = 8'b01110011; //  939 : 115 - 0x73
      10'h3AC: dout  = 8'b01110011; //  940 : 115 - 0x73
      10'h3AD: dout  = 8'b01110011; //  941 : 115 - 0x73
      10'h3AE: dout  = 8'b01110011; //  942 : 115 - 0x73
      10'h3AF: dout  = 8'b01110011; //  943 : 115 - 0x73
      10'h3B0: dout  = 8'b01110011; //  944 : 115 - 0x73
      10'h3B1: dout  = 8'b01110011; //  945 : 115 - 0x73
      10'h3B2: dout  = 8'b01110011; //  946 : 115 - 0x73
      10'h3B3: dout  = 8'b01110011; //  947 : 115 - 0x73
      10'h3B4: dout  = 8'b01110011; //  948 : 115 - 0x73
      10'h3B5: dout  = 8'b01110011; //  949 : 115 - 0x73
      10'h3B6: dout  = 8'b01110011; //  950 : 115 - 0x73
      10'h3B7: dout  = 8'b01110011; //  951 : 115 - 0x73
      10'h3B8: dout  = 8'b01110011; //  952 : 115 - 0x73
      10'h3B9: dout  = 8'b01110011; //  953 : 115 - 0x73
      10'h3BA: dout  = 8'b01110011; //  954 : 115 - 0x73
      10'h3BB: dout  = 8'b01110011; //  955 : 115 - 0x73
      10'h3BC: dout  = 8'b01110011; //  956 : 115 - 0x73
      10'h3BD: dout  = 8'b01110011; //  957 : 115 - 0x73
      10'h3BE: dout  = 8'b01110011; //  958 : 115 - 0x73
      10'h3BF: dout  = 8'b01110011; //  959 : 115 - 0x73
        //-- Attribute Table 0----
      10'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0
      10'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      10'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      10'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      10'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      10'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      10'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      10'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      10'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      10'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      10'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      10'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      10'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      10'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      10'h3CE: dout  = 8'b00001000; //  974 :   8 - 0x8
      10'h3CF: dout  = 8'b00001000; //  975 :   8 - 0x8
      10'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0
      10'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      10'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      10'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      10'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      10'h3D5: dout  = 8'b01010001; //  981 :  81 - 0x51
      10'h3D6: dout  = 8'b01010000; //  982 :  80 - 0x50
      10'h3D7: dout  = 8'b01010000; //  983 :  80 - 0x50
      10'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0
      10'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      10'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      10'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      10'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      10'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      10'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      10'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      10'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0
      10'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      10'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      10'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      10'h3E4: dout  = 8'b10100000; //  996 : 160 - 0xa0
      10'h3E5: dout  = 8'b10100000; //  997 : 160 - 0xa0
      10'h3E6: dout  = 8'b10100000; //  998 : 160 - 0xa0
      10'h3E7: dout  = 8'b10100000; //  999 : 160 - 0xa0
      10'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      10'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      10'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      10'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      10'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      10'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      10'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      10'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      10'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0
      10'h3F1: dout  = 8'b00000010; // 1009 :   2 - 0x2
      10'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      10'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      10'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      10'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      10'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      10'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      10'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0
      10'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      10'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      10'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      10'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      10'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      10'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      10'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
    endcase
  end

endmodule
