--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN_color1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN_color1;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN_color1 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Sprite 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Sprite 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Sprite 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Sprite 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x11
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x12
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- Sprite 0x15
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Sprite 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000011", --  194 - 0xc2  :    3 - 0x3
    "00000011", --  195 - 0xc3  :    3 - 0x3
    "00010011", --  196 - 0xc4  :   19 - 0x13
    "00111111", --  197 - 0xc5  :   63 - 0x3f
    "00111111", --  198 - 0xc6  :   63 - 0x3f
    "01111111", --  199 - 0xc7  :  127 - 0x7f
    "01111111", --  200 - 0xc8  :  127 - 0x7f -- Sprite 0x19
    "01111111", --  201 - 0xc9  :  127 - 0x7f
    "01111111", --  202 - 0xca  :  127 - 0x7f
    "01111111", --  203 - 0xcb  :  127 - 0x7f
    "01101110", --  204 - 0xcc  :  110 - 0x6e
    "01000110", --  205 - 0xcd  :   70 - 0x46
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "01111111", --  208 - 0xd0  :  127 - 0x7f -- Sprite 0x1a
    "01111111", --  209 - 0xd1  :  127 - 0x7f
    "01111111", --  210 - 0xd2  :  127 - 0x7f
    "01111111", --  211 - 0xd3  :  127 - 0x7f
    "01111011", --  212 - 0xd4  :  123 - 0x7b
    "00110001", --  213 - 0xd5  :   49 - 0x31
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "00000011", --  217 - 0xd9  :    3 - 0x3
    "00001111", --  218 - 0xda  :   15 - 0xf
    "00011111", --  219 - 0xdb  :   31 - 0x1f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00111111", --  221 - 0xdd  :   63 - 0x3f
    "00001111", --  222 - 0xde  :   15 - 0xf
    "01001111", --  223 - 0xdf  :   79 - 0x4f
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0x1c
    "11000000", --  225 - 0xe1  :  192 - 0xc0
    "11110000", --  226 - 0xe2  :  240 - 0xf0
    "11111000", --  227 - 0xe3  :  248 - 0xf8
    "11111100", --  228 - 0xe4  :  252 - 0xfc
    "11111100", --  229 - 0xe5  :  252 - 0xfc
    "00111100", --  230 - 0xe6  :   60 - 0x3c
    "00111110", --  231 - 0xe7  :   62 - 0x3e
    "01111111", --  232 - 0xe8  :  127 - 0x7f -- Sprite 0x1d
    "01111111", --  233 - 0xe9  :  127 - 0x7f
    "01111111", --  234 - 0xea  :  127 - 0x7f
    "01111111", --  235 - 0xeb  :  127 - 0x7f
    "01101110", --  236 - 0xec  :  110 - 0x6e
    "01000110", --  237 - 0xed  :   70 - 0x46
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "01111111", --  240 - 0xf0  :  127 - 0x7f -- Sprite 0x1e
    "01111111", --  241 - 0xf1  :  127 - 0x7f
    "01111111", --  242 - 0xf2  :  127 - 0x7f
    "01111111", --  243 - 0xf3  :  127 - 0x7f
    "01111011", --  244 - 0xf4  :  123 - 0x7b
    "00110001", --  245 - 0xf5  :   49 - 0x31
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "11111110", --  248 - 0xf8  :  254 - 0xfe -- Sprite 0x1f
    "11111110", --  249 - 0xf9  :  254 - 0xfe
    "11111110", --  250 - 0xfa  :  254 - 0xfe
    "11111110", --  251 - 0xfb  :  254 - 0xfe
    "01110110", --  252 - 0xfc  :  118 - 0x76
    "01100010", --  253 - 0xfd  :   98 - 0x62
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "11111110", --  256 - 0x100  :  254 - 0xfe -- Sprite 0x20
    "11111110", --  257 - 0x101  :  254 - 0xfe
    "11111110", --  258 - 0x102  :  254 - 0xfe
    "11111110", --  259 - 0x103  :  254 - 0xfe
    "11011110", --  260 - 0x104  :  222 - 0xde
    "10001100", --  261 - 0x105  :  140 - 0x8c
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000011", --  265 - 0x109  :    3 - 0x3
    "00001111", --  266 - 0x10a  :   15 - 0xf
    "00011111", --  267 - 0x10b  :   31 - 0x1f
    "00111111", --  268 - 0x10c  :   63 - 0x3f
    "00111111", --  269 - 0x10d  :   63 - 0x3f
    "00111111", --  270 - 0x10e  :   63 - 0x3f
    "01111111", --  271 - 0x10f  :  127 - 0x7f
    "01110011", --  272 - 0x110  :  115 - 0x73 -- Sprite 0x22
    "01110011", --  273 - 0x111  :  115 - 0x73
    "01111111", --  274 - 0x112  :  127 - 0x7f
    "01111111", --  275 - 0x113  :  127 - 0x7f
    "01101110", --  276 - 0x114  :  110 - 0x6e
    "01000110", --  277 - 0x115  :   70 - 0x46
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "01110011", --  280 - 0x118  :  115 - 0x73 -- Sprite 0x23
    "01110011", --  281 - 0x119  :  115 - 0x73
    "01111111", --  282 - 0x11a  :  127 - 0x7f
    "01111111", --  283 - 0x11b  :  127 - 0x7f
    "01110111", --  284 - 0x11c  :  119 - 0x77
    "00100011", --  285 - 0x11d  :   35 - 0x23
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000110", --  293 - 0x125  :    6 - 0x6
    "00000110", --  294 - 0x126  :    6 - 0x6
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- Sprite 0x25
    "00011001", --  297 - 0x129  :   25 - 0x19
    "00100110", --  298 - 0x12a  :   38 - 0x26
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "00011001", --  305 - 0x131  :   25 - 0x19
    "00100110", --  306 - 0x132  :   38 - 0x26
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Sprite 0x27
    "00001100", --  313 - 0x139  :   12 - 0xc
    "00010010", --  314 - 0x13a  :   18 - 0x12
    "00010010", --  315 - 0x13b  :   18 - 0x12
    "00011110", --  316 - 0x13c  :   30 - 0x1e
    "00001100", --  317 - 0x13d  :   12 - 0xc
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00111000", --  325 - 0x145  :   56 - 0x38
    "01001101", --  326 - 0x146  :   77 - 0x4d
    "01001101", --  327 - 0x147  :   77 - 0x4d
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Sprite 0x29
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "11100000", --  333 - 0x14d  :  224 - 0xe0
    "00110000", --  334 - 0x14e  :   48 - 0x30
    "00110000", --  335 - 0x14f  :   48 - 0x30
    "00111000", --  336 - 0x150  :   56 - 0x38 -- Sprite 0x2a
    "00000000", --  337 - 0x151  :    0 - 0x0
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "11100000", --  344 - 0x158  :  224 - 0xe0 -- Sprite 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00001100", --  358 - 0x166  :   12 - 0xc
    "00011110", --  359 - 0x167  :   30 - 0x1e
    "00010010", --  360 - 0x168  :   18 - 0x12 -- Sprite 0x2d
    "00010010", --  361 - 0x169  :   18 - 0x12
    "00001100", --  362 - 0x16a  :   12 - 0xc
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00010001", --  371 - 0x173  :   17 - 0x11
    "00110010", --  372 - 0x174  :   50 - 0x32
    "00010010", --  373 - 0x175  :   18 - 0x12
    "00010010", --  374 - 0x176  :   18 - 0x12
    "00010010", --  375 - 0x177  :   18 - 0x12
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "10001100", --  379 - 0x17b  :  140 - 0x8c
    "01010010", --  380 - 0x17c  :   82 - 0x52
    "01010010", --  381 - 0x17d  :   82 - 0x52
    "01010010", --  382 - 0x17e  :   82 - 0x52
    "01010010", --  383 - 0x17f  :   82 - 0x52
    "00010010", --  384 - 0x180  :   18 - 0x12 -- Sprite 0x30
    "00111001", --  385 - 0x181  :   57 - 0x39
    "00000000", --  386 - 0x182  :    0 - 0x0
    "00000000", --  387 - 0x183  :    0 - 0x0
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00000000", --  389 - 0x185  :    0 - 0x0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "01010010", --  392 - 0x188  :   82 - 0x52 -- Sprite 0x31
    "10001100", --  393 - 0x189  :  140 - 0x8c
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "01110001", --  403 - 0x193  :  113 - 0x71
    "10001010", --  404 - 0x194  :  138 - 0x8a
    "00001010", --  405 - 0x195  :   10 - 0xa
    "00010010", --  406 - 0x196  :   18 - 0x12
    "00100010", --  407 - 0x197  :   34 - 0x22
    "01000010", --  408 - 0x198  :   66 - 0x42 -- Sprite 0x33
    "11111001", --  409 - 0x199  :  249 - 0xf9
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00110001", --  419 - 0x1a3  :   49 - 0x31
    "01001010", --  420 - 0x1a4  :   74 - 0x4a
    "00001010", --  421 - 0x1a5  :   10 - 0xa
    "00110010", --  422 - 0x1a6  :   50 - 0x32
    "00001010", --  423 - 0x1a7  :   10 - 0xa
    "01001010", --  424 - 0x1a8  :   74 - 0x4a -- Sprite 0x35
    "00110001", --  425 - 0x1a9  :   49 - 0x31
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00010001", --  435 - 0x1b3  :   17 - 0x11
    "00110010", --  436 - 0x1b4  :   50 - 0x32
    "01010010", --  437 - 0x1b5  :   82 - 0x52
    "10010010", --  438 - 0x1b6  :  146 - 0x92
    "11111010", --  439 - 0x1b7  :  250 - 0xfa
    "00010010", --  440 - 0x1b8  :   18 - 0x12 -- Sprite 0x37
    "00010001", --  441 - 0x1b9  :   17 - 0x11
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "01110001", --  451 - 0x1c3  :  113 - 0x71
    "01000010", --  452 - 0x1c4  :   66 - 0x42
    "01000010", --  453 - 0x1c5  :   66 - 0x42
    "01110010", --  454 - 0x1c6  :  114 - 0x72
    "00001010", --  455 - 0x1c7  :   10 - 0xa
    "00001010", --  456 - 0x1c8  :   10 - 0xa -- Sprite 0x39
    "01110001", --  457 - 0x1c9  :  113 - 0x71
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "01110001", --  467 - 0x1d3  :  113 - 0x71
    "00001010", --  468 - 0x1d4  :   10 - 0xa
    "00010010", --  469 - 0x1d5  :   18 - 0x12
    "00010010", --  470 - 0x1d6  :   18 - 0x12
    "00100010", --  471 - 0x1d7  :   34 - 0x22
    "00100010", --  472 - 0x1d8  :   34 - 0x22 -- Sprite 0x3b
    "00100001", --  473 - 0x1d9  :   33 - 0x21
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "01110001", --  483 - 0x1e3  :  113 - 0x71
    "10001010", --  484 - 0x1e4  :  138 - 0x8a
    "10001010", --  485 - 0x1e5  :  138 - 0x8a
    "01110010", --  486 - 0x1e6  :  114 - 0x72
    "10001010", --  487 - 0x1e7  :  138 - 0x8a
    "10001010", --  488 - 0x1e8  :  138 - 0x8a -- Sprite 0x3d
    "01110001", --  489 - 0x1e9  :  113 - 0x71
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "10011000", --  499 - 0x1f3  :  152 - 0x98
    "10100101", --  500 - 0x1f4  :  165 - 0xa5
    "10100101", --  501 - 0x1f5  :  165 - 0xa5
    "10100101", --  502 - 0x1f6  :  165 - 0xa5
    "10100101", --  503 - 0x1f7  :  165 - 0xa5
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "11000110", --  507 - 0x1fb  :  198 - 0xc6
    "00101001", --  508 - 0x1fc  :   41 - 0x29
    "00101001", --  509 - 0x1fd  :   41 - 0x29
    "00101001", --  510 - 0x1fe  :   41 - 0x29
    "00101001", --  511 - 0x1ff  :   41 - 0x29
    "10100101", --  512 - 0x200  :  165 - 0xa5 -- Sprite 0x40
    "10011000", --  513 - 0x201  :  152 - 0x98
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00101001", --  520 - 0x208  :   41 - 0x29 -- Sprite 0x41
    "11000110", --  521 - 0x209  :  198 - 0xc6
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Sprite 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "10011100", --  531 - 0x213  :  156 - 0x9c
    "10100001", --  532 - 0x214  :  161 - 0xa1
    "10100001", --  533 - 0x215  :  161 - 0xa1
    "10111101", --  534 - 0x216  :  189 - 0xbd
    "10100101", --  535 - 0x217  :  165 - 0xa5
    "10100101", --  536 - 0x218  :  165 - 0xa5 -- Sprite 0x43
    "10011000", --  537 - 0x219  :  152 - 0x98
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Sprite 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "01100010", --  547 - 0x223  :   98 - 0x62
    "10010101", --  548 - 0x224  :  149 - 0x95
    "00010101", --  549 - 0x225  :   21 - 0x15
    "00100101", --  550 - 0x226  :   37 - 0x25
    "01000101", --  551 - 0x227  :   69 - 0x45
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Sprite 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00100010", --  555 - 0x22b  :   34 - 0x22
    "01010101", --  556 - 0x22c  :   85 - 0x55
    "01010101", --  557 - 0x22d  :   85 - 0x55
    "01010101", --  558 - 0x22e  :   85 - 0x55
    "01010101", --  559 - 0x22f  :   85 - 0x55
    "10000101", --  560 - 0x230  :  133 - 0x85 -- Sprite 0x46
    "11110010", --  561 - 0x231  :  242 - 0xf2
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "01010101", --  568 - 0x238  :   85 - 0x55 -- Sprite 0x47
    "00100010", --  569 - 0x239  :   34 - 0x22
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "01100010", --  579 - 0x243  :   98 - 0x62
    "10010101", --  580 - 0x244  :  149 - 0x95
    "00010101", --  581 - 0x245  :   21 - 0x15
    "01100101", --  582 - 0x246  :  101 - 0x65
    "00010101", --  583 - 0x247  :   21 - 0x15
    "10010101", --  584 - 0x248  :  149 - 0x95 -- Sprite 0x49
    "01100010", --  585 - 0x249  :   98 - 0x62
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Sprite 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "11100010", --  595 - 0x253  :  226 - 0xe2
    "10000101", --  596 - 0x254  :  133 - 0x85
    "10000101", --  597 - 0x255  :  133 - 0x85
    "11100101", --  598 - 0x256  :  229 - 0xe5
    "00010101", --  599 - 0x257  :   21 - 0x15
    "00010101", --  600 - 0x258  :   21 - 0x15 -- Sprite 0x4b
    "11100010", --  601 - 0x259  :  226 - 0xe2
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Sprite 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Sprite 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Sprite 0x56
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Sprite 0x57
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000100", --  703 - 0x2bf  :    4 - 0x4
    "00000110", --  704 - 0x2c0  :    6 - 0x6 -- Sprite 0x58
    "00000110", --  705 - 0x2c1  :    6 - 0x6
    "00000111", --  706 - 0x2c2  :    7 - 0x7
    "00000111", --  707 - 0x2c3  :    7 - 0x7
    "00000111", --  708 - 0x2c4  :    7 - 0x7
    "00000111", --  709 - 0x2c5  :    7 - 0x7
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Sprite 0x59
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00010000", --  719 - 0x2cf  :   16 - 0x10
    "00011100", --  720 - 0x2d0  :   28 - 0x1c -- Sprite 0x5a
    "00011110", --  721 - 0x2d1  :   30 - 0x1e
    "00011111", --  722 - 0x2d2  :   31 - 0x1f
    "00011111", --  723 - 0x2d3  :   31 - 0x1f
    "00011111", --  724 - 0x2d4  :   31 - 0x1f
    "00011111", --  725 - 0x2d5  :   31 - 0x1f
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "11000000", --  735 - 0x2df  :  192 - 0xc0
    "11110000", --  736 - 0x2e0  :  240 - 0xf0 -- Sprite 0x5c
    "11111100", --  737 - 0x2e1  :  252 - 0xfc
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Sprite 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000001", --  746 - 0x2ea  :    1 - 0x1
    "00000011", --  747 - 0x2eb  :    3 - 0x3
    "00001111", --  748 - 0x2ec  :   15 - 0xf
    "00001111", --  749 - 0x2ed  :   15 - 0xf
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "11111000", --  752 - 0x2f0  :  248 - 0xf8 -- Sprite 0x5e
    "11110000", --  753 - 0x2f1  :  240 - 0xf0
    "11100000", --  754 - 0x2f2  :  224 - 0xe0
    "11110000", --  755 - 0x2f3  :  240 - 0xf0
    "11100000", --  756 - 0x2f4  :  224 - 0xe0
    "11000000", --  757 - 0x2f5  :  192 - 0xc0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Sprite 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00000011", --  769 - 0x301  :    3 - 0x3
    "00001111", --  770 - 0x302  :   15 - 0xf
    "00011111", --  771 - 0x303  :   31 - 0x1f
    "00111111", --  772 - 0x304  :   63 - 0x3f
    "00111111", --  773 - 0x305  :   63 - 0x3f
    "00111001", --  774 - 0x306  :   57 - 0x39
    "01111011", --  775 - 0x307  :  123 - 0x7b
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "11000000", --  777 - 0x309  :  192 - 0xc0
    "11110000", --  778 - 0x30a  :  240 - 0xf0
    "11111000", --  779 - 0x30b  :  248 - 0xf8
    "11111100", --  780 - 0x30c  :  252 - 0xfc
    "11111100", --  781 - 0x30d  :  252 - 0xfc
    "11100100", --  782 - 0x30e  :  228 - 0xe4
    "11101110", --  783 - 0x30f  :  238 - 0xee
    "11111110", --  784 - 0x310  :  254 - 0xfe -- Sprite 0x62
    "11111110", --  785 - 0x311  :  254 - 0xfe
    "11111110", --  786 - 0x312  :  254 - 0xfe
    "11111110", --  787 - 0x313  :  254 - 0xfe
    "11111110", --  788 - 0x314  :  254 - 0xfe
    "01100110", --  789 - 0x315  :  102 - 0x66
    "01000010", --  790 - 0x316  :   66 - 0x42
    "00000000", --  791 - 0x317  :    0 - 0x0
    "11111110", --  792 - 0x318  :  254 - 0xfe -- Sprite 0x63
    "11111110", --  793 - 0x319  :  254 - 0xfe
    "11111110", --  794 - 0x31a  :  254 - 0xfe
    "11111110", --  795 - 0x31b  :  254 - 0xfe
    "11111110", --  796 - 0x31c  :  254 - 0xfe
    "11011110", --  797 - 0x31d  :  222 - 0xde
    "10001100", --  798 - 0x31e  :  140 - 0x8c
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Sprite 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "01101100", --  812 - 0x32c  :  108 - 0x6c
    "11111110", --  813 - 0x32d  :  254 - 0xfe
    "11111110", --  814 - 0x32e  :  254 - 0xfe
    "11111100", --  815 - 0x32f  :  252 - 0xfc
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Sprite 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00011111", --  849 - 0x351  :   31 - 0x1f
    "01111111", --  850 - 0x352  :  127 - 0x7f
    "00111111", --  851 - 0x353  :   63 - 0x3f
    "00001111", --  852 - 0x354  :   15 - 0xf
    "00000111", --  853 - 0x355  :    7 - 0x7
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "11000000", --  858 - 0x35a  :  192 - 0xc0
    "11110000", --  859 - 0x35b  :  240 - 0xf0
    "11111000", --  860 - 0x35c  :  248 - 0xf8
    "11111000", --  861 - 0x35d  :  248 - 0xf8
    "11100000", --  862 - 0x35e  :  224 - 0xe0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "00000000", --  868 - 0x364  :    0 - 0x0
    "00000000", --  869 - 0x365  :    0 - 0x0
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00000000", --  888 - 0x378  :    0 - 0x0 -- Sprite 0x6f
    "00000000", --  889 - 0x379  :    0 - 0x0
    "00000000", --  890 - 0x37a  :    0 - 0x0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "11111111", --  896 - 0x380  :  255 - 0xff -- Sprite 0x70
    "11111111", --  897 - 0x381  :  255 - 0xff
    "11111111", --  898 - 0x382  :  255 - 0xff
    "11111111", --  899 - 0x383  :  255 - 0xff
    "11111111", --  900 - 0x384  :  255 - 0xff
    "11111111", --  901 - 0x385  :  255 - 0xff
    "11111111", --  902 - 0x386  :  255 - 0xff
    "11111111", --  903 - 0x387  :  255 - 0xff
    "11111111", --  904 - 0x388  :  255 - 0xff -- Sprite 0x71
    "11111111", --  905 - 0x389  :  255 - 0xff
    "11111111", --  906 - 0x38a  :  255 - 0xff
    "11111111", --  907 - 0x38b  :  255 - 0xff
    "11111111", --  908 - 0x38c  :  255 - 0xff
    "11111111", --  909 - 0x38d  :  255 - 0xff
    "11111111", --  910 - 0x38e  :  255 - 0xff
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "11111111", --  912 - 0x390  :  255 - 0xff -- Sprite 0x72
    "11111111", --  913 - 0x391  :  255 - 0xff
    "11111111", --  914 - 0x392  :  255 - 0xff
    "11111111", --  915 - 0x393  :  255 - 0xff
    "11111111", --  916 - 0x394  :  255 - 0xff
    "11111111", --  917 - 0x395  :  255 - 0xff
    "11111111", --  918 - 0x396  :  255 - 0xff
    "11111111", --  919 - 0x397  :  255 - 0xff
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111111", --  927 - 0x39f  :  255 - 0xff
    "11111111", --  928 - 0x3a0  :  255 - 0xff -- Sprite 0x74
    "11111111", --  929 - 0x3a1  :  255 - 0xff
    "11111111", --  930 - 0x3a2  :  255 - 0xff
    "11111111", --  931 - 0x3a3  :  255 - 0xff
    "11111111", --  932 - 0x3a4  :  255 - 0xff
    "11111111", --  933 - 0x3a5  :  255 - 0xff
    "11111111", --  934 - 0x3a6  :  255 - 0xff
    "11111111", --  935 - 0x3a7  :  255 - 0xff
    "11111111", --  936 - 0x3a8  :  255 - 0xff -- Sprite 0x75
    "11111111", --  937 - 0x3a9  :  255 - 0xff
    "11111111", --  938 - 0x3aa  :  255 - 0xff
    "11111111", --  939 - 0x3ab  :  255 - 0xff
    "11111111", --  940 - 0x3ac  :  255 - 0xff
    "11111111", --  941 - 0x3ad  :  255 - 0xff
    "11111111", --  942 - 0x3ae  :  255 - 0xff
    "11111111", --  943 - 0x3af  :  255 - 0xff
    "11111111", --  944 - 0x3b0  :  255 - 0xff -- Sprite 0x76
    "11111111", --  945 - 0x3b1  :  255 - 0xff
    "11111111", --  946 - 0x3b2  :  255 - 0xff
    "11111111", --  947 - 0x3b3  :  255 - 0xff
    "11111111", --  948 - 0x3b4  :  255 - 0xff
    "11111111", --  949 - 0x3b5  :  255 - 0xff
    "11111111", --  950 - 0x3b6  :  255 - 0xff
    "11111111", --  951 - 0x3b7  :  255 - 0xff
    "11111111", --  952 - 0x3b8  :  255 - 0xff -- Sprite 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111111", --  954 - 0x3ba  :  255 - 0xff
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "11111111", --  956 - 0x3bc  :  255 - 0xff
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Sprite 0x78
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "11111111", --  966 - 0x3c6  :  255 - 0xff
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Sprite 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "11111111", --  971 - 0x3cb  :  255 - 0xff
    "11111111", --  972 - 0x3cc  :  255 - 0xff
    "11111111", --  973 - 0x3cd  :  255 - 0xff
    "11111111", --  974 - 0x3ce  :  255 - 0xff
    "11111111", --  975 - 0x3cf  :  255 - 0xff
    "11111111", --  976 - 0x3d0  :  255 - 0xff -- Sprite 0x7a
    "11111111", --  977 - 0x3d1  :  255 - 0xff
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "11111111", --  980 - 0x3d4  :  255 - 0xff
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "11111111", --  982 - 0x3d6  :  255 - 0xff
    "11111111", --  983 - 0x3d7  :  255 - 0xff
    "11111111", --  984 - 0x3d8  :  255 - 0xff -- Sprite 0x7b
    "11111111", --  985 - 0x3d9  :  255 - 0xff
    "11111111", --  986 - 0x3da  :  255 - 0xff
    "11111111", --  987 - 0x3db  :  255 - 0xff
    "11111111", --  988 - 0x3dc  :  255 - 0xff
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "11111111", --  991 - 0x3df  :  255 - 0xff
    "11111111", --  992 - 0x3e0  :  255 - 0xff -- Sprite 0x7c
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111111", --  996 - 0x3e4  :  255 - 0xff
    "11111111", --  997 - 0x3e5  :  255 - 0xff
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "11111111", -- 1000 - 0x3e8  :  255 - 0xff -- Sprite 0x7d
    "11111111", -- 1001 - 0x3e9  :  255 - 0xff
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111111", -- 1004 - 0x3ec  :  255 - 0xff
    "11111111", -- 1005 - 0x3ed  :  255 - 0xff
    "11111111", -- 1006 - 0x3ee  :  255 - 0xff
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "11111111", -- 1008 - 0x3f0  :  255 - 0xff -- Sprite 0x7e
    "11111111", -- 1009 - 0x3f1  :  255 - 0xff
    "11111111", -- 1010 - 0x3f2  :  255 - 0xff
    "11111111", -- 1011 - 0x3f3  :  255 - 0xff
    "11111111", -- 1012 - 0x3f4  :  255 - 0xff
    "11111111", -- 1013 - 0x3f5  :  255 - 0xff
    "11111111", -- 1014 - 0x3f6  :  255 - 0xff
    "11111111", -- 1015 - 0x3f7  :  255 - 0xff
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Sprite 0x7f
    "11111111", -- 1017 - 0x3f9  :  255 - 0xff
    "11111111", -- 1018 - 0x3fa  :  255 - 0xff
    "11111111", -- 1019 - 0x3fb  :  255 - 0xff
    "11111111", -- 1020 - 0x3fc  :  255 - 0xff
    "11111111", -- 1021 - 0x3fd  :  255 - 0xff
    "11111111", -- 1022 - 0x3fe  :  255 - 0xff
    "11111111", -- 1023 - 0x3ff  :  255 - 0xff
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Sprite 0x80
    "11111111", -- 1025 - 0x401  :  255 - 0xff
    "11111111", -- 1026 - 0x402  :  255 - 0xff
    "11111111", -- 1027 - 0x403  :  255 - 0xff
    "11111111", -- 1028 - 0x404  :  255 - 0xff
    "11111111", -- 1029 - 0x405  :  255 - 0xff
    "11111111", -- 1030 - 0x406  :  255 - 0xff
    "11111111", -- 1031 - 0x407  :  255 - 0xff
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Sprite 0x81
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11111111", -- 1035 - 0x40b  :  255 - 0xff
    "11111111", -- 1036 - 0x40c  :  255 - 0xff
    "11111111", -- 1037 - 0x40d  :  255 - 0xff
    "11111111", -- 1038 - 0x40e  :  255 - 0xff
    "11111111", -- 1039 - 0x40f  :  255 - 0xff
    "11111111", -- 1040 - 0x410  :  255 - 0xff -- Sprite 0x82
    "11111111", -- 1041 - 0x411  :  255 - 0xff
    "11111111", -- 1042 - 0x412  :  255 - 0xff
    "11111111", -- 1043 - 0x413  :  255 - 0xff
    "11111111", -- 1044 - 0x414  :  255 - 0xff
    "11111111", -- 1045 - 0x415  :  255 - 0xff
    "11111111", -- 1046 - 0x416  :  255 - 0xff
    "11111111", -- 1047 - 0x417  :  255 - 0xff
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- Sprite 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "11111111", -- 1051 - 0x41b  :  255 - 0xff
    "11111111", -- 1052 - 0x41c  :  255 - 0xff
    "11111111", -- 1053 - 0x41d  :  255 - 0xff
    "11111111", -- 1054 - 0x41e  :  255 - 0xff
    "11111111", -- 1055 - 0x41f  :  255 - 0xff
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Sprite 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111111", -- 1061 - 0x425  :  255 - 0xff
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111111", -- 1067 - 0x42b  :  255 - 0xff
    "11111111", -- 1068 - 0x42c  :  255 - 0xff
    "11111111", -- 1069 - 0x42d  :  255 - 0xff
    "11111111", -- 1070 - 0x42e  :  255 - 0xff
    "11111111", -- 1071 - 0x42f  :  255 - 0xff
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "11111111", -- 1076 - 0x434  :  255 - 0xff
    "11111111", -- 1077 - 0x435  :  255 - 0xff
    "11111111", -- 1078 - 0x436  :  255 - 0xff
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "11111111", -- 1080 - 0x438  :  255 - 0xff -- Sprite 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "11111111", -- 1086 - 0x43e  :  255 - 0xff
    "11111111", -- 1087 - 0x43f  :  255 - 0xff
    "11111111", -- 1088 - 0x440  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "11111111", -- 1090 - 0x442  :  255 - 0xff
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- Sprite 0x89
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11111111", -- 1100 - 0x44c  :  255 - 0xff
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "11111111", -- 1104 - 0x450  :  255 - 0xff -- Sprite 0x8a
    "11111111", -- 1105 - 0x451  :  255 - 0xff
    "11111111", -- 1106 - 0x452  :  255 - 0xff
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "11111111", -- 1108 - 0x454  :  255 - 0xff
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- Sprite 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "11111111", -- 1117 - 0x45d  :  255 - 0xff
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11111111", -- 1119 - 0x45f  :  255 - 0xff
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Sprite 0x8c
    "11111111", -- 1121 - 0x461  :  255 - 0xff
    "11111111", -- 1122 - 0x462  :  255 - 0xff
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "11111111", -- 1125 - 0x465  :  255 - 0xff
    "11111111", -- 1126 - 0x466  :  255 - 0xff
    "11111111", -- 1127 - 0x467  :  255 - 0xff
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- Sprite 0x8d
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "11111111", -- 1130 - 0x46a  :  255 - 0xff
    "11111111", -- 1131 - 0x46b  :  255 - 0xff
    "11111111", -- 1132 - 0x46c  :  255 - 0xff
    "11111111", -- 1133 - 0x46d  :  255 - 0xff
    "11111111", -- 1134 - 0x46e  :  255 - 0xff
    "11111111", -- 1135 - 0x46f  :  255 - 0xff
    "11111111", -- 1136 - 0x470  :  255 - 0xff -- Sprite 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111111", -- 1138 - 0x472  :  255 - 0xff
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11111111", -- 1140 - 0x474  :  255 - 0xff
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- Sprite 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111111", -- 1146 - 0x47a  :  255 - 0xff
    "11111111", -- 1147 - 0x47b  :  255 - 0xff
    "11111111", -- 1148 - 0x47c  :  255 - 0xff
    "11111111", -- 1149 - 0x47d  :  255 - 0xff
    "11111111", -- 1150 - 0x47e  :  255 - 0xff
    "11111111", -- 1151 - 0x47f  :  255 - 0xff
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- Sprite 0x91
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0 -- Sprite 0x92
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- Sprite 0x93
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0 -- Sprite 0x95
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- Sprite 0x97
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x98
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- Sprite 0x99
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- Sprite 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Sprite 0x9c
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- Sprite 0x9d
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x9e
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000000", -- 1269 - 0x4f5  :    0 - 0x0
    "00000000", -- 1270 - 0x4f6  :    0 - 0x0
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0xa0
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- Sprite 0xa1
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0 -- Sprite 0xa2
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- Sprite 0xa3
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0xa4
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00000000", -- 1317 - 0x525  :    0 - 0x0
    "00000000", -- 1318 - 0x526  :    0 - 0x0
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0 -- Sprite 0xa7
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0 -- Sprite 0xa9
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Sprite 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Sprite 0xad
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "01111110", -- 1408 - 0x580  :  126 - 0x7e -- Sprite 0xb0
    "01100011", -- 1409 - 0x581  :   99 - 0x63
    "01100011", -- 1410 - 0x582  :   99 - 0x63
    "01100011", -- 1411 - 0x583  :   99 - 0x63
    "01111110", -- 1412 - 0x584  :  126 - 0x7e
    "01100000", -- 1413 - 0x585  :   96 - 0x60
    "01100000", -- 1414 - 0x586  :   96 - 0x60
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "01100000", -- 1416 - 0x588  :   96 - 0x60 -- Sprite 0xb1
    "01100000", -- 1417 - 0x589  :   96 - 0x60
    "01100000", -- 1418 - 0x58a  :   96 - 0x60
    "01100000", -- 1419 - 0x58b  :   96 - 0x60
    "01100000", -- 1420 - 0x58c  :   96 - 0x60
    "01100000", -- 1421 - 0x58d  :   96 - 0x60
    "01111111", -- 1422 - 0x58e  :  127 - 0x7f
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00011100", -- 1424 - 0x590  :   28 - 0x1c -- Sprite 0xb2
    "00110110", -- 1425 - 0x591  :   54 - 0x36
    "01100011", -- 1426 - 0x592  :   99 - 0x63
    "01100011", -- 1427 - 0x593  :   99 - 0x63
    "01111111", -- 1428 - 0x594  :  127 - 0x7f
    "01100011", -- 1429 - 0x595  :   99 - 0x63
    "01100011", -- 1430 - 0x596  :   99 - 0x63
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00110011", -- 1432 - 0x598  :   51 - 0x33 -- Sprite 0xb3
    "00110011", -- 1433 - 0x599  :   51 - 0x33
    "00110011", -- 1434 - 0x59a  :   51 - 0x33
    "00011110", -- 1435 - 0x59b  :   30 - 0x1e
    "00001100", -- 1436 - 0x59c  :   12 - 0xc
    "00001100", -- 1437 - 0x59d  :   12 - 0xc
    "00001100", -- 1438 - 0x59e  :   12 - 0xc
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01111111", -- 1440 - 0x5a0  :  127 - 0x7f -- Sprite 0xb4
    "01100000", -- 1441 - 0x5a1  :   96 - 0x60
    "01100000", -- 1442 - 0x5a2  :   96 - 0x60
    "01111110", -- 1443 - 0x5a3  :  126 - 0x7e
    "01100000", -- 1444 - 0x5a4  :   96 - 0x60
    "01100000", -- 1445 - 0x5a5  :   96 - 0x60
    "01111111", -- 1446 - 0x5a6  :  127 - 0x7f
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "01111110", -- 1448 - 0x5a8  :  126 - 0x7e -- Sprite 0xb5
    "01100011", -- 1449 - 0x5a9  :   99 - 0x63
    "01100011", -- 1450 - 0x5aa  :   99 - 0x63
    "01100111", -- 1451 - 0x5ab  :  103 - 0x67
    "01111100", -- 1452 - 0x5ac  :  124 - 0x7c
    "01101110", -- 1453 - 0x5ad  :  110 - 0x6e
    "01100111", -- 1454 - 0x5ae  :  103 - 0x67
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00111110", -- 1456 - 0x5b0  :   62 - 0x3e -- Sprite 0xb6
    "01100011", -- 1457 - 0x5b1  :   99 - 0x63
    "01100011", -- 1458 - 0x5b2  :   99 - 0x63
    "01100011", -- 1459 - 0x5b3  :   99 - 0x63
    "01100011", -- 1460 - 0x5b4  :   99 - 0x63
    "01100011", -- 1461 - 0x5b5  :   99 - 0x63
    "00111110", -- 1462 - 0x5b6  :   62 - 0x3e
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "01100011", -- 1464 - 0x5b8  :   99 - 0x63 -- Sprite 0xb7
    "01110011", -- 1465 - 0x5b9  :  115 - 0x73
    "01111011", -- 1466 - 0x5ba  :  123 - 0x7b
    "01111111", -- 1467 - 0x5bb  :  127 - 0x7f
    "01101111", -- 1468 - 0x5bc  :  111 - 0x6f
    "01100111", -- 1469 - 0x5bd  :  103 - 0x67
    "01100011", -- 1470 - 0x5be  :   99 - 0x63
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00111111", -- 1472 - 0x5c0  :   63 - 0x3f -- Sprite 0xb8
    "00001100", -- 1473 - 0x5c1  :   12 - 0xc
    "00001100", -- 1474 - 0x5c2  :   12 - 0xc
    "00001100", -- 1475 - 0x5c3  :   12 - 0xc
    "00001100", -- 1476 - 0x5c4  :   12 - 0xc
    "00001100", -- 1477 - 0x5c5  :   12 - 0xc
    "00001100", -- 1478 - 0x5c6  :   12 - 0xc
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "01100011", -- 1480 - 0x5c8  :   99 - 0x63 -- Sprite 0xb9
    "01100011", -- 1481 - 0x5c9  :   99 - 0x63
    "01101011", -- 1482 - 0x5ca  :  107 - 0x6b
    "01111111", -- 1483 - 0x5cb  :  127 - 0x7f
    "01111111", -- 1484 - 0x5cc  :  127 - 0x7f
    "01110111", -- 1485 - 0x5cd  :  119 - 0x77
    "01100011", -- 1486 - 0x5ce  :   99 - 0x63
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0 -- Sprite 0xba
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000000", -- 1490 - 0x5d2  :    0 - 0x0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00011111", -- 1504 - 0x5e0  :   31 - 0x1f -- Sprite 0xbc
    "00110000", -- 1505 - 0x5e1  :   48 - 0x30
    "01100000", -- 1506 - 0x5e2  :   96 - 0x60
    "01100111", -- 1507 - 0x5e3  :  103 - 0x67
    "01100011", -- 1508 - 0x5e4  :   99 - 0x63
    "00110011", -- 1509 - 0x5e5  :   51 - 0x33
    "00011111", -- 1510 - 0x5e6  :   31 - 0x1f
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "01100011", -- 1512 - 0x5e8  :   99 - 0x63 -- Sprite 0xbd
    "01110111", -- 1513 - 0x5e9  :  119 - 0x77
    "01111111", -- 1514 - 0x5ea  :  127 - 0x7f
    "01111111", -- 1515 - 0x5eb  :  127 - 0x7f
    "01101011", -- 1516 - 0x5ec  :  107 - 0x6b
    "01100011", -- 1517 - 0x5ed  :   99 - 0x63
    "01100011", -- 1518 - 0x5ee  :   99 - 0x63
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "01100011", -- 1520 - 0x5f0  :   99 - 0x63 -- Sprite 0xbe
    "01100011", -- 1521 - 0x5f1  :   99 - 0x63
    "01100011", -- 1522 - 0x5f2  :   99 - 0x63
    "01110111", -- 1523 - 0x5f3  :  119 - 0x77
    "00111110", -- 1524 - 0x5f4  :   62 - 0x3e
    "00011100", -- 1525 - 0x5f5  :   28 - 0x1c
    "00001000", -- 1526 - 0x5f6  :    8 - 0x8
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- Sprite 0xc5
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0 -- Sprite 0xc7
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- Sprite 0xc9
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "11111111", -- 1664 - 0x680  :  255 - 0xff -- Sprite 0xd0
    "11111111", -- 1665 - 0x681  :  255 - 0xff
    "11111111", -- 1666 - 0x682  :  255 - 0xff
    "11111111", -- 1667 - 0x683  :  255 - 0xff
    "11111111", -- 1668 - 0x684  :  255 - 0xff
    "11111111", -- 1669 - 0x685  :  255 - 0xff
    "11111111", -- 1670 - 0x686  :  255 - 0xff
    "11111111", -- 1671 - 0x687  :  255 - 0xff
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Sprite 0xd1
    "11111111", -- 1673 - 0x689  :  255 - 0xff
    "11111111", -- 1674 - 0x68a  :  255 - 0xff
    "11111111", -- 1675 - 0x68b  :  255 - 0xff
    "11111111", -- 1676 - 0x68c  :  255 - 0xff
    "11111111", -- 1677 - 0x68d  :  255 - 0xff
    "11111111", -- 1678 - 0x68e  :  255 - 0xff
    "11111111", -- 1679 - 0x68f  :  255 - 0xff
    "11111111", -- 1680 - 0x690  :  255 - 0xff -- Sprite 0xd2
    "11111111", -- 1681 - 0x691  :  255 - 0xff
    "11111111", -- 1682 - 0x692  :  255 - 0xff
    "11111111", -- 1683 - 0x693  :  255 - 0xff
    "11111111", -- 1684 - 0x694  :  255 - 0xff
    "11111111", -- 1685 - 0x695  :  255 - 0xff
    "11111111", -- 1686 - 0x696  :  255 - 0xff
    "11111111", -- 1687 - 0x697  :  255 - 0xff
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111111", -- 1692 - 0x69c  :  255 - 0xff
    "11111111", -- 1693 - 0x69d  :  255 - 0xff
    "11111111", -- 1694 - 0x69e  :  255 - 0xff
    "11111111", -- 1695 - 0x69f  :  255 - 0xff
    "11111111", -- 1696 - 0x6a0  :  255 - 0xff -- Sprite 0xd4
    "11111111", -- 1697 - 0x6a1  :  255 - 0xff
    "11111111", -- 1698 - 0x6a2  :  255 - 0xff
    "11111111", -- 1699 - 0x6a3  :  255 - 0xff
    "11111111", -- 1700 - 0x6a4  :  255 - 0xff
    "11111111", -- 1701 - 0x6a5  :  255 - 0xff
    "11111111", -- 1702 - 0x6a6  :  255 - 0xff
    "11111111", -- 1703 - 0x6a7  :  255 - 0xff
    "11111111", -- 1704 - 0x6a8  :  255 - 0xff -- Sprite 0xd5
    "11111111", -- 1705 - 0x6a9  :  255 - 0xff
    "11111111", -- 1706 - 0x6aa  :  255 - 0xff
    "11111111", -- 1707 - 0x6ab  :  255 - 0xff
    "11111111", -- 1708 - 0x6ac  :  255 - 0xff
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "11111111", -- 1712 - 0x6b0  :  255 - 0xff -- Sprite 0xd6
    "11111111", -- 1713 - 0x6b1  :  255 - 0xff
    "11111111", -- 1714 - 0x6b2  :  255 - 0xff
    "11111111", -- 1715 - 0x6b3  :  255 - 0xff
    "11111111", -- 1716 - 0x6b4  :  255 - 0xff
    "11111111", -- 1717 - 0x6b5  :  255 - 0xff
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111111", -- 1723 - 0x6bb  :  255 - 0xff
    "11111111", -- 1724 - 0x6bc  :  255 - 0xff
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11111111", -- 1732 - 0x6c4  :  255 - 0xff
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111111", -- 1734 - 0x6c6  :  255 - 0xff
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- Sprite 0xd9
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11111111", -- 1740 - 0x6cc  :  255 - 0xff
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111111", -- 1742 - 0x6ce  :  255 - 0xff
    "11111111", -- 1743 - 0x6cf  :  255 - 0xff
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Sprite 0xda
    "11111111", -- 1745 - 0x6d1  :  255 - 0xff
    "11111111", -- 1746 - 0x6d2  :  255 - 0xff
    "11111111", -- 1747 - 0x6d3  :  255 - 0xff
    "11111111", -- 1748 - 0x6d4  :  255 - 0xff
    "11111111", -- 1749 - 0x6d5  :  255 - 0xff
    "11111111", -- 1750 - 0x6d6  :  255 - 0xff
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "11111111", -- 1752 - 0x6d8  :  255 - 0xff -- Sprite 0xdb
    "11111111", -- 1753 - 0x6d9  :  255 - 0xff
    "11111111", -- 1754 - 0x6da  :  255 - 0xff
    "11111111", -- 1755 - 0x6db  :  255 - 0xff
    "11111111", -- 1756 - 0x6dc  :  255 - 0xff
    "11111111", -- 1757 - 0x6dd  :  255 - 0xff
    "11111111", -- 1758 - 0x6de  :  255 - 0xff
    "11111111", -- 1759 - 0x6df  :  255 - 0xff
    "11111111", -- 1760 - 0x6e0  :  255 - 0xff -- Sprite 0xdc
    "11111111", -- 1761 - 0x6e1  :  255 - 0xff
    "11111111", -- 1762 - 0x6e2  :  255 - 0xff
    "11111111", -- 1763 - 0x6e3  :  255 - 0xff
    "11111111", -- 1764 - 0x6e4  :  255 - 0xff
    "11111111", -- 1765 - 0x6e5  :  255 - 0xff
    "11111111", -- 1766 - 0x6e6  :  255 - 0xff
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "11111111", -- 1768 - 0x6e8  :  255 - 0xff -- Sprite 0xdd
    "11111111", -- 1769 - 0x6e9  :  255 - 0xff
    "11111111", -- 1770 - 0x6ea  :  255 - 0xff
    "11111111", -- 1771 - 0x6eb  :  255 - 0xff
    "11111111", -- 1772 - 0x6ec  :  255 - 0xff
    "11111111", -- 1773 - 0x6ed  :  255 - 0xff
    "11111111", -- 1774 - 0x6ee  :  255 - 0xff
    "11111111", -- 1775 - 0x6ef  :  255 - 0xff
    "11111111", -- 1776 - 0x6f0  :  255 - 0xff -- Sprite 0xde
    "11111111", -- 1777 - 0x6f1  :  255 - 0xff
    "11111111", -- 1778 - 0x6f2  :  255 - 0xff
    "11111111", -- 1779 - 0x6f3  :  255 - 0xff
    "11111111", -- 1780 - 0x6f4  :  255 - 0xff
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "11111111", -- 1784 - 0x6f8  :  255 - 0xff -- Sprite 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11111111", -- 1788 - 0x6fc  :  255 - 0xff
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111111", -- 1791 - 0x6ff  :  255 - 0xff
    "11111111", -- 1792 - 0x700  :  255 - 0xff -- Sprite 0xe0
    "11111111", -- 1793 - 0x701  :  255 - 0xff
    "11111111", -- 1794 - 0x702  :  255 - 0xff
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "11111111", -- 1796 - 0x704  :  255 - 0xff
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "11111111", -- 1802 - 0x70a  :  255 - 0xff
    "11111111", -- 1803 - 0x70b  :  255 - 0xff
    "11111111", -- 1804 - 0x70c  :  255 - 0xff
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Sprite 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11111111", -- 1816 - 0x718  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "11111111", -- 1818 - 0x71a  :  255 - 0xff
    "11111111", -- 1819 - 0x71b  :  255 - 0xff
    "11111111", -- 1820 - 0x71c  :  255 - 0xff
    "11111111", -- 1821 - 0x71d  :  255 - 0xff
    "11111111", -- 1822 - 0x71e  :  255 - 0xff
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "11111111", -- 1824 - 0x720  :  255 - 0xff -- Sprite 0xe4
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "11111111", -- 1826 - 0x722  :  255 - 0xff
    "11111111", -- 1827 - 0x723  :  255 - 0xff
    "11111111", -- 1828 - 0x724  :  255 - 0xff
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "11111111", -- 1834 - 0x72a  :  255 - 0xff
    "11111111", -- 1835 - 0x72b  :  255 - 0xff
    "11111111", -- 1836 - 0x72c  :  255 - 0xff
    "11111111", -- 1837 - 0x72d  :  255 - 0xff
    "11111111", -- 1838 - 0x72e  :  255 - 0xff
    "11111111", -- 1839 - 0x72f  :  255 - 0xff
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Sprite 0xe6
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11111111", -- 1843 - 0x733  :  255 - 0xff
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11111111", -- 1845 - 0x735  :  255 - 0xff
    "11111111", -- 1846 - 0x736  :  255 - 0xff
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "11111111", -- 1850 - 0x73a  :  255 - 0xff
    "11111111", -- 1851 - 0x73b  :  255 - 0xff
    "11111111", -- 1852 - 0x73c  :  255 - 0xff
    "11111111", -- 1853 - 0x73d  :  255 - 0xff
    "11111111", -- 1854 - 0x73e  :  255 - 0xff
    "11111111", -- 1855 - 0x73f  :  255 - 0xff
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11111111", -- 1864 - 0x748  :  255 - 0xff -- Sprite 0xe9
    "11111111", -- 1865 - 0x749  :  255 - 0xff
    "11111111", -- 1866 - 0x74a  :  255 - 0xff
    "11111111", -- 1867 - 0x74b  :  255 - 0xff
    "11111111", -- 1868 - 0x74c  :  255 - 0xff
    "11111111", -- 1869 - 0x74d  :  255 - 0xff
    "11111111", -- 1870 - 0x74e  :  255 - 0xff
    "11111111", -- 1871 - 0x74f  :  255 - 0xff
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "11111111", -- 1880 - 0x758  :  255 - 0xff -- Sprite 0xeb
    "11111111", -- 1881 - 0x759  :  255 - 0xff
    "11111111", -- 1882 - 0x75a  :  255 - 0xff
    "11111111", -- 1883 - 0x75b  :  255 - 0xff
    "11111111", -- 1884 - 0x75c  :  255 - 0xff
    "11111111", -- 1885 - 0x75d  :  255 - 0xff
    "11111111", -- 1886 - 0x75e  :  255 - 0xff
    "11111111", -- 1887 - 0x75f  :  255 - 0xff
    "11111111", -- 1888 - 0x760  :  255 - 0xff -- Sprite 0xec
    "11111111", -- 1889 - 0x761  :  255 - 0xff
    "11111111", -- 1890 - 0x762  :  255 - 0xff
    "11111111", -- 1891 - 0x763  :  255 - 0xff
    "11111111", -- 1892 - 0x764  :  255 - 0xff
    "11111111", -- 1893 - 0x765  :  255 - 0xff
    "11111111", -- 1894 - 0x766  :  255 - 0xff
    "11111111", -- 1895 - 0x767  :  255 - 0xff
    "11111111", -- 1896 - 0x768  :  255 - 0xff -- Sprite 0xed
    "11111111", -- 1897 - 0x769  :  255 - 0xff
    "11111111", -- 1898 - 0x76a  :  255 - 0xff
    "11111111", -- 1899 - 0x76b  :  255 - 0xff
    "11111111", -- 1900 - 0x76c  :  255 - 0xff
    "11111111", -- 1901 - 0x76d  :  255 - 0xff
    "11111111", -- 1902 - 0x76e  :  255 - 0xff
    "11111111", -- 1903 - 0x76f  :  255 - 0xff
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Sprite 0xee
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "11111111", -- 1906 - 0x772  :  255 - 0xff
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111111", -- 1909 - 0x775  :  255 - 0xff
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "11111111", -- 1912 - 0x778  :  255 - 0xff -- Sprite 0xef
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111111", -- 1914 - 0x77a  :  255 - 0xff
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111111", -- 1916 - 0x77c  :  255 - 0xff
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11111111", -- 1919 - 0x77f  :  255 - 0xff
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- Sprite 0xf3
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Sprite 0xf4
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- Sprite 0xf5
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Sprite 0xf6
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff -- Sprite 0xf7
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Sprite 0xfc
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff -- Sprite 0xfd
    "11111111", -- 2025 - 0x7e9  :  255 - 0xff
    "11111111", -- 2026 - 0x7ea  :  255 - 0xff
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111111", -- 2028 - 0x7ec  :  255 - 0xff
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Sprite 0xfe
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111", -- 2047 - 0x7ff  :  255 - 0xff
          -- Background pattern Table
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Background 0x0
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000000", -- 2050 - 0x802  :    0 - 0x0
    "00000000", -- 2051 - 0x803  :    0 - 0x0
    "00000000", -- 2052 - 0x804  :    0 - 0x0
    "00000000", -- 2053 - 0x805  :    0 - 0x0
    "00000000", -- 2054 - 0x806  :    0 - 0x0
    "00000000", -- 2055 - 0x807  :    0 - 0x0
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- Background 0x1
    "00111000", -- 2057 - 0x809  :   56 - 0x38
    "01111100", -- 2058 - 0x80a  :  124 - 0x7c
    "11111110", -- 2059 - 0x80b  :  254 - 0xfe
    "11111110", -- 2060 - 0x80c  :  254 - 0xfe
    "11111110", -- 2061 - 0x80d  :  254 - 0xfe
    "01111100", -- 2062 - 0x80e  :  124 - 0x7c
    "00111000", -- 2063 - 0x80f  :   56 - 0x38
    "00000000", -- 2064 - 0x810  :    0 - 0x0 -- Background 0x2
    "00000000", -- 2065 - 0x811  :    0 - 0x0
    "00000000", -- 2066 - 0x812  :    0 - 0x0
    "00000000", -- 2067 - 0x813  :    0 - 0x0
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- Background 0x3
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00011000", -- 2075 - 0x81b  :   24 - 0x18
    "00011000", -- 2076 - 0x81c  :   24 - 0x18
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Background 0x4
    "11111111", -- 2081 - 0x821  :  255 - 0xff
    "11111111", -- 2082 - 0x822  :  255 - 0xff
    "11111111", -- 2083 - 0x823  :  255 - 0xff
    "11111111", -- 2084 - 0x824  :  255 - 0xff
    "11111111", -- 2085 - 0x825  :  255 - 0xff
    "11111111", -- 2086 - 0x826  :  255 - 0xff
    "11111111", -- 2087 - 0x827  :  255 - 0xff
    "00001111", -- 2088 - 0x828  :   15 - 0xf -- Background 0x5
    "00001111", -- 2089 - 0x829  :   15 - 0xf
    "00001111", -- 2090 - 0x82a  :   15 - 0xf
    "00001111", -- 2091 - 0x82b  :   15 - 0xf
    "00001111", -- 2092 - 0x82c  :   15 - 0xf
    "00001111", -- 2093 - 0x82d  :   15 - 0xf
    "00001111", -- 2094 - 0x82e  :   15 - 0xf
    "00001111", -- 2095 - 0x82f  :   15 - 0xf
    "11110000", -- 2096 - 0x830  :  240 - 0xf0 -- Background 0x6
    "11110000", -- 2097 - 0x831  :  240 - 0xf0
    "11110000", -- 2098 - 0x832  :  240 - 0xf0
    "11110000", -- 2099 - 0x833  :  240 - 0xf0
    "11110000", -- 2100 - 0x834  :  240 - 0xf0
    "11110000", -- 2101 - 0x835  :  240 - 0xf0
    "11110000", -- 2102 - 0x836  :  240 - 0xf0
    "11110000", -- 2103 - 0x837  :  240 - 0xf0
    "00000000", -- 2104 - 0x838  :    0 - 0x0 -- Background 0x7
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00000000", -- 2108 - 0x83c  :    0 - 0x0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0 -- Background 0x8
    "00000000", -- 2113 - 0x841  :    0 - 0x0
    "00000000", -- 2114 - 0x842  :    0 - 0x0
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000000", -- 2116 - 0x844  :    0 - 0x0
    "00000000", -- 2117 - 0x845  :    0 - 0x0
    "00000000", -- 2118 - 0x846  :    0 - 0x0
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- Background 0x9
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00011000", -- 2123 - 0x84b  :   24 - 0x18
    "00011000", -- 2124 - 0x84c  :   24 - 0x18
    "00000000", -- 2125 - 0x84d  :    0 - 0x0
    "00000000", -- 2126 - 0x84e  :    0 - 0x0
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "00000000", -- 2128 - 0x850  :    0 - 0x0 -- Background 0xa
    "00000000", -- 2129 - 0x851  :    0 - 0x0
    "00000000", -- 2130 - 0x852  :    0 - 0x0
    "00000000", -- 2131 - 0x853  :    0 - 0x0
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00000000", -- 2136 - 0x858  :    0 - 0x0 -- Background 0xb
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Background 0xc
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "00000000", -- 2148 - 0x864  :    0 - 0x0
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00000000", -- 2150 - 0x866  :    0 - 0x0
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- Background 0xd
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "00000000", -- 2157 - 0x86d  :    0 - 0x0
    "00000000", -- 2158 - 0x86e  :    0 - 0x0
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0 -- Background 0xe
    "00000000", -- 2161 - 0x871  :    0 - 0x0
    "00000000", -- 2162 - 0x872  :    0 - 0x0
    "00000000", -- 2163 - 0x873  :    0 - 0x0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- Background 0xf
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Background 0x10
    "00000000", -- 2177 - 0x881  :    0 - 0x0
    "00000000", -- 2178 - 0x882  :    0 - 0x0
    "00000000", -- 2179 - 0x883  :    0 - 0x0
    "00000000", -- 2180 - 0x884  :    0 - 0x0
    "00000000", -- 2181 - 0x885  :    0 - 0x0
    "00000000", -- 2182 - 0x886  :    0 - 0x0
    "00000000", -- 2183 - 0x887  :    0 - 0x0
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- Background 0x11
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000000", -- 2187 - 0x88b  :    0 - 0x0
    "00000000", -- 2188 - 0x88c  :    0 - 0x0
    "00000000", -- 2189 - 0x88d  :    0 - 0x0
    "00000000", -- 2190 - 0x88e  :    0 - 0x0
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "00000000", -- 2192 - 0x890  :    0 - 0x0 -- Background 0x12
    "00000000", -- 2193 - 0x891  :    0 - 0x0
    "00000000", -- 2194 - 0x892  :    0 - 0x0
    "00000000", -- 2195 - 0x893  :    0 - 0x0
    "00000000", -- 2196 - 0x894  :    0 - 0x0
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000000", -- 2200 - 0x898  :    0 - 0x0 -- Background 0x13
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000000", -- 2202 - 0x89a  :    0 - 0x0
    "00000000", -- 2203 - 0x89b  :    0 - 0x0
    "00000000", -- 2204 - 0x89c  :    0 - 0x0
    "00000000", -- 2205 - 0x89d  :    0 - 0x0
    "00000000", -- 2206 - 0x89e  :    0 - 0x0
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x14
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "00000000", -- 2212 - 0x8a4  :    0 - 0x0
    "00000000", -- 2213 - 0x8a5  :    0 - 0x0
    "00000000", -- 2214 - 0x8a6  :    0 - 0x0
    "00000000", -- 2215 - 0x8a7  :    0 - 0x0
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- Background 0x15
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00000000", -- 2222 - 0x8ae  :    0 - 0x0
    "00000000", -- 2223 - 0x8af  :    0 - 0x0
    "00000000", -- 2224 - 0x8b0  :    0 - 0x0 -- Background 0x16
    "00000000", -- 2225 - 0x8b1  :    0 - 0x0
    "00000000", -- 2226 - 0x8b2  :    0 - 0x0
    "00000000", -- 2227 - 0x8b3  :    0 - 0x0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "00000000", -- 2230 - 0x8b6  :    0 - 0x0
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00000000", -- 2232 - 0x8b8  :    0 - 0x0 -- Background 0x17
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00000000", -- 2234 - 0x8ba  :    0 - 0x0
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00000000", -- 2236 - 0x8bc  :    0 - 0x0
    "00000000", -- 2237 - 0x8bd  :    0 - 0x0
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Background 0x18
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000000", -- 2244 - 0x8c4  :    0 - 0x0
    "00000000", -- 2245 - 0x8c5  :    0 - 0x0
    "00000000", -- 2246 - 0x8c6  :    0 - 0x0
    "00000000", -- 2247 - 0x8c7  :    0 - 0x0
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- Background 0x19
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000000", -- 2251 - 0x8cb  :    0 - 0x0
    "00000000", -- 2252 - 0x8cc  :    0 - 0x0
    "00000000", -- 2253 - 0x8cd  :    0 - 0x0
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "00000000", -- 2256 - 0x8d0  :    0 - 0x0 -- Background 0x1a
    "00000000", -- 2257 - 0x8d1  :    0 - 0x0
    "00000000", -- 2258 - 0x8d2  :    0 - 0x0
    "00000000", -- 2259 - 0x8d3  :    0 - 0x0
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- Background 0x1b
    "00000000", -- 2265 - 0x8d9  :    0 - 0x0
    "00000000", -- 2266 - 0x8da  :    0 - 0x0
    "00000000", -- 2267 - 0x8db  :    0 - 0x0
    "00000000", -- 2268 - 0x8dc  :    0 - 0x0
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000000", -- 2270 - 0x8de  :    0 - 0x0
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Background 0x1c
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "00000000", -- 2276 - 0x8e4  :    0 - 0x0
    "00000000", -- 2277 - 0x8e5  :    0 - 0x0
    "00000000", -- 2278 - 0x8e6  :    0 - 0x0
    "00000000", -- 2279 - 0x8e7  :    0 - 0x0
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- Background 0x1d
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "00000000", -- 2283 - 0x8eb  :    0 - 0x0
    "00000000", -- 2284 - 0x8ec  :    0 - 0x0
    "00000000", -- 2285 - 0x8ed  :    0 - 0x0
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "00000000", -- 2288 - 0x8f0  :    0 - 0x0 -- Background 0x1e
    "00000000", -- 2289 - 0x8f1  :    0 - 0x0
    "00000000", -- 2290 - 0x8f2  :    0 - 0x0
    "00000000", -- 2291 - 0x8f3  :    0 - 0x0
    "00000000", -- 2292 - 0x8f4  :    0 - 0x0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0 -- Background 0x1f
    "00000000", -- 2297 - 0x8f9  :    0 - 0x0
    "00000000", -- 2298 - 0x8fa  :    0 - 0x0
    "00000000", -- 2299 - 0x8fb  :    0 - 0x0
    "00000000", -- 2300 - 0x8fc  :    0 - 0x0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x20
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00000000", -- 2307 - 0x903  :    0 - 0x0
    "00000000", -- 2308 - 0x904  :    0 - 0x0
    "00000000", -- 2309 - 0x905  :    0 - 0x0
    "00000000", -- 2310 - 0x906  :    0 - 0x0
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "00001111", -- 2312 - 0x908  :   15 - 0xf -- Background 0x21
    "00001111", -- 2313 - 0x909  :   15 - 0xf
    "00001111", -- 2314 - 0x90a  :   15 - 0xf
    "00000111", -- 2315 - 0x90b  :    7 - 0x7
    "00000111", -- 2316 - 0x90c  :    7 - 0x7
    "00001111", -- 2317 - 0x90d  :   15 - 0xf
    "00001111", -- 2318 - 0x90e  :   15 - 0xf
    "00001111", -- 2319 - 0x90f  :   15 - 0xf
    "11110000", -- 2320 - 0x910  :  240 - 0xf0 -- Background 0x22
    "11110000", -- 2321 - 0x911  :  240 - 0xf0
    "11110000", -- 2322 - 0x912  :  240 - 0xf0
    "11100000", -- 2323 - 0x913  :  224 - 0xe0
    "11100000", -- 2324 - 0x914  :  224 - 0xe0
    "11110000", -- 2325 - 0x915  :  240 - 0xf0
    "11110000", -- 2326 - 0x916  :  240 - 0xf0
    "11110000", -- 2327 - 0x917  :  240 - 0xf0
    "11111111", -- 2328 - 0x918  :  255 - 0xff -- Background 0x23
    "11111111", -- 2329 - 0x919  :  255 - 0xff
    "11100001", -- 2330 - 0x91a  :  225 - 0xe1
    "11100001", -- 2331 - 0x91b  :  225 - 0xe1
    "11100001", -- 2332 - 0x91c  :  225 - 0xe1
    "11100001", -- 2333 - 0x91d  :  225 - 0xe1
    "11100001", -- 2334 - 0x91e  :  225 - 0xe1
    "11100001", -- 2335 - 0x91f  :  225 - 0xe1
    "10000111", -- 2336 - 0x920  :  135 - 0x87 -- Background 0x24
    "11000111", -- 2337 - 0x921  :  199 - 0xc7
    "11000000", -- 2338 - 0x922  :  192 - 0xc0
    "11000111", -- 2339 - 0x923  :  199 - 0xc7
    "11001111", -- 2340 - 0x924  :  207 - 0xcf
    "11001110", -- 2341 - 0x925  :  206 - 0xce
    "11001111", -- 2342 - 0x926  :  207 - 0xcf
    "11000111", -- 2343 - 0x927  :  199 - 0xc7
    "11111000", -- 2344 - 0x928  :  248 - 0xf8 -- Background 0x25
    "11111100", -- 2345 - 0x929  :  252 - 0xfc
    "00011100", -- 2346 - 0x92a  :   28 - 0x1c
    "11111100", -- 2347 - 0x92b  :  252 - 0xfc
    "11111100", -- 2348 - 0x92c  :  252 - 0xfc
    "00011100", -- 2349 - 0x92d  :   28 - 0x1c
    "11111100", -- 2350 - 0x92e  :  252 - 0xfc
    "11111100", -- 2351 - 0x92f  :  252 - 0xfc
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Background 0x26
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "11100111", -- 2354 - 0x932  :  231 - 0xe7
    "11100111", -- 2355 - 0x933  :  231 - 0xe7
    "11100111", -- 2356 - 0x934  :  231 - 0xe7
    "11100111", -- 2357 - 0x935  :  231 - 0xe7
    "11100111", -- 2358 - 0x936  :  231 - 0xe7
    "11100111", -- 2359 - 0x937  :  231 - 0xe7
    "11110000", -- 2360 - 0x938  :  240 - 0xf0 -- Background 0x27
    "11111001", -- 2361 - 0x939  :  249 - 0xf9
    "00111001", -- 2362 - 0x93a  :   57 - 0x39
    "00111001", -- 2363 - 0x93b  :   57 - 0x39
    "00111001", -- 2364 - 0x93c  :   57 - 0x39
    "00111001", -- 2365 - 0x93d  :   57 - 0x39
    "00111001", -- 2366 - 0x93e  :   57 - 0x39
    "00111000", -- 2367 - 0x93f  :   56 - 0x38
    "11111111", -- 2368 - 0x940  :  255 - 0xff -- Background 0x28
    "11111111", -- 2369 - 0x941  :  255 - 0xff
    "11000000", -- 2370 - 0x942  :  192 - 0xc0
    "11000000", -- 2371 - 0x943  :  192 - 0xc0
    "11000000", -- 2372 - 0x944  :  192 - 0xc0
    "11000000", -- 2373 - 0x945  :  192 - 0xc0
    "11111111", -- 2374 - 0x946  :  255 - 0xff
    "11111111", -- 2375 - 0x947  :  255 - 0xff
    "00011111", -- 2376 - 0x948  :   31 - 0x1f -- Background 0x29
    "00111111", -- 2377 - 0x949  :   63 - 0x3f
    "00110000", -- 2378 - 0x94a  :   48 - 0x30
    "00110000", -- 2379 - 0x94b  :   48 - 0x30
    "00110000", -- 2380 - 0x94c  :   48 - 0x30
    "00110000", -- 2381 - 0x94d  :   48 - 0x30
    "00111111", -- 2382 - 0x94e  :   63 - 0x3f
    "00011111", -- 2383 - 0x94f  :   31 - 0x1f
    "11100011", -- 2384 - 0x950  :  227 - 0xe3 -- Background 0x2a
    "11110011", -- 2385 - 0x951  :  243 - 0xf3
    "01110000", -- 2386 - 0x952  :  112 - 0x70
    "01110000", -- 2387 - 0x953  :  112 - 0x70
    "01110000", -- 2388 - 0x954  :  112 - 0x70
    "01110000", -- 2389 - 0x955  :  112 - 0x70
    "11110000", -- 2390 - 0x956  :  240 - 0xf0
    "11100000", -- 2391 - 0x957  :  224 - 0xe0
    "11111110", -- 2392 - 0x958  :  254 - 0xfe -- Background 0x2b
    "11111110", -- 2393 - 0x959  :  254 - 0xfe
    "01110000", -- 2394 - 0x95a  :  112 - 0x70
    "01110000", -- 2395 - 0x95b  :  112 - 0x70
    "01110000", -- 2396 - 0x95c  :  112 - 0x70
    "01110000", -- 2397 - 0x95d  :  112 - 0x70
    "01110000", -- 2398 - 0x95e  :  112 - 0x70
    "01110000", -- 2399 - 0x95f  :  112 - 0x70
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "11111111", -- 2408 - 0x968  :  255 - 0xff -- Background 0x2d
    "11111111", -- 2409 - 0x969  :  255 - 0xff
    "11111111", -- 2410 - 0x96a  :  255 - 0xff
    "11111111", -- 2411 - 0x96b  :  255 - 0xff
    "11111111", -- 2412 - 0x96c  :  255 - 0xff
    "11111111", -- 2413 - 0x96d  :  255 - 0xff
    "11111111", -- 2414 - 0x96e  :  255 - 0xff
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000000", -- 2424 - 0x978  :    0 - 0x0 -- Background 0x2f
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "00000000", -- 2426 - 0x97a  :    0 - 0x0
    "00011000", -- 2427 - 0x97b  :   24 - 0x18
    "00011000", -- 2428 - 0x97c  :   24 - 0x18
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Background 0x30
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "00000000", -- 2436 - 0x984  :    0 - 0x0
    "00000000", -- 2437 - 0x985  :    0 - 0x0
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- Background 0x31
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Background 0x32
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "00000000", -- 2453 - 0x995  :    0 - 0x0
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "00000000", -- 2456 - 0x998  :    0 - 0x0 -- Background 0x33
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Background 0x34
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00000000", -- 2466 - 0x9a2  :    0 - 0x0
    "00000000", -- 2467 - 0x9a3  :    0 - 0x0
    "00000000", -- 2468 - 0x9a4  :    0 - 0x0
    "00000000", -- 2469 - 0x9a5  :    0 - 0x0
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- Background 0x35
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0 -- Background 0x36
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "00000000", -- 2485 - 0x9b5  :    0 - 0x0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0 -- Background 0x37
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000111", -- 2529 - 0x9e1  :    7 - 0x7
    "00011111", -- 2530 - 0x9e2  :   31 - 0x1f
    "00111111", -- 2531 - 0x9e3  :   63 - 0x3f
    "00111111", -- 2532 - 0x9e4  :   63 - 0x3f
    "00001111", -- 2533 - 0x9e5  :   15 - 0xf
    "00000011", -- 2534 - 0x9e6  :    3 - 0x3
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "11000000", -- 2537 - 0x9e9  :  192 - 0xc0
    "11110000", -- 2538 - 0x9ea  :  240 - 0xf0
    "11111000", -- 2539 - 0x9eb  :  248 - 0xf8
    "11111000", -- 2540 - 0x9ec  :  248 - 0xf8
    "11111100", -- 2541 - 0x9ed  :  252 - 0xfc
    "11111100", -- 2542 - 0x9ee  :  252 - 0xfc
    "11111100", -- 2543 - 0x9ef  :  252 - 0xfc
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "00000011", -- 2545 - 0x9f1  :    3 - 0x3
    "00001111", -- 2546 - 0x9f2  :   15 - 0xf
    "00111111", -- 2547 - 0x9f3  :   63 - 0x3f
    "00111111", -- 2548 - 0x9f4  :   63 - 0x3f
    "00011111", -- 2549 - 0x9f5  :   31 - 0x1f
    "00000111", -- 2550 - 0x9f6  :    7 - 0x7
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "11111100", -- 2552 - 0x9f8  :  252 - 0xfc -- Background 0x3f
    "11111100", -- 2553 - 0x9f9  :  252 - 0xfc
    "11111100", -- 2554 - 0x9fa  :  252 - 0xfc
    "11111000", -- 2555 - 0x9fb  :  248 - 0xf8
    "11111000", -- 2556 - 0x9fc  :  248 - 0xf8
    "11110000", -- 2557 - 0x9fd  :  240 - 0xf0
    "11000000", -- 2558 - 0x9fe  :  192 - 0xc0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Background 0x40
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- Background 0x41
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Background 0x42
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "00000000", -- 2580 - 0xa14  :    0 - 0x0
    "00000000", -- 2581 - 0xa15  :    0 - 0x0
    "00000000", -- 2582 - 0xa16  :    0 - 0x0
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00000000", -- 2584 - 0xa18  :    0 - 0x0 -- Background 0x43
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Background 0x44
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "00000000", -- 2594 - 0xa22  :    0 - 0x0
    "00000000", -- 2595 - 0xa23  :    0 - 0x0
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "00000000", -- 2598 - 0xa26  :    0 - 0x0
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- Background 0x45
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00000000", -- 2608 - 0xa30  :    0 - 0x0 -- Background 0x46
    "00000000", -- 2609 - 0xa31  :    0 - 0x0
    "00000000", -- 2610 - 0xa32  :    0 - 0x0
    "00000000", -- 2611 - 0xa33  :    0 - 0x0
    "00000000", -- 2612 - 0xa34  :    0 - 0x0
    "00000000", -- 2613 - 0xa35  :    0 - 0x0
    "00000000", -- 2614 - 0xa36  :    0 - 0x0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- Background 0x47
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0x48
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- Background 0x49
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "00000000", -- 2648 - 0xa58  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00000000", -- 2658 - 0xa62  :    0 - 0x0
    "00000000", -- 2659 - 0xa63  :    0 - 0x0
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00000000", -- 2669 - 0xa6d  :    0 - 0x0
    "00000000", -- 2670 - 0xa6e  :    0 - 0x0
    "00000000", -- 2671 - 0xa6f  :    0 - 0x0
    "00000000", -- 2672 - 0xa70  :    0 - 0x0 -- Background 0x4e
    "00000000", -- 2673 - 0xa71  :    0 - 0x0
    "00000000", -- 2674 - 0xa72  :    0 - 0x0
    "00000000", -- 2675 - 0xa73  :    0 - 0x0
    "00000000", -- 2676 - 0xa74  :    0 - 0x0
    "00000000", -- 2677 - 0xa75  :    0 - 0x0
    "00000000", -- 2678 - 0xa76  :    0 - 0x0
    "00000000", -- 2679 - 0xa77  :    0 - 0x0
    "00000000", -- 2680 - 0xa78  :    0 - 0x0 -- Background 0x4f
    "00000000", -- 2681 - 0xa79  :    0 - 0x0
    "00000000", -- 2682 - 0xa7a  :    0 - 0x0
    "00000000", -- 2683 - 0xa7b  :    0 - 0x0
    "00000000", -- 2684 - 0xa7c  :    0 - 0x0
    "00000000", -- 2685 - 0xa7d  :    0 - 0x0
    "00000000", -- 2686 - 0xa7e  :    0 - 0x0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Background 0x50
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00000000", -- 2693 - 0xa85  :    0 - 0x0
    "00000000", -- 2694 - 0xa86  :    0 - 0x0
    "00000000", -- 2695 - 0xa87  :    0 - 0x0
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- Background 0x51
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000000", -- 2702 - 0xa8e  :    0 - 0x0
    "00000000", -- 2703 - 0xa8f  :    0 - 0x0
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00000000", -- 2706 - 0xa92  :    0 - 0x0
    "00000000", -- 2707 - 0xa93  :    0 - 0x0
    "00000000", -- 2708 - 0xa94  :    0 - 0x0
    "00000000", -- 2709 - 0xa95  :    0 - 0x0
    "00000000", -- 2710 - 0xa96  :    0 - 0x0
    "00000000", -- 2711 - 0xa97  :    0 - 0x0
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- Background 0x53
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Background 0x54
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "00000000", -- 2724 - 0xaa4  :    0 - 0x0
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- Background 0x55
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "00000000", -- 2733 - 0xaad  :    0 - 0x0
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "00000000", -- 2736 - 0xab0  :    0 - 0x0 -- Background 0x56
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- Background 0x57
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Background 0x58
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- Background 0x59
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 2769 - 0xad1  :    0 - 0x0
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "00000000", -- 2771 - 0xad3  :    0 - 0x0
    "00000000", -- 2772 - 0xad4  :    0 - 0x0
    "00000000", -- 2773 - 0xad5  :    0 - 0x0
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000000", -- 2786 - 0xae2  :    0 - 0x0
    "00000000", -- 2787 - 0xae3  :    0 - 0x0
    "00000000", -- 2788 - 0xae4  :    0 - 0x0
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "00000000", -- 2800 - 0xaf0  :    0 - 0x0 -- Background 0x5e
    "00000000", -- 2801 - 0xaf1  :    0 - 0x0
    "00010000", -- 2802 - 0xaf2  :   16 - 0x10
    "00010000", -- 2803 - 0xaf3  :   16 - 0x10
    "00010000", -- 2804 - 0xaf4  :   16 - 0x10
    "00010000", -- 2805 - 0xaf5  :   16 - 0x10
    "00000000", -- 2806 - 0xaf6  :    0 - 0x0
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Background 0x60
    "00000000", -- 2817 - 0xb01  :    0 - 0x0
    "00000000", -- 2818 - 0xb02  :    0 - 0x0
    "00000000", -- 2819 - 0xb03  :    0 - 0x0
    "00000000", -- 2820 - 0xb04  :    0 - 0x0
    "00000000", -- 2821 - 0xb05  :    0 - 0x0
    "00000000", -- 2822 - 0xb06  :    0 - 0x0
    "00000000", -- 2823 - 0xb07  :    0 - 0x0
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- Background 0x61
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "00000000", -- 2826 - 0xb0a  :    0 - 0x0
    "00000000", -- 2827 - 0xb0b  :    0 - 0x0
    "00000000", -- 2828 - 0xb0c  :    0 - 0x0
    "00000000", -- 2829 - 0xb0d  :    0 - 0x0
    "00000000", -- 2830 - 0xb0e  :    0 - 0x0
    "00000000", -- 2831 - 0xb0f  :    0 - 0x0
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Background 0x62
    "00000000", -- 2833 - 0xb11  :    0 - 0x0
    "00000000", -- 2834 - 0xb12  :    0 - 0x0
    "00000000", -- 2835 - 0xb13  :    0 - 0x0
    "00000000", -- 2836 - 0xb14  :    0 - 0x0
    "00000000", -- 2837 - 0xb15  :    0 - 0x0
    "00000000", -- 2838 - 0xb16  :    0 - 0x0
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "00000000", -- 2840 - 0xb18  :    0 - 0x0 -- Background 0x63
    "00000000", -- 2841 - 0xb19  :    0 - 0x0
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "00000000", -- 2845 - 0xb1d  :    0 - 0x0
    "00000000", -- 2846 - 0xb1e  :    0 - 0x0
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0x64
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000000", -- 2851 - 0xb23  :    0 - 0x0
    "00000000", -- 2852 - 0xb24  :    0 - 0x0
    "00000000", -- 2853 - 0xb25  :    0 - 0x0
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00000000", -- 2856 - 0xb28  :    0 - 0x0 -- Background 0x65
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000000", -- 2858 - 0xb2a  :    0 - 0x0
    "00000000", -- 2859 - 0xb2b  :    0 - 0x0
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00000000", -- 2861 - 0xb2d  :    0 - 0x0
    "00000000", -- 2862 - 0xb2e  :    0 - 0x0
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00000000", -- 2864 - 0xb30  :    0 - 0x0 -- Background 0x66
    "00000000", -- 2865 - 0xb31  :    0 - 0x0
    "00000000", -- 2866 - 0xb32  :    0 - 0x0
    "00000000", -- 2867 - 0xb33  :    0 - 0x0
    "00000000", -- 2868 - 0xb34  :    0 - 0x0
    "00000000", -- 2869 - 0xb35  :    0 - 0x0
    "00000000", -- 2870 - 0xb36  :    0 - 0x0
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "00000000", -- 2872 - 0xb38  :    0 - 0x0 -- Background 0x67
    "00000000", -- 2873 - 0xb39  :    0 - 0x0
    "00000000", -- 2874 - 0xb3a  :    0 - 0x0
    "00000000", -- 2875 - 0xb3b  :    0 - 0x0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Background 0x68
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000001", -- 2883 - 0xb43  :    1 - 0x1
    "00000001", -- 2884 - 0xb44  :    1 - 0x1
    "00001011", -- 2885 - 0xb45  :   11 - 0xb
    "00011100", -- 2886 - 0xb46  :   28 - 0x1c
    "00111111", -- 2887 - 0xb47  :   63 - 0x3f
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- Background 0x69
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00110000", -- 2890 - 0xb4a  :   48 - 0x30
    "01111000", -- 2891 - 0xb4b  :  120 - 0x78
    "10000000", -- 2892 - 0xb4c  :  128 - 0x80
    "11110000", -- 2893 - 0xb4d  :  240 - 0xf0
    "11111000", -- 2894 - 0xb4e  :  248 - 0xf8
    "11111100", -- 2895 - 0xb4f  :  252 - 0xfc
    "00111111", -- 2896 - 0xb50  :   63 - 0x3f -- Background 0x6a
    "00111111", -- 2897 - 0xb51  :   63 - 0x3f
    "00111111", -- 2898 - 0xb52  :   63 - 0x3f
    "00011111", -- 2899 - 0xb53  :   31 - 0x1f
    "00011111", -- 2900 - 0xb54  :   31 - 0x1f
    "00000111", -- 2901 - 0xb55  :    7 - 0x7
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "11111100", -- 2904 - 0xb58  :  252 - 0xfc -- Background 0x6b
    "11101100", -- 2905 - 0xb59  :  236 - 0xec
    "11101100", -- 2906 - 0xb5a  :  236 - 0xec
    "11011000", -- 2907 - 0xb5b  :  216 - 0xd8
    "11111000", -- 2908 - 0xb5c  :  248 - 0xf8
    "11100000", -- 2909 - 0xb5d  :  224 - 0xe0
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000001", -- 2914 - 0xb62  :    1 - 0x1
    "00011101", -- 2915 - 0xb63  :   29 - 0x1d
    "00111110", -- 2916 - 0xb64  :   62 - 0x3e
    "00111111", -- 2917 - 0xb65  :   63 - 0x3f
    "00111111", -- 2918 - 0xb66  :   63 - 0x3f
    "00111111", -- 2919 - 0xb67  :   63 - 0x3f
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "10000000", -- 2921 - 0xb69  :  128 - 0x80
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "01110000", -- 2923 - 0xb6b  :  112 - 0x70
    "11111000", -- 2924 - 0xb6c  :  248 - 0xf8
    "11111100", -- 2925 - 0xb6d  :  252 - 0xfc
    "11111100", -- 2926 - 0xb6e  :  252 - 0xfc
    "11111100", -- 2927 - 0xb6f  :  252 - 0xfc
    "00111111", -- 2928 - 0xb70  :   63 - 0x3f -- Background 0x6e
    "00111111", -- 2929 - 0xb71  :   63 - 0x3f
    "00011111", -- 2930 - 0xb72  :   31 - 0x1f
    "00011111", -- 2931 - 0xb73  :   31 - 0x1f
    "00001111", -- 2932 - 0xb74  :   15 - 0xf
    "00000110", -- 2933 - 0xb75  :    6 - 0x6
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "11101100", -- 2936 - 0xb78  :  236 - 0xec -- Background 0x6f
    "11101100", -- 2937 - 0xb79  :  236 - 0xec
    "11011000", -- 2938 - 0xb7a  :  216 - 0xd8
    "11111000", -- 2939 - 0xb7b  :  248 - 0xf8
    "11110000", -- 2940 - 0xb7c  :  240 - 0xf0
    "11100000", -- 2941 - 0xb7d  :  224 - 0xe0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0x70
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000000", -- 2946 - 0xb82  :    0 - 0x0
    "00000000", -- 2947 - 0xb83  :    0 - 0x0
    "00000000", -- 2948 - 0xb84  :    0 - 0x0
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- Background 0x71
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "00000000", -- 2957 - 0xb8d  :    0 - 0x0
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Background 0x72
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "00000000", -- 2962 - 0xb92  :    0 - 0x0
    "00000000", -- 2963 - 0xb93  :    0 - 0x0
    "00000000", -- 2964 - 0xb94  :    0 - 0x0
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- Background 0x73
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Background 0x74
    "00000000", -- 2977 - 0xba1  :    0 - 0x0
    "00000000", -- 2978 - 0xba2  :    0 - 0x0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00010001", -- 2980 - 0xba4  :   17 - 0x11
    "00010011", -- 2981 - 0xba5  :   19 - 0x13
    "00011111", -- 2982 - 0xba6  :   31 - 0x1f
    "00011111", -- 2983 - 0xba7  :   31 - 0x1f
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- Background 0x75
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "10000000", -- 2987 - 0xbab  :  128 - 0x80
    "11000100", -- 2988 - 0xbac  :  196 - 0xc4
    "11100100", -- 2989 - 0xbad  :  228 - 0xe4
    "11111100", -- 2990 - 0xbae  :  252 - 0xfc
    "11111100", -- 2991 - 0xbaf  :  252 - 0xfc
    "00011111", -- 2992 - 0xbb0  :   31 - 0x1f -- Background 0x76
    "00001110", -- 2993 - 0xbb1  :   14 - 0xe
    "00000110", -- 2994 - 0xbb2  :    6 - 0x6
    "00000010", -- 2995 - 0xbb3  :    2 - 0x2
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "11111100", -- 3000 - 0xbb8  :  252 - 0xfc -- Background 0x77
    "10111000", -- 3001 - 0xbb9  :  184 - 0xb8
    "10110000", -- 3002 - 0xbba  :  176 - 0xb0
    "10100000", -- 3003 - 0xbbb  :  160 - 0xa0
    "10000000", -- 3004 - 0xbbc  :  128 - 0x80
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000001", -- 3011 - 0xbc3  :    1 - 0x1
    "00000011", -- 3012 - 0xbc4  :    3 - 0x3
    "00000110", -- 3013 - 0xbc5  :    6 - 0x6
    "00000110", -- 3014 - 0xbc6  :    6 - 0x6
    "00001111", -- 3015 - 0xbc7  :   15 - 0xf
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- Background 0x79
    "00011000", -- 3017 - 0xbc9  :   24 - 0x18
    "11110100", -- 3018 - 0xbca  :  244 - 0xf4
    "11111000", -- 3019 - 0xbcb  :  248 - 0xf8
    "00111000", -- 3020 - 0xbcc  :   56 - 0x38
    "01111100", -- 3021 - 0xbcd  :  124 - 0x7c
    "11111100", -- 3022 - 0xbce  :  252 - 0xfc
    "11111100", -- 3023 - 0xbcf  :  252 - 0xfc
    "00001111", -- 3024 - 0xbd0  :   15 - 0xf -- Background 0x7a
    "00011111", -- 3025 - 0xbd1  :   31 - 0x1f
    "00110000", -- 3026 - 0xbd2  :   48 - 0x30
    "00111000", -- 3027 - 0xbd3  :   56 - 0x38
    "00011101", -- 3028 - 0xbd4  :   29 - 0x1d
    "00000011", -- 3029 - 0xbd5  :    3 - 0x3
    "00000011", -- 3030 - 0xbd6  :    3 - 0x3
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "11111100", -- 3032 - 0xbd8  :  252 - 0xfc -- Background 0x7b
    "11111100", -- 3033 - 0xbd9  :  252 - 0xfc
    "01111100", -- 3034 - 0xbda  :  124 - 0x7c
    "10001110", -- 3035 - 0xbdb  :  142 - 0x8e
    "10000110", -- 3036 - 0xbdc  :  134 - 0x86
    "10011100", -- 3037 - 0xbdd  :  156 - 0x9c
    "01111000", -- 3038 - 0xbde  :  120 - 0x78
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Background 0x7c
    "00000001", -- 3041 - 0xbe1  :    1 - 0x1
    "00000110", -- 3042 - 0xbe2  :    6 - 0x6
    "00000111", -- 3043 - 0xbe3  :    7 - 0x7
    "00000111", -- 3044 - 0xbe4  :    7 - 0x7
    "00000111", -- 3045 - 0xbe5  :    7 - 0x7
    "00000001", -- 3046 - 0xbe6  :    1 - 0x1
    "00000011", -- 3047 - 0xbe7  :    3 - 0x3
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- Background 0x7d
    "11000000", -- 3049 - 0xbe9  :  192 - 0xc0
    "00110000", -- 3050 - 0xbea  :   48 - 0x30
    "11110000", -- 3051 - 0xbeb  :  240 - 0xf0
    "11110000", -- 3052 - 0xbec  :  240 - 0xf0
    "11110000", -- 3053 - 0xbed  :  240 - 0xf0
    "01000000", -- 3054 - 0xbee  :   64 - 0x40
    "01000000", -- 3055 - 0xbef  :   64 - 0x40
    "00000001", -- 3056 - 0xbf0  :    1 - 0x1 -- Background 0x7e
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000001", -- 3058 - 0xbf2  :    1 - 0x1
    "00000011", -- 3059 - 0xbf3  :    3 - 0x3
    "00000001", -- 3060 - 0xbf4  :    1 - 0x1
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "01000000", -- 3064 - 0xbf8  :   64 - 0x40 -- Background 0x7f
    "01000000", -- 3065 - 0xbf9  :   64 - 0x40
    "01000000", -- 3066 - 0xbfa  :   64 - 0x40
    "01000000", -- 3067 - 0xbfb  :   64 - 0x40
    "01000000", -- 3068 - 0xbfc  :   64 - 0x40
    "10000000", -- 3069 - 0xbfd  :  128 - 0x80
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0x80
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00000000", -- 3074 - 0xc02  :    0 - 0x0
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000000", -- 3076 - 0xc04  :    0 - 0x0
    "00011111", -- 3077 - 0xc05  :   31 - 0x1f
    "00010000", -- 3078 - 0xc06  :   16 - 0x10
    "00010111", -- 3079 - 0xc07  :   23 - 0x17
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- Background 0x81
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "11111111", -- 3085 - 0xc0d  :  255 - 0xff
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "11111111", -- 3087 - 0xc0f  :  255 - 0xff
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Background 0x82
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "10000000", -- 3093 - 0xc15  :  128 - 0x80
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "11000000", -- 3095 - 0xc17  :  192 - 0xc0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0 -- Background 0x83
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00001000", -- 3101 - 0xc1d  :    8 - 0x8
    "00001000", -- 3102 - 0xc1e  :    8 - 0x8
    "00010110", -- 3103 - 0xc1f  :   22 - 0x16
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0x84
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "01000000", -- 3110 - 0xc26  :   64 - 0x40
    "11000000", -- 3111 - 0xc27  :  192 - 0xc0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- Background 0x85
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000001", -- 3117 - 0xc2d  :    1 - 0x1
    "00000111", -- 3118 - 0xc2e  :    7 - 0x7
    "00001100", -- 3119 - 0xc2f  :   12 - 0xc
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0x86
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "11000000", -- 3125 - 0xc35  :  192 - 0xc0
    "00111111", -- 3126 - 0xc36  :   63 - 0x3f
    "11111111", -- 3127 - 0xc37  :  255 - 0xff
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- Background 0x87
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "11000000", -- 3135 - 0xc3f  :  192 - 0xc0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0x88
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0 -- Background 0x89
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "01000100", -- 3149 - 0xc4d  :   68 - 0x44
    "01010110", -- 3150 - 0xc4e  :   86 - 0x56
    "01011011", -- 3151 - 0xc4f  :   91 - 0x5b
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00000000", -- 3154 - 0xc52  :    0 - 0x0
    "00000000", -- 3155 - 0xc53  :    0 - 0x0
    "00000000", -- 3156 - 0xc54  :    0 - 0x0
    "00000000", -- 3157 - 0xc55  :    0 - 0x0
    "00000000", -- 3158 - 0xc56  :    0 - 0x0
    "00000000", -- 3159 - 0xc57  :    0 - 0x0
    "00000000", -- 3160 - 0xc58  :    0 - 0x0 -- Background 0x8b
    "00000000", -- 3161 - 0xc59  :    0 - 0x0
    "00000000", -- 3162 - 0xc5a  :    0 - 0x0
    "00000000", -- 3163 - 0xc5b  :    0 - 0x0
    "00000000", -- 3164 - 0xc5c  :    0 - 0x0
    "00010000", -- 3165 - 0xc5d  :   16 - 0x10
    "00110100", -- 3166 - 0xc5e  :   52 - 0x34
    "01101101", -- 3167 - 0xc5f  :  109 - 0x6d
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "00000000", -- 3174 - 0xc66  :    0 - 0x0
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0 -- Background 0x8d
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "01000000", -- 3180 - 0xc6c  :   64 - 0x40
    "01001000", -- 3181 - 0xc6d  :   72 - 0x48
    "10101000", -- 3182 - 0xc6e  :  168 - 0xa8
    "10101100", -- 3183 - 0xc6f  :  172 - 0xac
    "00000000", -- 3184 - 0xc70  :    0 - 0x0 -- Background 0x8e
    "00000000", -- 3185 - 0xc71  :    0 - 0x0
    "00000000", -- 3186 - 0xc72  :    0 - 0x0
    "00000000", -- 3187 - 0xc73  :    0 - 0x0
    "00000010", -- 3188 - 0xc74  :    2 - 0x2
    "00000010", -- 3189 - 0xc75  :    2 - 0x2
    "00000010", -- 3190 - 0xc76  :    2 - 0x2
    "00000010", -- 3191 - 0xc77  :    2 - 0x2
    "00000000", -- 3192 - 0xc78  :    0 - 0x0 -- Background 0x8f
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000011", -- 3195 - 0xc7b  :    3 - 0x3
    "01000011", -- 3196 - 0xc7c  :   67 - 0x43
    "01100010", -- 3197 - 0xc7d  :   98 - 0x62
    "10110010", -- 3198 - 0xc7e  :  178 - 0xb2
    "11011010", -- 3199 - 0xc7f  :  218 - 0xda
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "11111100", -- 3203 - 0xc83  :  252 - 0xfc
    "11111100", -- 3204 - 0xc84  :  252 - 0xfc
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "11111111", -- 3206 - 0xc86  :  255 - 0xff
    "11111111", -- 3207 - 0xc87  :  255 - 0xff
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- Background 0x91
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000000", -- 3213 - 0xc8d  :    0 - 0x0
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00010111", -- 3216 - 0xc90  :   23 - 0x17 -- Background 0x92
    "00010111", -- 3217 - 0xc91  :   23 - 0x17
    "00010111", -- 3218 - 0xc92  :   23 - 0x17
    "00010111", -- 3219 - 0xc93  :   23 - 0x17
    "00010111", -- 3220 - 0xc94  :   23 - 0x17
    "00010111", -- 3221 - 0xc95  :   23 - 0x17
    "00010111", -- 3222 - 0xc96  :   23 - 0x17
    "00010111", -- 3223 - 0xc97  :   23 - 0x17
    "11111111", -- 3224 - 0xc98  :  255 - 0xff -- Background 0x93
    "11111111", -- 3225 - 0xc99  :  255 - 0xff
    "11111111", -- 3226 - 0xc9a  :  255 - 0xff
    "11111111", -- 3227 - 0xc9b  :  255 - 0xff
    "11111001", -- 3228 - 0xc9c  :  249 - 0xf9
    "11111001", -- 3229 - 0xc9d  :  249 - 0xf9
    "11111111", -- 3230 - 0xc9e  :  255 - 0xff
    "11111111", -- 3231 - 0xc9f  :  255 - 0xff
    "11110000", -- 3232 - 0xca0  :  240 - 0xf0 -- Background 0x94
    "11111000", -- 3233 - 0xca1  :  248 - 0xf8
    "11111000", -- 3234 - 0xca2  :  248 - 0xf8
    "11111100", -- 3235 - 0xca3  :  252 - 0xfc
    "11111100", -- 3236 - 0xca4  :  252 - 0xfc
    "11111100", -- 3237 - 0xca5  :  252 - 0xfc
    "01111100", -- 3238 - 0xca6  :  124 - 0x7c
    "01111100", -- 3239 - 0xca7  :  124 - 0x7c
    "00010111", -- 3240 - 0xca8  :   23 - 0x17 -- Background 0x95
    "00101111", -- 3241 - 0xca9  :   47 - 0x2f
    "00101111", -- 3242 - 0xcaa  :   47 - 0x2f
    "01011111", -- 3243 - 0xcab  :   95 - 0x5f
    "01011111", -- 3244 - 0xcac  :   95 - 0x5f
    "10111111", -- 3245 - 0xcad  :  191 - 0xbf
    "10111111", -- 3246 - 0xcae  :  191 - 0xbf
    "01111111", -- 3247 - 0xcaf  :  127 - 0x7f
    "01100000", -- 3248 - 0xcb0  :   96 - 0x60 -- Background 0x96
    "01100000", -- 3249 - 0xcb1  :   96 - 0x60
    "10110000", -- 3250 - 0xcb2  :  176 - 0xb0
    "10110000", -- 3251 - 0xcb3  :  176 - 0xb0
    "11011000", -- 3252 - 0xcb4  :  216 - 0xd8
    "11011000", -- 3253 - 0xcb5  :  216 - 0xd8
    "11101100", -- 3254 - 0xcb6  :  236 - 0xec
    "11101100", -- 3255 - 0xcb7  :  236 - 0xec
    "00110011", -- 3256 - 0xcb8  :   51 - 0x33 -- Background 0x97
    "00101111", -- 3257 - 0xcb9  :   47 - 0x2f
    "01101111", -- 3258 - 0xcba  :  111 - 0x6f
    "01011111", -- 3259 - 0xcbb  :   95 - 0x5f
    "11011111", -- 3260 - 0xcbc  :  223 - 0xdf
    "10111111", -- 3261 - 0xcbd  :  191 - 0xbf
    "10111111", -- 3262 - 0xcbe  :  191 - 0xbf
    "10111111", -- 3263 - 0xcbf  :  191 - 0xbf
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff -- Background 0x98
    "11111111", -- 3265 - 0xcc1  :  255 - 0xff
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111110", -- 3267 - 0xcc3  :  254 - 0xfe
    "11111001", -- 3268 - 0xcc4  :  249 - 0xf9
    "11100111", -- 3269 - 0xcc5  :  231 - 0xe7
    "11111100", -- 3270 - 0xcc6  :  252 - 0xfc
    "11110011", -- 3271 - 0xcc7  :  243 - 0xf3
    "11110000", -- 3272 - 0xcc8  :  240 - 0xf0 -- Background 0x99
    "11111000", -- 3273 - 0xcc9  :  248 - 0xf8
    "11111000", -- 3274 - 0xcca  :  248 - 0xf8
    "01110000", -- 3275 - 0xccb  :  112 - 0x70
    "11001100", -- 3276 - 0xccc  :  204 - 0xcc
    "00110000", -- 3277 - 0xccd  :   48 - 0x30
    "11000000", -- 3278 - 0xcce  :  192 - 0xc0
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000000", -- 3283 - 0xcd3  :    0 - 0x0
    "00111111", -- 3284 - 0xcd4  :   63 - 0x3f
    "00100000", -- 3285 - 0xcd5  :   32 - 0x20
    "00101111", -- 3286 - 0xcd6  :   47 - 0x2f
    "00101111", -- 3287 - 0xcd7  :   47 - 0x2f
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0 -- Background 0x9b
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "11100000", -- 3292 - 0xcdc  :  224 - 0xe0
    "00000000", -- 3293 - 0xcdd  :    0 - 0x0
    "11110000", -- 3294 - 0xcde  :  240 - 0xf0
    "11110000", -- 3295 - 0xcdf  :  240 - 0xf0
    "01011101", -- 3296 - 0xce0  :   93 - 0x5d -- Background 0x9c
    "01011110", -- 3297 - 0xce1  :   94 - 0x5e
    "01011111", -- 3298 - 0xce2  :   95 - 0x5f
    "01011111", -- 3299 - 0xce3  :   95 - 0x5f
    "01011111", -- 3300 - 0xce4  :   95 - 0x5f
    "01011111", -- 3301 - 0xce5  :   95 - 0x5f
    "01011111", -- 3302 - 0xce6  :   95 - 0x5f
    "01011111", -- 3303 - 0xce7  :   95 - 0x5f
    "10000000", -- 3304 - 0xce8  :  128 - 0x80 -- Background 0x9d
    "11000001", -- 3305 - 0xce9  :  193 - 0xc1
    "01100011", -- 3306 - 0xcea  :   99 - 0x63
    "10110110", -- 3307 - 0xceb  :  182 - 0xb6
    "11011001", -- 3308 - 0xcec  :  217 - 0xd9
    "11101011", -- 3309 - 0xced  :  235 - 0xeb
    "11110111", -- 3310 - 0xcee  :  247 - 0xf7
    "11111111", -- 3311 - 0xcef  :  255 - 0xff
    "11011101", -- 3312 - 0xcf0  :  221 - 0xdd -- Background 0x9e
    "10111101", -- 3313 - 0xcf1  :  189 - 0xbd
    "01111101", -- 3314 - 0xcf2  :  125 - 0x7d
    "11111101", -- 3315 - 0xcf3  :  253 - 0xfd
    "11111101", -- 3316 - 0xcf4  :  253 - 0xfd
    "11111101", -- 3317 - 0xcf5  :  253 - 0xfd
    "11111101", -- 3318 - 0xcf6  :  253 - 0xfd
    "11111101", -- 3319 - 0xcf7  :  253 - 0xfd
    "00000001", -- 3320 - 0xcf8  :    1 - 0x1 -- Background 0x9f
    "00000001", -- 3321 - 0xcf9  :    1 - 0x1
    "00000010", -- 3322 - 0xcfa  :    2 - 0x2
    "00000010", -- 3323 - 0xcfb  :    2 - 0x2
    "00000101", -- 3324 - 0xcfc  :    5 - 0x5
    "00000101", -- 3325 - 0xcfd  :    5 - 0x5
    "00001011", -- 3326 - 0xcfe  :   11 - 0xb
    "00001011", -- 3327 - 0xcff  :   11 - 0xb
    "01110100", -- 3328 - 0xd00  :  116 - 0x74 -- Background 0xa0
    "01110110", -- 3329 - 0xd01  :  118 - 0x76
    "11111010", -- 3330 - 0xd02  :  250 - 0xfa
    "11111011", -- 3331 - 0xd03  :  251 - 0xfb
    "11111101", -- 3332 - 0xd04  :  253 - 0xfd
    "11111101", -- 3333 - 0xd05  :  253 - 0xfd
    "11111110", -- 3334 - 0xd06  :  254 - 0xfe
    "11111110", -- 3335 - 0xd07  :  254 - 0xfe
    "00000010", -- 3336 - 0xd08  :    2 - 0x2 -- Background 0xa1
    "00000010", -- 3337 - 0xd09  :    2 - 0x2
    "00000010", -- 3338 - 0xd0a  :    2 - 0x2
    "00000010", -- 3339 - 0xd0b  :    2 - 0x2
    "00000010", -- 3340 - 0xd0c  :    2 - 0x2
    "10000010", -- 3341 - 0xd0d  :  130 - 0x82
    "10000010", -- 3342 - 0xd0e  :  130 - 0x82
    "11000010", -- 3343 - 0xd0f  :  194 - 0xc2
    "11101010", -- 3344 - 0xd10  :  234 - 0xea -- Background 0xa2
    "11110110", -- 3345 - 0xd11  :  246 - 0xf6
    "11111010", -- 3346 - 0xd12  :  250 - 0xfa
    "11111010", -- 3347 - 0xd13  :  250 - 0xfa
    "11111100", -- 3348 - 0xd14  :  252 - 0xfc
    "11111100", -- 3349 - 0xd15  :  252 - 0xfc
    "11111110", -- 3350 - 0xd16  :  254 - 0xfe
    "11111111", -- 3351 - 0xd17  :  255 - 0xff
    "11111111", -- 3352 - 0xd18  :  255 - 0xff -- Background 0xa3
    "11111111", -- 3353 - 0xd19  :  255 - 0xff
    "11111111", -- 3354 - 0xd1a  :  255 - 0xff
    "11111111", -- 3355 - 0xd1b  :  255 - 0xff
    "11111111", -- 3356 - 0xd1c  :  255 - 0xff
    "11111111", -- 3357 - 0xd1d  :  255 - 0xff
    "11111111", -- 3358 - 0xd1e  :  255 - 0xff
    "11111111", -- 3359 - 0xd1f  :  255 - 0xff
    "01000000", -- 3360 - 0xd20  :   64 - 0x40 -- Background 0xa4
    "01000000", -- 3361 - 0xd21  :   64 - 0x40
    "01000000", -- 3362 - 0xd22  :   64 - 0x40
    "01000000", -- 3363 - 0xd23  :   64 - 0x40
    "01000000", -- 3364 - 0xd24  :   64 - 0x40
    "01000000", -- 3365 - 0xd25  :   64 - 0x40
    "01000000", -- 3366 - 0xd26  :   64 - 0x40
    "01000000", -- 3367 - 0xd27  :   64 - 0x40
    "11111000", -- 3368 - 0xd28  :  248 - 0xf8 -- Background 0xa5
    "11111111", -- 3369 - 0xd29  :  255 - 0xff
    "11111111", -- 3370 - 0xd2a  :  255 - 0xff
    "11111000", -- 3371 - 0xd2b  :  248 - 0xf8
    "11111011", -- 3372 - 0xd2c  :  251 - 0xfb
    "11111010", -- 3373 - 0xd2d  :  250 - 0xfa
    "11111010", -- 3374 - 0xd2e  :  250 - 0xfa
    "11111010", -- 3375 - 0xd2f  :  250 - 0xfa
    "11111100", -- 3376 - 0xd30  :  252 - 0xfc -- Background 0xa6
    "11111010", -- 3377 - 0xd31  :  250 - 0xfa
    "11110110", -- 3378 - 0xd32  :  246 - 0xf6
    "00001101", -- 3379 - 0xd33  :   13 - 0xd
    "11111001", -- 3380 - 0xd34  :  249 - 0xf9
    "00000011", -- 3381 - 0xd35  :    3 - 0x3
    "00010011", -- 3382 - 0xd36  :   19 - 0x13
    "00110111", -- 3383 - 0xd37  :   55 - 0x37
    "01111111", -- 3384 - 0xd38  :  127 - 0x7f -- Background 0xa7
    "11111001", -- 3385 - 0xd39  :  249 - 0xf9
    "11111001", -- 3386 - 0xd3a  :  249 - 0xf9
    "11111111", -- 3387 - 0xd3b  :  255 - 0xff
    "11111110", -- 3388 - 0xd3c  :  254 - 0xfe
    "11111100", -- 3389 - 0xd3d  :  252 - 0xfc
    "11111111", -- 3390 - 0xd3e  :  255 - 0xff
    "11111111", -- 3391 - 0xd3f  :  255 - 0xff
    "11110110", -- 3392 - 0xd40  :  246 - 0xf6 -- Background 0xa8
    "11110110", -- 3393 - 0xd41  :  246 - 0xf6
    "11111011", -- 3394 - 0xd42  :  251 - 0xfb
    "01111011", -- 3395 - 0xd43  :  123 - 0x7b
    "11111101", -- 3396 - 0xd44  :  253 - 0xfd
    "11110101", -- 3397 - 0xd45  :  245 - 0xf5
    "11110110", -- 3398 - 0xd46  :  246 - 0xf6
    "11111010", -- 3399 - 0xd47  :  250 - 0xfa
    "10111111", -- 3400 - 0xd48  :  191 - 0xbf -- Background 0xa9
    "10111111", -- 3401 - 0xd49  :  191 - 0xbf
    "00111111", -- 3402 - 0xd4a  :   63 - 0x3f
    "00111111", -- 3403 - 0xd4b  :   63 - 0x3f
    "10111111", -- 3404 - 0xd4c  :  191 - 0xbf
    "10011111", -- 3405 - 0xd4d  :  159 - 0x9f
    "11001111", -- 3406 - 0xd4e  :  207 - 0xcf
    "11010111", -- 3407 - 0xd4f  :  215 - 0xd7
    "11100100", -- 3408 - 0xd50  :  228 - 0xe4 -- Background 0xaa
    "11111000", -- 3409 - 0xd51  :  248 - 0xf8
    "11111111", -- 3410 - 0xd52  :  255 - 0xff
    "11110011", -- 3411 - 0xd53  :  243 - 0xf3
    "11111100", -- 3412 - 0xd54  :  252 - 0xfc
    "11111111", -- 3413 - 0xd55  :  255 - 0xff
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- Background 0xab
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "11000000", -- 3419 - 0xd5b  :  192 - 0xc0
    "11110000", -- 3420 - 0xd5c  :  240 - 0xf0
    "00111100", -- 3421 - 0xd5d  :   60 - 0x3c
    "11011000", -- 3422 - 0xd5e  :  216 - 0xd8
    "10110110", -- 3423 - 0xd5f  :  182 - 0xb6
    "00001111", -- 3424 - 0xd60  :   15 - 0xf -- Background 0xac
    "00001111", -- 3425 - 0xd61  :   15 - 0xf
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "00000011", -- 3427 - 0xd63  :    3 - 0x3
    "00000000", -- 3428 - 0xd64  :    0 - 0x0
    "00000000", -- 3429 - 0xd65  :    0 - 0x0
    "00000000", -- 3430 - 0xd66  :    0 - 0x0
    "00000000", -- 3431 - 0xd67  :    0 - 0x0
    "11110100", -- 3432 - 0xd68  :  244 - 0xf4 -- Background 0xad
    "11110100", -- 3433 - 0xd69  :  244 - 0xf4
    "00000100", -- 3434 - 0xd6a  :    4 - 0x4
    "11111100", -- 3435 - 0xd6b  :  252 - 0xfc
    "00000000", -- 3436 - 0xd6c  :    0 - 0x0
    "00000000", -- 3437 - 0xd6d  :    0 - 0x0
    "00000000", -- 3438 - 0xd6e  :    0 - 0x0
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "01011111", -- 3440 - 0xd70  :   95 - 0x5f -- Background 0xae
    "01011111", -- 3441 - 0xd71  :   95 - 0x5f
    "01011111", -- 3442 - 0xd72  :   95 - 0x5f
    "01011111", -- 3443 - 0xd73  :   95 - 0x5f
    "01011111", -- 3444 - 0xd74  :   95 - 0x5f
    "01011111", -- 3445 - 0xd75  :   95 - 0x5f
    "01011111", -- 3446 - 0xd76  :   95 - 0x5f
    "01011111", -- 3447 - 0xd77  :   95 - 0x5f
    "11111101", -- 3448 - 0xd78  :  253 - 0xfd -- Background 0xaf
    "11111101", -- 3449 - 0xd79  :  253 - 0xfd
    "11111101", -- 3450 - 0xd7a  :  253 - 0xfd
    "11111101", -- 3451 - 0xd7b  :  253 - 0xfd
    "11110101", -- 3452 - 0xd7c  :  245 - 0xf5
    "11110101", -- 3453 - 0xd7d  :  245 - 0xf5
    "11110101", -- 3454 - 0xd7e  :  245 - 0xf5
    "11110101", -- 3455 - 0xd7f  :  245 - 0xf5
    "00001100", -- 3456 - 0xd80  :   12 - 0xc -- Background 0xb0
    "00011100", -- 3457 - 0xd81  :   28 - 0x1c
    "00001100", -- 3458 - 0xd82  :   12 - 0xc
    "00001100", -- 3459 - 0xd83  :   12 - 0xc
    "00001100", -- 3460 - 0xd84  :   12 - 0xc
    "00001100", -- 3461 - 0xd85  :   12 - 0xc
    "00111111", -- 3462 - 0xd86  :   63 - 0x3f
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00111110", -- 3464 - 0xd88  :   62 - 0x3e -- Background 0xb1
    "01100011", -- 3465 - 0xd89  :   99 - 0x63
    "00000111", -- 3466 - 0xd8a  :    7 - 0x7
    "00011110", -- 3467 - 0xd8b  :   30 - 0x1e
    "00111100", -- 3468 - 0xd8c  :   60 - 0x3c
    "01110000", -- 3469 - 0xd8d  :  112 - 0x70
    "01111111", -- 3470 - 0xd8e  :  127 - 0x7f
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "01111110", -- 3472 - 0xd90  :  126 - 0x7e -- Background 0xb2
    "01100011", -- 3473 - 0xd91  :   99 - 0x63
    "01100011", -- 3474 - 0xd92  :   99 - 0x63
    "01100011", -- 3475 - 0xd93  :   99 - 0x63
    "01111110", -- 3476 - 0xd94  :  126 - 0x7e
    "01100000", -- 3477 - 0xd95  :   96 - 0x60
    "01100000", -- 3478 - 0xd96  :   96 - 0x60
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "01100011", -- 3480 - 0xd98  :   99 - 0x63 -- Background 0xb3
    "01100011", -- 3481 - 0xd99  :   99 - 0x63
    "01100011", -- 3482 - 0xd9a  :   99 - 0x63
    "01100011", -- 3483 - 0xd9b  :   99 - 0x63
    "01100011", -- 3484 - 0xd9c  :   99 - 0x63
    "01100011", -- 3485 - 0xd9d  :   99 - 0x63
    "00111110", -- 3486 - 0xd9e  :   62 - 0x3e
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "01100011", -- 3488 - 0xda0  :   99 - 0x63 -- Background 0xb4
    "01100011", -- 3489 - 0xda1  :   99 - 0x63
    "01100011", -- 3490 - 0xda2  :   99 - 0x63
    "01111111", -- 3491 - 0xda3  :  127 - 0x7f
    "01100011", -- 3492 - 0xda4  :   99 - 0x63
    "01100011", -- 3493 - 0xda5  :   99 - 0x63
    "01100011", -- 3494 - 0xda6  :   99 - 0x63
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00111111", -- 3496 - 0xda8  :   63 - 0x3f -- Background 0xb5
    "00001100", -- 3497 - 0xda9  :   12 - 0xc
    "00001100", -- 3498 - 0xdaa  :   12 - 0xc
    "00001100", -- 3499 - 0xdab  :   12 - 0xc
    "00001100", -- 3500 - 0xdac  :   12 - 0xc
    "00001100", -- 3501 - 0xdad  :   12 - 0xc
    "00111111", -- 3502 - 0xdae  :   63 - 0x3f
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 3505 - 0xdb1  :    0 - 0x0
    "00000000", -- 3506 - 0xdb2  :    0 - 0x0
    "01111110", -- 3507 - 0xdb3  :  126 - 0x7e
    "00000000", -- 3508 - 0xdb4  :    0 - 0x0
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000000", -- 3510 - 0xdb6  :    0 - 0x0
    "00000000", -- 3511 - 0xdb7  :    0 - 0x0
    "00111100", -- 3512 - 0xdb8  :   60 - 0x3c -- Background 0xb7
    "01100110", -- 3513 - 0xdb9  :  102 - 0x66
    "01100000", -- 3514 - 0xdba  :   96 - 0x60
    "00111110", -- 3515 - 0xdbb  :   62 - 0x3e
    "00000011", -- 3516 - 0xdbc  :    3 - 0x3
    "01100011", -- 3517 - 0xdbd  :   99 - 0x63
    "00111110", -- 3518 - 0xdbe  :   62 - 0x3e
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00011110", -- 3520 - 0xdc0  :   30 - 0x1e -- Background 0xb8
    "00110011", -- 3521 - 0xdc1  :   51 - 0x33
    "01100000", -- 3522 - 0xdc2  :   96 - 0x60
    "01100000", -- 3523 - 0xdc3  :   96 - 0x60
    "01100000", -- 3524 - 0xdc4  :   96 - 0x60
    "00110011", -- 3525 - 0xdc5  :   51 - 0x33
    "00011110", -- 3526 - 0xdc6  :   30 - 0x1e
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "00111110", -- 3528 - 0xdc8  :   62 - 0x3e -- Background 0xb9
    "01100011", -- 3529 - 0xdc9  :   99 - 0x63
    "01100011", -- 3530 - 0xdca  :   99 - 0x63
    "01100011", -- 3531 - 0xdcb  :   99 - 0x63
    "01100011", -- 3532 - 0xdcc  :   99 - 0x63
    "01100011", -- 3533 - 0xdcd  :   99 - 0x63
    "00111110", -- 3534 - 0xdce  :   62 - 0x3e
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "01111110", -- 3536 - 0xdd0  :  126 - 0x7e -- Background 0xba
    "01100011", -- 3537 - 0xdd1  :   99 - 0x63
    "01100011", -- 3538 - 0xdd2  :   99 - 0x63
    "01100111", -- 3539 - 0xdd3  :  103 - 0x67
    "01111100", -- 3540 - 0xdd4  :  124 - 0x7c
    "01101110", -- 3541 - 0xdd5  :  110 - 0x6e
    "01100111", -- 3542 - 0xdd6  :  103 - 0x67
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "01111111", -- 3544 - 0xdd8  :  127 - 0x7f -- Background 0xbb
    "01100000", -- 3545 - 0xdd9  :   96 - 0x60
    "01100000", -- 3546 - 0xdda  :   96 - 0x60
    "01111110", -- 3547 - 0xddb  :  126 - 0x7e
    "01100000", -- 3548 - 0xddc  :   96 - 0x60
    "01100000", -- 3549 - 0xddd  :   96 - 0x60
    "01111111", -- 3550 - 0xdde  :  127 - 0x7f
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00000000", -- 3552 - 0xde0  :    0 - 0x0 -- Background 0xbc
    "00000000", -- 3553 - 0xde1  :    0 - 0x0
    "00000000", -- 3554 - 0xde2  :    0 - 0x0
    "00000000", -- 3555 - 0xde3  :    0 - 0x0
    "00000000", -- 3556 - 0xde4  :    0 - 0x0
    "00000000", -- 3557 - 0xde5  :    0 - 0x0
    "00000000", -- 3558 - 0xde6  :    0 - 0x0
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "00000000", -- 3560 - 0xde8  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 3561 - 0xde9  :    0 - 0x0
    "00000000", -- 3562 - 0xdea  :    0 - 0x0
    "00000000", -- 3563 - 0xdeb  :    0 - 0x0
    "00000000", -- 3564 - 0xdec  :    0 - 0x0
    "00000000", -- 3565 - 0xded  :    0 - 0x0
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "00000000", -- 3568 - 0xdf0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 3569 - 0xdf1  :    0 - 0x0
    "00000000", -- 3570 - 0xdf2  :    0 - 0x0
    "00000000", -- 3571 - 0xdf3  :    0 - 0x0
    "00000000", -- 3572 - 0xdf4  :    0 - 0x0
    "00000000", -- 3573 - 0xdf5  :    0 - 0x0
    "00000000", -- 3574 - 0xdf6  :    0 - 0x0
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "01100011", -- 3584 - 0xe00  :   99 - 0x63 -- Background 0xc0
    "01100110", -- 3585 - 0xe01  :  102 - 0x66
    "01101100", -- 3586 - 0xe02  :  108 - 0x6c
    "01111000", -- 3587 - 0xe03  :  120 - 0x78
    "01111100", -- 3588 - 0xe04  :  124 - 0x7c
    "01100110", -- 3589 - 0xe05  :  102 - 0x66
    "01100011", -- 3590 - 0xe06  :   99 - 0x63
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00111111", -- 3592 - 0xe08  :   63 - 0x3f -- Background 0xc1
    "00001100", -- 3593 - 0xe09  :   12 - 0xc
    "00001100", -- 3594 - 0xe0a  :   12 - 0xc
    "00001100", -- 3595 - 0xe0b  :   12 - 0xc
    "00001100", -- 3596 - 0xe0c  :   12 - 0xc
    "00001100", -- 3597 - 0xe0d  :   12 - 0xc
    "00111111", -- 3598 - 0xe0e  :   63 - 0x3f
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "01100011", -- 3600 - 0xe10  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 3601 - 0xe11  :  119 - 0x77
    "01111111", -- 3602 - 0xe12  :  127 - 0x7f
    "01111111", -- 3603 - 0xe13  :  127 - 0x7f
    "01101011", -- 3604 - 0xe14  :  107 - 0x6b
    "01100011", -- 3605 - 0xe15  :   99 - 0x63
    "01100011", -- 3606 - 0xe16  :   99 - 0x63
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00011100", -- 3608 - 0xe18  :   28 - 0x1c -- Background 0xc3
    "00110110", -- 3609 - 0xe19  :   54 - 0x36
    "01100011", -- 3610 - 0xe1a  :   99 - 0x63
    "01100011", -- 3611 - 0xe1b  :   99 - 0x63
    "01111111", -- 3612 - 0xe1c  :  127 - 0x7f
    "01100011", -- 3613 - 0xe1d  :   99 - 0x63
    "01100011", -- 3614 - 0xe1e  :   99 - 0x63
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00011111", -- 3616 - 0xe20  :   31 - 0x1f -- Background 0xc4
    "00110000", -- 3617 - 0xe21  :   48 - 0x30
    "01100000", -- 3618 - 0xe22  :   96 - 0x60
    "01100111", -- 3619 - 0xe23  :  103 - 0x67
    "01100011", -- 3620 - 0xe24  :   99 - 0x63
    "00110011", -- 3621 - 0xe25  :   51 - 0x33
    "00011111", -- 3622 - 0xe26  :   31 - 0x1f
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "01100011", -- 3624 - 0xe28  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 3625 - 0xe29  :   99 - 0x63
    "01100011", -- 3626 - 0xe2a  :   99 - 0x63
    "01100011", -- 3627 - 0xe2b  :   99 - 0x63
    "01100011", -- 3628 - 0xe2c  :   99 - 0x63
    "01100011", -- 3629 - 0xe2d  :   99 - 0x63
    "00111110", -- 3630 - 0xe2e  :   62 - 0x3e
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "01111110", -- 3632 - 0xe30  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 3633 - 0xe31  :   99 - 0x63
    "01100011", -- 3634 - 0xe32  :   99 - 0x63
    "01100111", -- 3635 - 0xe33  :  103 - 0x67
    "01111100", -- 3636 - 0xe34  :  124 - 0x7c
    "01101110", -- 3637 - 0xe35  :  110 - 0x6e
    "01100111", -- 3638 - 0xe36  :  103 - 0x67
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "01111111", -- 3640 - 0xe38  :  127 - 0x7f -- Background 0xc7
    "01100000", -- 3641 - 0xe39  :   96 - 0x60
    "01100000", -- 3642 - 0xe3a  :   96 - 0x60
    "01111110", -- 3643 - 0xe3b  :  126 - 0x7e
    "01100000", -- 3644 - 0xe3c  :   96 - 0x60
    "01100000", -- 3645 - 0xe3d  :   96 - 0x60
    "01111111", -- 3646 - 0xe3e  :  127 - 0x7f
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00110110", -- 3648 - 0xe40  :   54 - 0x36 -- Background 0xc8
    "00110110", -- 3649 - 0xe41  :   54 - 0x36
    "00010010", -- 3650 - 0xe42  :   18 - 0x12
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00111110", -- 3656 - 0xe48  :   62 - 0x3e -- Background 0xc9
    "01100011", -- 3657 - 0xe49  :   99 - 0x63
    "01100011", -- 3658 - 0xe4a  :   99 - 0x63
    "01100011", -- 3659 - 0xe4b  :   99 - 0x63
    "01100011", -- 3660 - 0xe4c  :   99 - 0x63
    "01100011", -- 3661 - 0xe4d  :   99 - 0x63
    "00111110", -- 3662 - 0xe4e  :   62 - 0x3e
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00111100", -- 3664 - 0xe50  :   60 - 0x3c -- Background 0xca
    "01100110", -- 3665 - 0xe51  :  102 - 0x66
    "01100000", -- 3666 - 0xe52  :   96 - 0x60
    "00111110", -- 3667 - 0xe53  :   62 - 0x3e
    "00000011", -- 3668 - 0xe54  :    3 - 0x3
    "01100011", -- 3669 - 0xe55  :   99 - 0x63
    "00111110", -- 3670 - 0xe56  :   62 - 0x3e
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- Background 0xcb
    "00111000", -- 3673 - 0xe59  :   56 - 0x38
    "01111100", -- 3674 - 0xe5a  :  124 - 0x7c
    "11111110", -- 3675 - 0xe5b  :  254 - 0xfe
    "11111110", -- 3676 - 0xe5c  :  254 - 0xfe
    "11111110", -- 3677 - 0xe5d  :  254 - 0xfe
    "01111100", -- 3678 - 0xe5e  :  124 - 0x7c
    "00111000", -- 3679 - 0xe5f  :   56 - 0x38
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "00000000", -- 3685 - 0xe65  :    0 - 0x0
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "00000000", -- 3691 - 0xe6b  :    0 - 0x0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "00000000", -- 3702 - 0xe76  :    0 - 0x0
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00000000", -- 3704 - 0xe78  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00010111", -- 3712 - 0xe80  :   23 - 0x17 -- Background 0xd0
    "00010111", -- 3713 - 0xe81  :   23 - 0x17
    "00101111", -- 3714 - 0xe82  :   47 - 0x2f
    "00101111", -- 3715 - 0xe83  :   47 - 0x2f
    "01011111", -- 3716 - 0xe84  :   95 - 0x5f
    "01011111", -- 3717 - 0xe85  :   95 - 0x5f
    "00111111", -- 3718 - 0xe86  :   63 - 0x3f
    "00111111", -- 3719 - 0xe87  :   63 - 0x3f
    "11111111", -- 3720 - 0xe88  :  255 - 0xff -- Background 0xd1
    "11001111", -- 3721 - 0xe89  :  207 - 0xcf
    "11001111", -- 3722 - 0xe8a  :  207 - 0xcf
    "11111011", -- 3723 - 0xe8b  :  251 - 0xfb
    "11110111", -- 3724 - 0xe8c  :  247 - 0xf7
    "11100111", -- 3725 - 0xe8d  :  231 - 0xe7
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "01000010", -- 3728 - 0xe90  :   66 - 0x42 -- Background 0xd2
    "01100010", -- 3729 - 0xe91  :   98 - 0x62
    "10100010", -- 3730 - 0xe92  :  162 - 0xa2
    "10110010", -- 3731 - 0xe93  :  178 - 0xb2
    "01010010", -- 3732 - 0xe94  :   82 - 0x52
    "01011010", -- 3733 - 0xe95  :   90 - 0x5a
    "10101010", -- 3734 - 0xe96  :  170 - 0xaa
    "10101100", -- 3735 - 0xe97  :  172 - 0xac
    "11111111", -- 3736 - 0xe98  :  255 - 0xff -- Background 0xd3
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111101", -- 3740 - 0xe9c  :  253 - 0xfd
    "11111101", -- 3741 - 0xe9d  :  253 - 0xfd
    "11111101", -- 3742 - 0xe9e  :  253 - 0xfd
    "11111101", -- 3743 - 0xe9f  :  253 - 0xfd
    "00000111", -- 3744 - 0xea0  :    7 - 0x7 -- Background 0xd4
    "00000111", -- 3745 - 0xea1  :    7 - 0x7
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000011", -- 3747 - 0xea3  :    3 - 0x3
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "11111010", -- 3752 - 0xea8  :  250 - 0xfa -- Background 0xd5
    "11111010", -- 3753 - 0xea9  :  250 - 0xfa
    "00000010", -- 3754 - 0xeaa  :    2 - 0x2
    "11111110", -- 3755 - 0xeab  :  254 - 0xfe
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00001111", -- 3760 - 0xeb0  :   15 - 0xf -- Background 0xd6
    "00001111", -- 3761 - 0xeb1  :   15 - 0xf
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "00000111", -- 3763 - 0xeb3  :    7 - 0x7
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "00000000", -- 3770 - 0xeba  :    0 - 0x0
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "11000011", -- 3776 - 0xec0  :  195 - 0xc3 -- Background 0xd8
    "11111111", -- 3777 - 0xec1  :  255 - 0xff
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "11111111", -- 3779 - 0xec3  :  255 - 0xff
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "01101011", -- 3784 - 0xec8  :  107 - 0x6b -- Background 0xd9
    "10110101", -- 3785 - 0xec9  :  181 - 0xb5
    "00110110", -- 3786 - 0xeca  :   54 - 0x36
    "11111000", -- 3787 - 0xecb  :  248 - 0xf8
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "11111111", -- 3792 - 0xed0  :  255 - 0xff -- Background 0xda
    "11111111", -- 3793 - 0xed1  :  255 - 0xff
    "01111110", -- 3794 - 0xed2  :  126 - 0x7e
    "10000001", -- 3795 - 0xed3  :  129 - 0x81
    "00011111", -- 3796 - 0xed4  :   31 - 0x1f
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "01101100", -- 3800 - 0xed8  :  108 - 0x6c -- Background 0xdb
    "11011000", -- 3801 - 0xed9  :  216 - 0xd8
    "00110000", -- 3802 - 0xeda  :   48 - 0x30
    "11100000", -- 3803 - 0xedb  :  224 - 0xe0
    "10000000", -- 3804 - 0xedc  :  128 - 0x80
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00011111", -- 3808 - 0xee0  :   31 - 0x1f -- Background 0xdc
    "00011111", -- 3809 - 0xee1  :   31 - 0x1f
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000111", -- 3811 - 0xee3  :    7 - 0x7
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "10000101", -- 3816 - 0xee8  :  133 - 0x85 -- Background 0xdd
    "11111101", -- 3817 - 0xee9  :  253 - 0xfd
    "00000001", -- 3818 - 0xeea  :    1 - 0x1
    "11111111", -- 3819 - 0xeeb  :  255 - 0xff
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "01111111", -- 3824 - 0xef0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 3825 - 0xef1  :  127 - 0x7f
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "01011111", -- 3827 - 0xef3  :   95 - 0x5f
    "00000000", -- 3828 - 0xef4  :    0 - 0x0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "00000000", -- 3830 - 0xef6  :    0 - 0x0
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "11111100", -- 3832 - 0xef8  :  252 - 0xfc -- Background 0xdf
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00110100", -- 3840 - 0xf00  :   52 - 0x34 -- Background 0xe0
    "11110110", -- 3841 - 0xf01  :  246 - 0xf6
    "00000010", -- 3842 - 0xf02  :    2 - 0x2
    "11111111", -- 3843 - 0xf03  :  255 - 0xff
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "11111111", -- 3848 - 0xf08  :  255 - 0xff -- Background 0xe1
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "01111111", -- 3851 - 0xf0b  :  127 - 0x7f
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "11100001", -- 3856 - 0xf10  :  225 - 0xe1 -- Background 0xe2
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "01000000", -- 3864 - 0xf18  :   64 - 0x40 -- Background 0xe3
    "01000000", -- 3865 - 0xf19  :   64 - 0x40
    "01000000", -- 3866 - 0xf1a  :   64 - 0x40
    "11000000", -- 3867 - 0xf1b  :  192 - 0xc0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000111", -- 3876 - 0xf24  :    7 - 0x7
    "00001111", -- 3877 - 0xf25  :   15 - 0xf
    "00001111", -- 3878 - 0xf26  :   15 - 0xf
    "00001111", -- 3879 - 0xf27  :   15 - 0xf
    "00000000", -- 3880 - 0xf28  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "11100000", -- 3884 - 0xf2c  :  224 - 0xe0
    "11110000", -- 3885 - 0xf2d  :  240 - 0xf0
    "11110000", -- 3886 - 0xf2e  :  240 - 0xf0
    "11110000", -- 3887 - 0xf2f  :  240 - 0xf0
    "11110000", -- 3888 - 0xf30  :  240 - 0xf0 -- Background 0xe6
    "11110000", -- 3889 - 0xf31  :  240 - 0xf0
    "11110000", -- 3890 - 0xf32  :  240 - 0xf0
    "11100000", -- 3891 - 0xf33  :  224 - 0xe0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00001111", -- 3896 - 0xf38  :   15 - 0xf -- Background 0xe7
    "00001111", -- 3897 - 0xf39  :   15 - 0xf
    "00001111", -- 3898 - 0xf3a  :   15 - 0xf
    "00000111", -- 3899 - 0xf3b  :    7 - 0x7
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "11111111", -- 3908 - 0xf44  :  255 - 0xff
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "11110000", -- 3912 - 0xf48  :  240 - 0xf0 -- Background 0xe9
    "11110000", -- 3913 - 0xf49  :  240 - 0xf0
    "11110000", -- 3914 - 0xf4a  :  240 - 0xf0
    "11110000", -- 3915 - 0xf4b  :  240 - 0xf0
    "11110000", -- 3916 - 0xf4c  :  240 - 0xf0
    "11110000", -- 3917 - 0xf4d  :  240 - 0xf0
    "11110000", -- 3918 - 0xf4e  :  240 - 0xf0
    "11110000", -- 3919 - 0xf4f  :  240 - 0xf0
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Background 0xea
    "11111111", -- 3921 - 0xf51  :  255 - 0xff
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "11111111", -- 3923 - 0xf53  :  255 - 0xff
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00001111", -- 3928 - 0xf58  :   15 - 0xf -- Background 0xeb
    "00001111", -- 3929 - 0xf59  :   15 - 0xf
    "00001111", -- 3930 - 0xf5a  :   15 - 0xf
    "00001111", -- 3931 - 0xf5b  :   15 - 0xf
    "00001111", -- 3932 - 0xf5c  :   15 - 0xf
    "00001111", -- 3933 - 0xf5d  :   15 - 0xf
    "00001111", -- 3934 - 0xf5e  :   15 - 0xf
    "00001111", -- 3935 - 0xf5f  :   15 - 0xf
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- Background 0xed
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0 -- Background 0xef
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "11111111", -- 3968 - 0xf80  :  255 - 0xff -- Background 0xf0
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "11111111", -- 3970 - 0xf82  :  255 - 0xff
    "11111111", -- 3971 - 0xf83  :  255 - 0xff
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "11111111", -- 3974 - 0xf86  :  255 - 0xff
    "11111111", -- 3975 - 0xf87  :  255 - 0xff
    "11111111", -- 3976 - 0xf88  :  255 - 0xff -- Background 0xf1
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111111", -- 3982 - 0xf8e  :  255 - 0xff
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Background 0xf2
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "11111111", -- 3992 - 0xf98  :  255 - 0xff -- Background 0xf3
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111111", -- 3999 - 0xf9f  :  255 - 0xff
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Background 0xf4
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "11111111", -- 4007 - 0xfa7  :  255 - 0xff
    "11111111", -- 4008 - 0xfa8  :  255 - 0xff -- Background 0xf5
    "11111111", -- 4009 - 0xfa9  :  255 - 0xff
    "11111111", -- 4010 - 0xfaa  :  255 - 0xff
    "11111111", -- 4011 - 0xfab  :  255 - 0xff
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "11111111", -- 4015 - 0xfaf  :  255 - 0xff
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Background 0xf6
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "11111111", -- 4024 - 0xfb8  :  255 - 0xff -- Background 0xf7
    "11111111", -- 4025 - 0xfb9  :  255 - 0xff
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "11111111", -- 4031 - 0xfbf  :  255 - 0xff
    "11111111", -- 4032 - 0xfc0  :  255 - 0xff -- Background 0xf8
    "11111111", -- 4033 - 0xfc1  :  255 - 0xff
    "11111111", -- 4034 - 0xfc2  :  255 - 0xff
    "11111111", -- 4035 - 0xfc3  :  255 - 0xff
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "11111111", -- 4040 - 0xfc8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 4041 - 0xfc9  :  255 - 0xff
    "11111111", -- 4042 - 0xfca  :  255 - 0xff
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "11111111", -- 4048 - 0xfd0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 4049 - 0xfd1  :  255 - 0xff
    "11111111", -- 4050 - 0xfd2  :  255 - 0xff
    "11111111", -- 4051 - 0xfd3  :  255 - 0xff
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff -- Background 0xfb
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "11111111", -- 4064 - 0xfe0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 4065 - 0xfe1  :  255 - 0xff
    "11111111", -- 4066 - 0xfe2  :  255 - 0xff
    "11111111", -- 4067 - 0xfe3  :  255 - 0xff
    "11111111", -- 4068 - 0xfe4  :  255 - 0xff
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff -- Background 0xfd
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11111111", -- 4075 - 0xfeb  :  255 - 0xff
    "11111111", -- 4076 - 0xfec  :  255 - 0xff
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff -- Background 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
