//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: smario_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_color0
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout  = 8'b00000011; //    0 :   3 - 0x3 -- Sprite 0x0
      12'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      12'h2: dout  = 8'b00011111; //    2 :  31 - 0x1f
      12'h3: dout  = 8'b00011111; //    3 :  31 - 0x1f
      12'h4: dout  = 8'b00011100; //    4 :  28 - 0x1c
      12'h5: dout  = 8'b00100100; //    5 :  36 - 0x24
      12'h6: dout  = 8'b00100110; //    6 :  38 - 0x26
      12'h7: dout  = 8'b01100110; //    7 : 102 - 0x66
      12'h8: dout  = 8'b11100000; //    8 : 224 - 0xe0 -- Sprite 0x1
      12'h9: dout  = 8'b11000000; //    9 : 192 - 0xc0
      12'hA: dout  = 8'b10000000; //   10 : 128 - 0x80
      12'hB: dout  = 8'b11111100; //   11 : 252 - 0xfc
      12'hC: dout  = 8'b10000000; //   12 : 128 - 0x80
      12'hD: dout  = 8'b11000000; //   13 : 192 - 0xc0
      12'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout  = 8'b00100000; //   15 :  32 - 0x20
      12'h10: dout  = 8'b01100000; //   16 :  96 - 0x60 -- Sprite 0x2
      12'h11: dout  = 8'b01110000; //   17 : 112 - 0x70
      12'h12: dout  = 8'b00011000; //   18 :  24 - 0x18
      12'h13: dout  = 8'b00000111; //   19 :   7 - 0x7
      12'h14: dout  = 8'b00001111; //   20 :  15 - 0xf
      12'h15: dout  = 8'b00011111; //   21 :  31 - 0x1f
      12'h16: dout  = 8'b00111111; //   22 :  63 - 0x3f
      12'h17: dout  = 8'b01111111; //   23 : 127 - 0x7f
      12'h18: dout  = 8'b11111100; //   24 : 252 - 0xfc -- Sprite 0x3
      12'h19: dout  = 8'b01111100; //   25 : 124 - 0x7c
      12'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout  = 8'b11100000; //   28 : 224 - 0xe0
      12'h1D: dout  = 8'b11110000; //   29 : 240 - 0xf0
      12'h1E: dout  = 8'b11111000; //   30 : 248 - 0xf8
      12'h1F: dout  = 8'b11111000; //   31 : 248 - 0xf8
      12'h20: dout  = 8'b01111111; //   32 : 127 - 0x7f -- Sprite 0x4
      12'h21: dout  = 8'b01111111; //   33 : 127 - 0x7f
      12'h22: dout  = 8'b11111111; //   34 : 255 - 0xff
      12'h23: dout  = 8'b11111111; //   35 : 255 - 0xff
      12'h24: dout  = 8'b00000111; //   36 :   7 - 0x7
      12'h25: dout  = 8'b00000111; //   37 :   7 - 0x7
      12'h26: dout  = 8'b00001111; //   38 :  15 - 0xf
      12'h27: dout  = 8'b00001111; //   39 :  15 - 0xf
      12'h28: dout  = 8'b11111101; //   40 : 253 - 0xfd -- Sprite 0x5
      12'h29: dout  = 8'b11111110; //   41 : 254 - 0xfe
      12'h2A: dout  = 8'b10110100; //   42 : 180 - 0xb4
      12'h2B: dout  = 8'b11111000; //   43 : 248 - 0xf8
      12'h2C: dout  = 8'b11111000; //   44 : 248 - 0xf8
      12'h2D: dout  = 8'b11111001; //   45 : 249 - 0xf9
      12'h2E: dout  = 8'b11111011; //   46 : 251 - 0xfb
      12'h2F: dout  = 8'b11111111; //   47 : 255 - 0xff
      12'h30: dout  = 8'b00011111; //   48 :  31 - 0x1f -- Sprite 0x6
      12'h31: dout  = 8'b00111111; //   49 :  63 - 0x3f
      12'h32: dout  = 8'b11111111; //   50 : 255 - 0xff
      12'h33: dout  = 8'b11111111; //   51 : 255 - 0xff
      12'h34: dout  = 8'b11111100; //   52 : 252 - 0xfc
      12'h35: dout  = 8'b01110000; //   53 : 112 - 0x70
      12'h36: dout  = 8'b01110000; //   54 : 112 - 0x70
      12'h37: dout  = 8'b00111000; //   55 :  56 - 0x38
      12'h38: dout  = 8'b11111111; //   56 : 255 - 0xff -- Sprite 0x7
      12'h39: dout  = 8'b11111111; //   57 : 255 - 0xff
      12'h3A: dout  = 8'b11111111; //   58 : 255 - 0xff
      12'h3B: dout  = 8'b00011111; //   59 :  31 - 0x1f
      12'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      12'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      12'h42: dout  = 8'b00000001; //   66 :   1 - 0x1
      12'h43: dout  = 8'b00000111; //   67 :   7 - 0x7
      12'h44: dout  = 8'b00001111; //   68 :  15 - 0xf
      12'h45: dout  = 8'b00001111; //   69 :  15 - 0xf
      12'h46: dout  = 8'b00001110; //   70 :  14 - 0xe
      12'h47: dout  = 8'b00010010; //   71 :  18 - 0x12
      12'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      12'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout  = 8'b11110000; //   74 : 240 - 0xf0
      12'h4B: dout  = 8'b11100000; //   75 : 224 - 0xe0
      12'h4C: dout  = 8'b11000000; //   76 : 192 - 0xc0
      12'h4D: dout  = 8'b11111110; //   77 : 254 - 0xfe
      12'h4E: dout  = 8'b01000000; //   78 :  64 - 0x40
      12'h4F: dout  = 8'b01100000; //   79 :  96 - 0x60
      12'h50: dout  = 8'b00010011; //   80 :  19 - 0x13 -- Sprite 0xa
      12'h51: dout  = 8'b00110011; //   81 :  51 - 0x33
      12'h52: dout  = 8'b00110000; //   82 :  48 - 0x30
      12'h53: dout  = 8'b00011000; //   83 :  24 - 0x18
      12'h54: dout  = 8'b00000100; //   84 :   4 - 0x4
      12'h55: dout  = 8'b00001111; //   85 :  15 - 0xf
      12'h56: dout  = 8'b00011111; //   86 :  31 - 0x1f
      12'h57: dout  = 8'b00011111; //   87 :  31 - 0x1f
      12'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- Sprite 0xb
      12'h59: dout  = 8'b00010000; //   89 :  16 - 0x10
      12'h5A: dout  = 8'b01111110; //   90 : 126 - 0x7e
      12'h5B: dout  = 8'b00111110; //   91 :  62 - 0x3e
      12'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout  = 8'b11000000; //   94 : 192 - 0xc0
      12'h5F: dout  = 8'b11100000; //   95 : 224 - 0xe0
      12'h60: dout  = 8'b00111111; //   96 :  63 - 0x3f -- Sprite 0xc
      12'h61: dout  = 8'b00111111; //   97 :  63 - 0x3f
      12'h62: dout  = 8'b00111111; //   98 :  63 - 0x3f
      12'h63: dout  = 8'b00011111; //   99 :  31 - 0x1f
      12'h64: dout  = 8'b00011111; //  100 :  31 - 0x1f
      12'h65: dout  = 8'b00011111; //  101 :  31 - 0x1f
      12'h66: dout  = 8'b00011111; //  102 :  31 - 0x1f
      12'h67: dout  = 8'b00011111; //  103 :  31 - 0x1f
      12'h68: dout  = 8'b11110000; //  104 : 240 - 0xf0 -- Sprite 0xd
      12'h69: dout  = 8'b11110000; //  105 : 240 - 0xf0
      12'h6A: dout  = 8'b11110000; //  106 : 240 - 0xf0
      12'h6B: dout  = 8'b11111000; //  107 : 248 - 0xf8
      12'h6C: dout  = 8'b11111000; //  108 : 248 - 0xf8
      12'h6D: dout  = 8'b11111000; //  109 : 248 - 0xf8
      12'h6E: dout  = 8'b11111000; //  110 : 248 - 0xf8
      12'h6F: dout  = 8'b11111000; //  111 : 248 - 0xf8
      12'h70: dout  = 8'b11111111; //  112 : 255 - 0xff -- Sprite 0xe
      12'h71: dout  = 8'b11111111; //  113 : 255 - 0xff
      12'h72: dout  = 8'b11111111; //  114 : 255 - 0xff
      12'h73: dout  = 8'b11111110; //  115 : 254 - 0xfe
      12'h74: dout  = 8'b11110000; //  116 : 240 - 0xf0
      12'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      12'h76: dout  = 8'b10000000; //  118 : 128 - 0x80
      12'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout  = 8'b11111100; //  120 : 252 - 0xfc -- Sprite 0xf
      12'h79: dout  = 8'b11111100; //  121 : 252 - 0xfc
      12'h7A: dout  = 8'b11111000; //  122 : 248 - 0xf8
      12'h7B: dout  = 8'b01111000; //  123 : 120 - 0x78
      12'h7C: dout  = 8'b01111000; //  124 : 120 - 0x78
      12'h7D: dout  = 8'b01111000; //  125 : 120 - 0x78
      12'h7E: dout  = 8'b01111110; //  126 : 126 - 0x7e
      12'h7F: dout  = 8'b01111110; //  127 : 126 - 0x7e
      12'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout  = 8'b00000011; //  129 :   3 - 0x3
      12'h82: dout  = 8'b00001111; //  130 :  15 - 0xf
      12'h83: dout  = 8'b00011111; //  131 :  31 - 0x1f
      12'h84: dout  = 8'b00011111; //  132 :  31 - 0x1f
      12'h85: dout  = 8'b00011100; //  133 :  28 - 0x1c
      12'h86: dout  = 8'b00100100; //  134 :  36 - 0x24
      12'h87: dout  = 8'b00100110; //  135 :  38 - 0x26
      12'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      12'h89: dout  = 8'b11100000; //  137 : 224 - 0xe0
      12'h8A: dout  = 8'b11000000; //  138 : 192 - 0xc0
      12'h8B: dout  = 8'b10000000; //  139 : 128 - 0x80
      12'h8C: dout  = 8'b11111100; //  140 : 252 - 0xfc
      12'h8D: dout  = 8'b10000000; //  141 : 128 - 0x80
      12'h8E: dout  = 8'b11000000; //  142 : 192 - 0xc0
      12'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout  = 8'b01100110; //  144 : 102 - 0x66 -- Sprite 0x12
      12'h91: dout  = 8'b01100000; //  145 :  96 - 0x60
      12'h92: dout  = 8'b00110000; //  146 :  48 - 0x30
      12'h93: dout  = 8'b00011000; //  147 :  24 - 0x18
      12'h94: dout  = 8'b00001111; //  148 :  15 - 0xf
      12'h95: dout  = 8'b00011111; //  149 :  31 - 0x1f
      12'h96: dout  = 8'b00111111; //  150 :  63 - 0x3f
      12'h97: dout  = 8'b00111111; //  151 :  63 - 0x3f
      12'h98: dout  = 8'b00100000; //  152 :  32 - 0x20 -- Sprite 0x13
      12'h99: dout  = 8'b11111100; //  153 : 252 - 0xfc
      12'h9A: dout  = 8'b01111100; //  154 : 124 - 0x7c
      12'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout  = 8'b11100000; //  157 : 224 - 0xe0
      12'h9E: dout  = 8'b11100000; //  158 : 224 - 0xe0
      12'h9F: dout  = 8'b11110000; //  159 : 240 - 0xf0
      12'hA0: dout  = 8'b00111111; //  160 :  63 - 0x3f -- Sprite 0x14
      12'hA1: dout  = 8'b00111111; //  161 :  63 - 0x3f
      12'hA2: dout  = 8'b00111111; //  162 :  63 - 0x3f
      12'hA3: dout  = 8'b00111111; //  163 :  63 - 0x3f
      12'hA4: dout  = 8'b00111111; //  164 :  63 - 0x3f
      12'hA5: dout  = 8'b00111111; //  165 :  63 - 0x3f
      12'hA6: dout  = 8'b00111111; //  166 :  63 - 0x3f
      12'hA7: dout  = 8'b00011111; //  167 :  31 - 0x1f
      12'hA8: dout  = 8'b11110000; //  168 : 240 - 0xf0 -- Sprite 0x15
      12'hA9: dout  = 8'b10010000; //  169 : 144 - 0x90
      12'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout  = 8'b00001000; //  171 :   8 - 0x8
      12'hAC: dout  = 8'b00001100; //  172 :  12 - 0xc
      12'hAD: dout  = 8'b00011100; //  173 :  28 - 0x1c
      12'hAE: dout  = 8'b11111100; //  174 : 252 - 0xfc
      12'hAF: dout  = 8'b11111000; //  175 : 248 - 0xf8
      12'hB0: dout  = 8'b00001111; //  176 :  15 - 0xf -- Sprite 0x16
      12'hB1: dout  = 8'b00001111; //  177 :  15 - 0xf
      12'hB2: dout  = 8'b00000111; //  178 :   7 - 0x7
      12'hB3: dout  = 8'b00000111; //  179 :   7 - 0x7
      12'hB4: dout  = 8'b00000111; //  180 :   7 - 0x7
      12'hB5: dout  = 8'b00001111; //  181 :  15 - 0xf
      12'hB6: dout  = 8'b00001111; //  182 :  15 - 0xf
      12'hB7: dout  = 8'b00000011; //  183 :   3 - 0x3
      12'hB8: dout  = 8'b11111000; //  184 : 248 - 0xf8 -- Sprite 0x17
      12'hB9: dout  = 8'b11110000; //  185 : 240 - 0xf0
      12'hBA: dout  = 8'b11100000; //  186 : 224 - 0xe0
      12'hBB: dout  = 8'b11110000; //  187 : 240 - 0xf0
      12'hBC: dout  = 8'b10110000; //  188 : 176 - 0xb0
      12'hBD: dout  = 8'b10000000; //  189 : 128 - 0x80
      12'hBE: dout  = 8'b11100000; //  190 : 224 - 0xe0
      12'hBF: dout  = 8'b11100000; //  191 : 224 - 0xe0
      12'hC0: dout  = 8'b00000011; //  192 :   3 - 0x3 -- Sprite 0x18
      12'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      12'hC2: dout  = 8'b01111111; //  194 : 127 - 0x7f
      12'hC3: dout  = 8'b00011001; //  195 :  25 - 0x19
      12'hC4: dout  = 8'b00001001; //  196 :   9 - 0x9
      12'hC5: dout  = 8'b00001001; //  197 :   9 - 0x9
      12'hC6: dout  = 8'b00101000; //  198 :  40 - 0x28
      12'hC7: dout  = 8'b01011100; //  199 :  92 - 0x5c
      12'hC8: dout  = 8'b11111000; //  200 : 248 - 0xf8 -- Sprite 0x19
      12'hC9: dout  = 8'b11100000; //  201 : 224 - 0xe0
      12'hCA: dout  = 8'b11100000; //  202 : 224 - 0xe0
      12'hCB: dout  = 8'b11111100; //  203 : 252 - 0xfc
      12'hCC: dout  = 8'b00100110; //  204 :  38 - 0x26
      12'hCD: dout  = 8'b00110000; //  205 :  48 - 0x30
      12'hCE: dout  = 8'b10000000; //  206 : 128 - 0x80
      12'hCF: dout  = 8'b00010000; //  207 :  16 - 0x10
      12'hD0: dout  = 8'b00111110; //  208 :  62 - 0x3e -- Sprite 0x1a
      12'hD1: dout  = 8'b00011110; //  209 :  30 - 0x1e
      12'hD2: dout  = 8'b00111111; //  210 :  63 - 0x3f
      12'hD3: dout  = 8'b00111000; //  211 :  56 - 0x38
      12'hD4: dout  = 8'b00110000; //  212 :  48 - 0x30
      12'hD5: dout  = 8'b00110000; //  213 :  48 - 0x30
      12'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout  = 8'b00111010; //  215 :  58 - 0x3a
      12'hD8: dout  = 8'b01111000; //  216 : 120 - 0x78 -- Sprite 0x1b
      12'hD9: dout  = 8'b00011110; //  217 :  30 - 0x1e
      12'hDA: dout  = 8'b10000000; //  218 : 128 - 0x80
      12'hDB: dout  = 8'b11111110; //  219 : 254 - 0xfe
      12'hDC: dout  = 8'b01111110; //  220 : 126 - 0x7e
      12'hDD: dout  = 8'b01111110; //  221 : 126 - 0x7e
      12'hDE: dout  = 8'b01111111; //  222 : 127 - 0x7f
      12'hDF: dout  = 8'b01111111; //  223 : 127 - 0x7f
      12'hE0: dout  = 8'b00111100; //  224 :  60 - 0x3c -- Sprite 0x1c
      12'hE1: dout  = 8'b00111111; //  225 :  63 - 0x3f
      12'hE2: dout  = 8'b00011111; //  226 :  31 - 0x1f
      12'hE3: dout  = 8'b00001111; //  227 :  15 - 0xf
      12'hE4: dout  = 8'b00000111; //  228 :   7 - 0x7
      12'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      12'hE6: dout  = 8'b00100001; //  230 :  33 - 0x21
      12'hE7: dout  = 8'b00100000; //  231 :  32 - 0x20
      12'hE8: dout  = 8'b11111111; //  232 : 255 - 0xff -- Sprite 0x1d
      12'hE9: dout  = 8'b11111111; //  233 : 255 - 0xff
      12'hEA: dout  = 8'b11111111; //  234 : 255 - 0xff
      12'hEB: dout  = 8'b11111110; //  235 : 254 - 0xfe
      12'hEC: dout  = 8'b11111110; //  236 : 254 - 0xfe
      12'hED: dout  = 8'b11111110; //  237 : 254 - 0xfe
      12'hEE: dout  = 8'b11111100; //  238 : 252 - 0xfc
      12'hEF: dout  = 8'b01110000; //  239 : 112 - 0x70
      12'hF0: dout  = 8'b00001111; //  240 :  15 - 0xf -- Sprite 0x1e
      12'hF1: dout  = 8'b10011111; //  241 : 159 - 0x9f
      12'hF2: dout  = 8'b11001111; //  242 : 207 - 0xcf
      12'hF3: dout  = 8'b11111111; //  243 : 255 - 0xff
      12'hF4: dout  = 8'b01111111; //  244 : 127 - 0x7f
      12'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      12'hF6: dout  = 8'b00011110; //  246 :  30 - 0x1e
      12'hF7: dout  = 8'b00001110; //  247 :  14 - 0xe
      12'hF8: dout  = 8'b00100000; //  248 :  32 - 0x20 -- Sprite 0x1f
      12'hF9: dout  = 8'b11000000; //  249 : 192 - 0xc0
      12'hFA: dout  = 8'b10000000; //  250 : 128 - 0x80
      12'hFB: dout  = 8'b10000000; //  251 : 128 - 0x80
      12'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout  = 8'b00000011; //  258 :   3 - 0x3
      12'h103: dout  = 8'b00001111; //  259 :  15 - 0xf
      12'h104: dout  = 8'b00011111; //  260 :  31 - 0x1f
      12'h105: dout  = 8'b00011111; //  261 :  31 - 0x1f
      12'h106: dout  = 8'b00011100; //  262 :  28 - 0x1c
      12'h107: dout  = 8'b00100100; //  263 :  36 - 0x24
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout  = 8'b00000100; //  265 :   4 - 0x4
      12'h10A: dout  = 8'b11100110; //  266 : 230 - 0xe6
      12'h10B: dout  = 8'b11100000; //  267 : 224 - 0xe0
      12'h10C: dout  = 8'b11111111; //  268 : 255 - 0xff
      12'h10D: dout  = 8'b11111111; //  269 : 255 - 0xff
      12'h10E: dout  = 8'b10001111; //  270 : 143 - 0x8f
      12'h10F: dout  = 8'b10000011; //  271 : 131 - 0x83
      12'h110: dout  = 8'b00100110; //  272 :  38 - 0x26 -- Sprite 0x22
      12'h111: dout  = 8'b00100110; //  273 :  38 - 0x26
      12'h112: dout  = 8'b01100000; //  274 :  96 - 0x60
      12'h113: dout  = 8'b01111000; //  275 : 120 - 0x78
      12'h114: dout  = 8'b00011000; //  276 :  24 - 0x18
      12'h115: dout  = 8'b00001111; //  277 :  15 - 0xf
      12'h116: dout  = 8'b01111111; //  278 : 127 - 0x7f
      12'h117: dout  = 8'b11111111; //  279 : 255 - 0xff
      12'h118: dout  = 8'b00000001; //  280 :   1 - 0x1 -- Sprite 0x23
      12'h119: dout  = 8'b00100001; //  281 :  33 - 0x21
      12'h11A: dout  = 8'b11111110; //  282 : 254 - 0xfe
      12'h11B: dout  = 8'b01111010; //  283 : 122 - 0x7a
      12'h11C: dout  = 8'b00000110; //  284 :   6 - 0x6
      12'h11D: dout  = 8'b11111110; //  285 : 254 - 0xfe
      12'h11E: dout  = 8'b11111100; //  286 : 252 - 0xfc
      12'h11F: dout  = 8'b11111100; //  287 : 252 - 0xfc
      12'h120: dout  = 8'b11111111; //  288 : 255 - 0xff -- Sprite 0x24
      12'h121: dout  = 8'b11001111; //  289 : 207 - 0xcf
      12'h122: dout  = 8'b10000111; //  290 : 135 - 0x87
      12'h123: dout  = 8'b00000111; //  291 :   7 - 0x7
      12'h124: dout  = 8'b00000111; //  292 :   7 - 0x7
      12'h125: dout  = 8'b00001111; //  293 :  15 - 0xf
      12'h126: dout  = 8'b00011111; //  294 :  31 - 0x1f
      12'h127: dout  = 8'b00011111; //  295 :  31 - 0x1f
      12'h128: dout  = 8'b11111000; //  296 : 248 - 0xf8 -- Sprite 0x25
      12'h129: dout  = 8'b11111000; //  297 : 248 - 0xf8
      12'h12A: dout  = 8'b11110000; //  298 : 240 - 0xf0
      12'h12B: dout  = 8'b10111000; //  299 : 184 - 0xb8
      12'h12C: dout  = 8'b11111000; //  300 : 248 - 0xf8
      12'h12D: dout  = 8'b11111001; //  301 : 249 - 0xf9
      12'h12E: dout  = 8'b11111011; //  302 : 251 - 0xfb
      12'h12F: dout  = 8'b11111111; //  303 : 255 - 0xff
      12'h130: dout  = 8'b00011111; //  304 :  31 - 0x1f -- Sprite 0x26
      12'h131: dout  = 8'b11111111; //  305 : 255 - 0xff
      12'h132: dout  = 8'b11111111; //  306 : 255 - 0xff
      12'h133: dout  = 8'b11111111; //  307 : 255 - 0xff
      12'h134: dout  = 8'b11111111; //  308 : 255 - 0xff
      12'h135: dout  = 8'b11111110; //  309 : 254 - 0xfe
      12'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      12'h137: dout  = 8'b10000000; //  311 : 128 - 0x80
      12'h138: dout  = 8'b11111111; //  312 : 255 - 0xff -- Sprite 0x27
      12'h139: dout  = 8'b11111111; //  313 : 255 - 0xff
      12'h13A: dout  = 8'b11111111; //  314 : 255 - 0xff
      12'h13B: dout  = 8'b00111111; //  315 :  63 - 0x3f
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b00010011; //  320 :  19 - 0x13 -- Sprite 0x28
      12'h141: dout  = 8'b00110011; //  321 :  51 - 0x33
      12'h142: dout  = 8'b00110000; //  322 :  48 - 0x30
      12'h143: dout  = 8'b00011000; //  323 :  24 - 0x18
      12'h144: dout  = 8'b00000100; //  324 :   4 - 0x4
      12'h145: dout  = 8'b00001111; //  325 :  15 - 0xf
      12'h146: dout  = 8'b00011111; //  326 :  31 - 0x1f
      12'h147: dout  = 8'b00011111; //  327 :  31 - 0x1f
      12'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Sprite 0x29
      12'h149: dout  = 8'b00010000; //  329 :  16 - 0x10
      12'h14A: dout  = 8'b01111110; //  330 : 126 - 0x7e
      12'h14B: dout  = 8'b00110000; //  331 :  48 - 0x30
      12'h14C: dout  = 8'b11100000; //  332 : 224 - 0xe0
      12'h14D: dout  = 8'b11110000; //  333 : 240 - 0xf0
      12'h14E: dout  = 8'b11110000; //  334 : 240 - 0xf0
      12'h14F: dout  = 8'b11100000; //  335 : 224 - 0xe0
      12'h150: dout  = 8'b00011111; //  336 :  31 - 0x1f -- Sprite 0x2a
      12'h151: dout  = 8'b00011111; //  337 :  31 - 0x1f
      12'h152: dout  = 8'b00001111; //  338 :  15 - 0xf
      12'h153: dout  = 8'b00001111; //  339 :  15 - 0xf
      12'h154: dout  = 8'b00001111; //  340 :  15 - 0xf
      12'h155: dout  = 8'b00011111; //  341 :  31 - 0x1f
      12'h156: dout  = 8'b00011111; //  342 :  31 - 0x1f
      12'h157: dout  = 8'b00011111; //  343 :  31 - 0x1f
      12'h158: dout  = 8'b11110000; //  344 : 240 - 0xf0 -- Sprite 0x2b
      12'h159: dout  = 8'b11110000; //  345 : 240 - 0xf0
      12'h15A: dout  = 8'b11111000; //  346 : 248 - 0xf8
      12'h15B: dout  = 8'b11111000; //  347 : 248 - 0xf8
      12'h15C: dout  = 8'b10111000; //  348 : 184 - 0xb8
      12'h15D: dout  = 8'b11111000; //  349 : 248 - 0xf8
      12'h15E: dout  = 8'b11111000; //  350 : 248 - 0xf8
      12'h15F: dout  = 8'b11111000; //  351 : 248 - 0xf8
      12'h160: dout  = 8'b00111111; //  352 :  63 - 0x3f -- Sprite 0x2c
      12'h161: dout  = 8'b11111111; //  353 : 255 - 0xff
      12'h162: dout  = 8'b11111111; //  354 : 255 - 0xff
      12'h163: dout  = 8'b11111111; //  355 : 255 - 0xff
      12'h164: dout  = 8'b11110110; //  356 : 246 - 0xf6
      12'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      12'h166: dout  = 8'b10000100; //  358 : 132 - 0x84
      12'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout  = 8'b11110000; //  360 : 240 - 0xf0 -- Sprite 0x2d
      12'h169: dout  = 8'b11100000; //  361 : 224 - 0xe0
      12'h16A: dout  = 8'b10000000; //  362 : 128 - 0x80
      12'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout  = 8'b00011111; //  368 :  31 - 0x1f -- Sprite 0x2e
      12'h171: dout  = 8'b00011111; //  369 :  31 - 0x1f
      12'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      12'h173: dout  = 8'b00111111; //  371 :  63 - 0x3f
      12'h174: dout  = 8'b00011111; //  372 :  31 - 0x1f
      12'h175: dout  = 8'b00001111; //  373 :  15 - 0xf
      12'h176: dout  = 8'b00001111; //  374 :  15 - 0xf
      12'h177: dout  = 8'b00011111; //  375 :  31 - 0x1f
      12'h178: dout  = 8'b11110000; //  376 : 240 - 0xf0 -- Sprite 0x2f
      12'h179: dout  = 8'b11110000; //  377 : 240 - 0xf0
      12'h17A: dout  = 8'b11111000; //  378 : 248 - 0xf8
      12'h17B: dout  = 8'b11111000; //  379 : 248 - 0xf8
      12'h17C: dout  = 8'b10111000; //  380 : 184 - 0xb8
      12'h17D: dout  = 8'b11111000; //  381 : 248 - 0xf8
      12'h17E: dout  = 8'b11111000; //  382 : 248 - 0xf8
      12'h17F: dout  = 8'b11110000; //  383 : 240 - 0xf0
      12'h180: dout  = 8'b11100000; //  384 : 224 - 0xe0 -- Sprite 0x30
      12'h181: dout  = 8'b11110000; //  385 : 240 - 0xf0
      12'h182: dout  = 8'b11110000; //  386 : 240 - 0xf0
      12'h183: dout  = 8'b11110000; //  387 : 240 - 0xf0
      12'h184: dout  = 8'b11110000; //  388 : 240 - 0xf0
      12'h185: dout  = 8'b11110000; //  389 : 240 - 0xf0
      12'h186: dout  = 8'b11111000; //  390 : 248 - 0xf8
      12'h187: dout  = 8'b11110000; //  391 : 240 - 0xf0
      12'h188: dout  = 8'b00011111; //  392 :  31 - 0x1f -- Sprite 0x31
      12'h189: dout  = 8'b00011111; //  393 :  31 - 0x1f
      12'h18A: dout  = 8'b00011111; //  394 :  31 - 0x1f
      12'h18B: dout  = 8'b00111111; //  395 :  63 - 0x3f
      12'h18C: dout  = 8'b00111110; //  396 :  62 - 0x3e
      12'h18D: dout  = 8'b00111100; //  397 :  60 - 0x3c
      12'h18E: dout  = 8'b00111000; //  398 :  56 - 0x38
      12'h18F: dout  = 8'b00011000; //  399 :  24 - 0x18
      12'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      12'h191: dout  = 8'b00000011; //  401 :   3 - 0x3
      12'h192: dout  = 8'b00000111; //  402 :   7 - 0x7
      12'h193: dout  = 8'b00000111; //  403 :   7 - 0x7
      12'h194: dout  = 8'b00001010; //  404 :  10 - 0xa
      12'h195: dout  = 8'b00001011; //  405 :  11 - 0xb
      12'h196: dout  = 8'b00001100; //  406 :  12 - 0xc
      12'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      12'h199: dout  = 8'b11100000; //  409 : 224 - 0xe0
      12'h19A: dout  = 8'b11111100; //  410 : 252 - 0xfc
      12'h19B: dout  = 8'b00100000; //  411 :  32 - 0x20
      12'h19C: dout  = 8'b00100000; //  412 :  32 - 0x20
      12'h19D: dout  = 8'b00010000; //  413 :  16 - 0x10
      12'h19E: dout  = 8'b00111100; //  414 :  60 - 0x3c
      12'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout  = 8'b00000111; //  416 :   7 - 0x7 -- Sprite 0x34
      12'h1A1: dout  = 8'b00000111; //  417 :   7 - 0x7
      12'h1A2: dout  = 8'b00000111; //  418 :   7 - 0x7
      12'h1A3: dout  = 8'b00011111; //  419 :  31 - 0x1f
      12'h1A4: dout  = 8'b00011111; //  420 :  31 - 0x1f
      12'h1A5: dout  = 8'b00111110; //  421 :  62 - 0x3e
      12'h1A6: dout  = 8'b00100001; //  422 :  33 - 0x21
      12'h1A7: dout  = 8'b00000001; //  423 :   1 - 0x1
      12'h1A8: dout  = 8'b11100000; //  424 : 224 - 0xe0 -- Sprite 0x35
      12'h1A9: dout  = 8'b11100000; //  425 : 224 - 0xe0
      12'h1AA: dout  = 8'b11100000; //  426 : 224 - 0xe0
      12'h1AB: dout  = 8'b11110000; //  427 : 240 - 0xf0
      12'h1AC: dout  = 8'b11110000; //  428 : 240 - 0xf0
      12'h1AD: dout  = 8'b11100000; //  429 : 224 - 0xe0
      12'h1AE: dout  = 8'b11000000; //  430 : 192 - 0xc0
      12'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      12'h1B0: dout  = 8'b00000111; //  432 :   7 - 0x7 -- Sprite 0x36
      12'h1B1: dout  = 8'b00001111; //  433 :  15 - 0xf
      12'h1B2: dout  = 8'b00001110; //  434 :  14 - 0xe
      12'h1B3: dout  = 8'b00010100; //  435 :  20 - 0x14
      12'h1B4: dout  = 8'b00010110; //  436 :  22 - 0x16
      12'h1B5: dout  = 8'b00011000; //  437 :  24 - 0x18
      12'h1B6: dout  = 8'b00000000; //  438 :   0 - 0x0
      12'h1B7: dout  = 8'b00111111; //  439 :  63 - 0x3f
      12'h1B8: dout  = 8'b11000000; //  440 : 192 - 0xc0 -- Sprite 0x37
      12'h1B9: dout  = 8'b11111000; //  441 : 248 - 0xf8
      12'h1BA: dout  = 8'b01000000; //  442 :  64 - 0x40
      12'h1BB: dout  = 8'b01000000; //  443 :  64 - 0x40
      12'h1BC: dout  = 8'b00100000; //  444 :  32 - 0x20
      12'h1BD: dout  = 8'b01111000; //  445 : 120 - 0x78
      12'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout  = 8'b11000000; //  447 : 192 - 0xc0
      12'h1C0: dout  = 8'b00111111; //  448 :  63 - 0x3f -- Sprite 0x38
      12'h1C1: dout  = 8'b00001110; //  449 :  14 - 0xe
      12'h1C2: dout  = 8'b00001111; //  450 :  15 - 0xf
      12'h1C3: dout  = 8'b00011111; //  451 :  31 - 0x1f
      12'h1C4: dout  = 8'b00111111; //  452 :  63 - 0x3f
      12'h1C5: dout  = 8'b01111100; //  453 : 124 - 0x7c
      12'h1C6: dout  = 8'b01110000; //  454 : 112 - 0x70
      12'h1C7: dout  = 8'b00111000; //  455 :  56 - 0x38
      12'h1C8: dout  = 8'b11110000; //  456 : 240 - 0xf0 -- Sprite 0x39
      12'h1C9: dout  = 8'b11111000; //  457 : 248 - 0xf8
      12'h1CA: dout  = 8'b11100100; //  458 : 228 - 0xe4
      12'h1CB: dout  = 8'b11111100; //  459 : 252 - 0xfc
      12'h1CC: dout  = 8'b11111100; //  460 : 252 - 0xfc
      12'h1CD: dout  = 8'b01111100; //  461 : 124 - 0x7c
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b00000111; //  464 :   7 - 0x7 -- Sprite 0x3a
      12'h1D1: dout  = 8'b00001111; //  465 :  15 - 0xf
      12'h1D2: dout  = 8'b00001110; //  466 :  14 - 0xe
      12'h1D3: dout  = 8'b00010100; //  467 :  20 - 0x14
      12'h1D4: dout  = 8'b00010110; //  468 :  22 - 0x16
      12'h1D5: dout  = 8'b00011000; //  469 :  24 - 0x18
      12'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout  = 8'b00001111; //  471 :  15 - 0xf
      12'h1D8: dout  = 8'b00011111; //  472 :  31 - 0x1f -- Sprite 0x3b
      12'h1D9: dout  = 8'b00011111; //  473 :  31 - 0x1f
      12'h1DA: dout  = 8'b00011111; //  474 :  31 - 0x1f
      12'h1DB: dout  = 8'b00011100; //  475 :  28 - 0x1c
      12'h1DC: dout  = 8'b00001100; //  476 :  12 - 0xc
      12'h1DD: dout  = 8'b00000111; //  477 :   7 - 0x7
      12'h1DE: dout  = 8'b00000111; //  478 :   7 - 0x7
      12'h1DF: dout  = 8'b00000111; //  479 :   7 - 0x7
      12'h1E0: dout  = 8'b11100000; //  480 : 224 - 0xe0 -- Sprite 0x3c
      12'h1E1: dout  = 8'b01100000; //  481 :  96 - 0x60
      12'h1E2: dout  = 8'b11110000; //  482 : 240 - 0xf0
      12'h1E3: dout  = 8'b01110000; //  483 : 112 - 0x70
      12'h1E4: dout  = 8'b11100000; //  484 : 224 - 0xe0
      12'h1E5: dout  = 8'b11100000; //  485 : 224 - 0xe0
      12'h1E6: dout  = 8'b11110000; //  486 : 240 - 0xf0
      12'h1E7: dout  = 8'b10000000; //  487 : 128 - 0x80
      12'h1E8: dout  = 8'b00000111; //  488 :   7 - 0x7 -- Sprite 0x3d
      12'h1E9: dout  = 8'b00011111; //  489 :  31 - 0x1f
      12'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      12'h1EB: dout  = 8'b00010010; //  491 :  18 - 0x12
      12'h1EC: dout  = 8'b00010011; //  492 :  19 - 0x13
      12'h1ED: dout  = 8'b00001000; //  493 :   8 - 0x8
      12'h1EE: dout  = 8'b00011111; //  494 :  31 - 0x1f
      12'h1EF: dout  = 8'b00110001; //  495 :  49 - 0x31
      12'h1F0: dout  = 8'b11000000; //  496 : 192 - 0xc0 -- Sprite 0x3e
      12'h1F1: dout  = 8'b11110000; //  497 : 240 - 0xf0
      12'h1F2: dout  = 8'b01000000; //  498 :  64 - 0x40
      12'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      12'h1F4: dout  = 8'b00110000; //  500 :  48 - 0x30
      12'h1F5: dout  = 8'b00011000; //  501 :  24 - 0x18
      12'h1F6: dout  = 8'b11000000; //  502 : 192 - 0xc0
      12'h1F7: dout  = 8'b11111000; //  503 : 248 - 0xf8
      12'h1F8: dout  = 8'b00110001; //  504 :  49 - 0x31 -- Sprite 0x3f
      12'h1F9: dout  = 8'b00111001; //  505 :  57 - 0x39
      12'h1FA: dout  = 8'b00011111; //  506 :  31 - 0x1f
      12'h1FB: dout  = 8'b00011111; //  507 :  31 - 0x1f
      12'h1FC: dout  = 8'b00001111; //  508 :  15 - 0xf
      12'h1FD: dout  = 8'b01011111; //  509 :  95 - 0x5f
      12'h1FE: dout  = 8'b01111110; //  510 : 126 - 0x7e
      12'h1FF: dout  = 8'b00111100; //  511 :  60 - 0x3c
      12'h200: dout  = 8'b11111000; //  512 : 248 - 0xf8 -- Sprite 0x40
      12'h201: dout  = 8'b11111000; //  513 : 248 - 0xf8
      12'h202: dout  = 8'b11110000; //  514 : 240 - 0xf0
      12'h203: dout  = 8'b11100000; //  515 : 224 - 0xe0
      12'h204: dout  = 8'b11100000; //  516 : 224 - 0xe0
      12'h205: dout  = 8'b11000000; //  517 : 192 - 0xc0
      12'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      12'h209: dout  = 8'b11100000; //  521 : 224 - 0xe0
      12'h20A: dout  = 8'b11111100; //  522 : 252 - 0xfc
      12'h20B: dout  = 8'b00100111; //  523 :  39 - 0x27
      12'h20C: dout  = 8'b00100111; //  524 :  39 - 0x27
      12'h20D: dout  = 8'b00010001; //  525 :  17 - 0x11
      12'h20E: dout  = 8'b00111110; //  526 :  62 - 0x3e
      12'h20F: dout  = 8'b00000100; //  527 :   4 - 0x4
      12'h210: dout  = 8'b00111111; //  528 :  63 - 0x3f -- Sprite 0x42
      12'h211: dout  = 8'b01111111; //  529 : 127 - 0x7f
      12'h212: dout  = 8'b00111111; //  530 :  63 - 0x3f
      12'h213: dout  = 8'b00001111; //  531 :  15 - 0xf
      12'h214: dout  = 8'b00011111; //  532 :  31 - 0x1f
      12'h215: dout  = 8'b00111111; //  533 :  63 - 0x3f
      12'h216: dout  = 8'b01111111; //  534 : 127 - 0x7f
      12'h217: dout  = 8'b01001111; //  535 :  79 - 0x4f
      12'h218: dout  = 8'b11111000; //  536 : 248 - 0xf8 -- Sprite 0x43
      12'h219: dout  = 8'b11111001; //  537 : 249 - 0xf9
      12'h21A: dout  = 8'b11111001; //  538 : 249 - 0xf9
      12'h21B: dout  = 8'b10110111; //  539 : 183 - 0xb7
      12'h21C: dout  = 8'b11111111; //  540 : 255 - 0xff
      12'h21D: dout  = 8'b11111111; //  541 : 255 - 0xff
      12'h21E: dout  = 8'b11100000; //  542 : 224 - 0xe0
      12'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout  = 8'b00000111; //  544 :   7 - 0x7 -- Sprite 0x44
      12'h221: dout  = 8'b00000111; //  545 :   7 - 0x7
      12'h222: dout  = 8'b00001111; //  546 :  15 - 0xf
      12'h223: dout  = 8'b00111111; //  547 :  63 - 0x3f
      12'h224: dout  = 8'b00111111; //  548 :  63 - 0x3f
      12'h225: dout  = 8'b00111111; //  549 :  63 - 0x3f
      12'h226: dout  = 8'b00100110; //  550 :  38 - 0x26
      12'h227: dout  = 8'b00000100; //  551 :   4 - 0x4
      12'h228: dout  = 8'b11110000; //  552 : 240 - 0xf0 -- Sprite 0x45
      12'h229: dout  = 8'b11110000; //  553 : 240 - 0xf0
      12'h22A: dout  = 8'b11110000; //  554 : 240 - 0xf0
      12'h22B: dout  = 8'b11100000; //  555 : 224 - 0xe0
      12'h22C: dout  = 8'b11000000; //  556 : 192 - 0xc0
      12'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout  = 8'b00000111; //  560 :   7 - 0x7 -- Sprite 0x46
      12'h231: dout  = 8'b00000111; //  561 :   7 - 0x7
      12'h232: dout  = 8'b00001111; //  562 :  15 - 0xf
      12'h233: dout  = 8'b00011111; //  563 :  31 - 0x1f
      12'h234: dout  = 8'b00111111; //  564 :  63 - 0x3f
      12'h235: dout  = 8'b00001111; //  565 :  15 - 0xf
      12'h236: dout  = 8'b00011100; //  566 :  28 - 0x1c
      12'h237: dout  = 8'b00011000; //  567 :  24 - 0x18
      12'h238: dout  = 8'b11100000; //  568 : 224 - 0xe0 -- Sprite 0x47
      12'h239: dout  = 8'b11100000; //  569 : 224 - 0xe0
      12'h23A: dout  = 8'b11100000; //  570 : 224 - 0xe0
      12'h23B: dout  = 8'b11100000; //  571 : 224 - 0xe0
      12'h23C: dout  = 8'b11000000; //  572 : 192 - 0xc0
      12'h23D: dout  = 8'b10000000; //  573 : 128 - 0x80
      12'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout  = 8'b00000111; //  576 :   7 - 0x7 -- Sprite 0x48
      12'h241: dout  = 8'b00001111; //  577 :  15 - 0xf
      12'h242: dout  = 8'b00011111; //  578 :  31 - 0x1f
      12'h243: dout  = 8'b00001111; //  579 :  15 - 0xf
      12'h244: dout  = 8'b00111111; //  580 :  63 - 0x3f
      12'h245: dout  = 8'b00001111; //  581 :  15 - 0xf
      12'h246: dout  = 8'b00011100; //  582 :  28 - 0x1c
      12'h247: dout  = 8'b00011000; //  583 :  24 - 0x18
      12'h248: dout  = 8'b11100000; //  584 : 224 - 0xe0 -- Sprite 0x49
      12'h249: dout  = 8'b11100000; //  585 : 224 - 0xe0
      12'h24A: dout  = 8'b11100000; //  586 : 224 - 0xe0
      12'h24B: dout  = 8'b01000000; //  587 :  64 - 0x40
      12'h24C: dout  = 8'b11000000; //  588 : 192 - 0xc0
      12'h24D: dout  = 8'b10000000; //  589 : 128 - 0x80
      12'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b01111111; //  592 : 127 - 0x7f -- Sprite 0x4a
      12'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      12'h252: dout  = 8'b11111111; //  594 : 255 - 0xff
      12'h253: dout  = 8'b11111011; //  595 : 251 - 0xfb
      12'h254: dout  = 8'b00001111; //  596 :  15 - 0xf
      12'h255: dout  = 8'b00001111; //  597 :  15 - 0xf
      12'h256: dout  = 8'b00001111; //  598 :  15 - 0xf
      12'h257: dout  = 8'b00011111; //  599 :  31 - 0x1f
      12'h258: dout  = 8'b00111111; //  600 :  63 - 0x3f -- Sprite 0x4b
      12'h259: dout  = 8'b01111110; //  601 : 126 - 0x7e
      12'h25A: dout  = 8'b01111100; //  602 : 124 - 0x7c
      12'h25B: dout  = 8'b01111100; //  603 : 124 - 0x7c
      12'h25C: dout  = 8'b00111100; //  604 :  60 - 0x3c
      12'h25D: dout  = 8'b00111100; //  605 :  60 - 0x3c
      12'h25E: dout  = 8'b11111100; //  606 : 252 - 0xfc
      12'h25F: dout  = 8'b11111100; //  607 : 252 - 0xfc
      12'h260: dout  = 8'b01100000; //  608 :  96 - 0x60 -- Sprite 0x4c
      12'h261: dout  = 8'b01110000; //  609 : 112 - 0x70
      12'h262: dout  = 8'b00011000; //  610 :  24 - 0x18
      12'h263: dout  = 8'b00001000; //  611 :   8 - 0x8
      12'h264: dout  = 8'b00001111; //  612 :  15 - 0xf
      12'h265: dout  = 8'b00011111; //  613 :  31 - 0x1f
      12'h266: dout  = 8'b00111111; //  614 :  63 - 0x3f
      12'h267: dout  = 8'b01111111; //  615 : 127 - 0x7f
      12'h268: dout  = 8'b11111100; //  616 : 252 - 0xfc -- Sprite 0x4d
      12'h269: dout  = 8'b01111100; //  617 : 124 - 0x7c
      12'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout  = 8'b00100000; //  619 :  32 - 0x20
      12'h26C: dout  = 8'b11110000; //  620 : 240 - 0xf0
      12'h26D: dout  = 8'b11111000; //  621 : 248 - 0xf8
      12'h26E: dout  = 8'b11111100; //  622 : 252 - 0xfc
      12'h26F: dout  = 8'b11111110; //  623 : 254 - 0xfe
      12'h270: dout  = 8'b00001011; //  624 :  11 - 0xb -- Sprite 0x4e
      12'h271: dout  = 8'b00001111; //  625 :  15 - 0xf
      12'h272: dout  = 8'b00011111; //  626 :  31 - 0x1f
      12'h273: dout  = 8'b00011110; //  627 :  30 - 0x1e
      12'h274: dout  = 8'b00111100; //  628 :  60 - 0x3c
      12'h275: dout  = 8'b00111100; //  629 :  60 - 0x3c
      12'h276: dout  = 8'b00111100; //  630 :  60 - 0x3c
      12'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      12'h278: dout  = 8'b00011111; //  632 :  31 - 0x1f -- Sprite 0x4f
      12'h279: dout  = 8'b00111111; //  633 :  63 - 0x3f
      12'h27A: dout  = 8'b00001101; //  634 :  13 - 0xd
      12'h27B: dout  = 8'b00000111; //  635 :   7 - 0x7
      12'h27C: dout  = 8'b00001111; //  636 :  15 - 0xf
      12'h27D: dout  = 8'b00001110; //  637 :  14 - 0xe
      12'h27E: dout  = 8'b00011100; //  638 :  28 - 0x1c
      12'h27F: dout  = 8'b00111100; //  639 :  60 - 0x3c
      12'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      12'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      12'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout  = 8'b00000111; //  649 :   7 - 0x7
      12'h28A: dout  = 8'b00011111; //  650 :  31 - 0x1f
      12'h28B: dout  = 8'b11111111; //  651 : 255 - 0xff
      12'h28C: dout  = 8'b00000111; //  652 :   7 - 0x7
      12'h28D: dout  = 8'b00011111; //  653 :  31 - 0x1f
      12'h28E: dout  = 8'b00001111; //  654 :  15 - 0xf
      12'h28F: dout  = 8'b00000110; //  655 :   6 - 0x6
      12'h290: dout  = 8'b00111111; //  656 :  63 - 0x3f -- Sprite 0x52
      12'h291: dout  = 8'b11111111; //  657 : 255 - 0xff
      12'h292: dout  = 8'b11111111; //  658 : 255 - 0xff
      12'h293: dout  = 8'b11111111; //  659 : 255 - 0xff
      12'h294: dout  = 8'b11111111; //  660 : 255 - 0xff
      12'h295: dout  = 8'b11111111; //  661 : 255 - 0xff
      12'h296: dout  = 8'b11111011; //  662 : 251 - 0xfb
      12'h297: dout  = 8'b01110110; //  663 : 118 - 0x76
      12'h298: dout  = 8'b00100000; //  664 :  32 - 0x20 -- Sprite 0x53
      12'h299: dout  = 8'b11111000; //  665 : 248 - 0xf8
      12'h29A: dout  = 8'b11111111; //  666 : 255 - 0xff
      12'h29B: dout  = 8'b11000011; //  667 : 195 - 0xc3
      12'h29C: dout  = 8'b11111101; //  668 : 253 - 0xfd
      12'h29D: dout  = 8'b11111110; //  669 : 254 - 0xfe
      12'h29E: dout  = 8'b11110000; //  670 : 240 - 0xf0
      12'h29F: dout  = 8'b01000000; //  671 :  64 - 0x40
      12'h2A0: dout  = 8'b01000000; //  672 :  64 - 0x40 -- Sprite 0x54
      12'h2A1: dout  = 8'b11100000; //  673 : 224 - 0xe0
      12'h2A2: dout  = 8'b01000000; //  674 :  64 - 0x40
      12'h2A3: dout  = 8'b01000000; //  675 :  64 - 0x40
      12'h2A4: dout  = 8'b01000001; //  676 :  65 - 0x41
      12'h2A5: dout  = 8'b01000001; //  677 :  65 - 0x41
      12'h2A6: dout  = 8'b01001111; //  678 :  79 - 0x4f
      12'h2A7: dout  = 8'b01000111; //  679 :  71 - 0x47
      12'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout  = 8'b11100000; //  686 : 224 - 0xe0
      12'h2AF: dout  = 8'b11000000; //  687 : 192 - 0xc0
      12'h2B0: dout  = 8'b01000011; //  688 :  67 - 0x43 -- Sprite 0x56
      12'h2B1: dout  = 8'b01000110; //  689 :  70 - 0x46
      12'h2B2: dout  = 8'b01000100; //  690 :  68 - 0x44
      12'h2B3: dout  = 8'b01000000; //  691 :  64 - 0x40
      12'h2B4: dout  = 8'b01000000; //  692 :  64 - 0x40
      12'h2B5: dout  = 8'b01000000; //  693 :  64 - 0x40
      12'h2B6: dout  = 8'b01000000; //  694 :  64 - 0x40
      12'h2B7: dout  = 8'b01000000; //  695 :  64 - 0x40
      12'h2B8: dout  = 8'b10000000; //  696 : 128 - 0x80 -- Sprite 0x57
      12'h2B9: dout  = 8'b11000000; //  697 : 192 - 0xc0
      12'h2BA: dout  = 8'b01000000; //  698 :  64 - 0x40
      12'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b00110001; //  704 :  49 - 0x31 -- Sprite 0x58
      12'h2C1: dout  = 8'b00110000; //  705 :  48 - 0x30
      12'h2C2: dout  = 8'b00111000; //  706 :  56 - 0x38
      12'h2C3: dout  = 8'b01111100; //  707 : 124 - 0x7c
      12'h2C4: dout  = 8'b01111111; //  708 : 127 - 0x7f
      12'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      12'h2C6: dout  = 8'b11111111; //  710 : 255 - 0xff
      12'h2C7: dout  = 8'b11111011; //  711 : 251 - 0xfb
      12'h2C8: dout  = 8'b00010000; //  712 :  16 - 0x10 -- Sprite 0x59
      12'h2C9: dout  = 8'b01111110; //  713 : 126 - 0x7e
      12'h2CA: dout  = 8'b00111110; //  714 :  62 - 0x3e
      12'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout  = 8'b00011110; //  716 :  30 - 0x1e
      12'h2CD: dout  = 8'b11111110; //  717 : 254 - 0xfe
      12'h2CE: dout  = 8'b11111111; //  718 : 255 - 0xff
      12'h2CF: dout  = 8'b11111111; //  719 : 255 - 0xff
      12'h2D0: dout  = 8'b11111111; //  720 : 255 - 0xff -- Sprite 0x5a
      12'h2D1: dout  = 8'b11111111; //  721 : 255 - 0xff
      12'h2D2: dout  = 8'b11100011; //  722 : 227 - 0xe3
      12'h2D3: dout  = 8'b11000011; //  723 : 195 - 0xc3
      12'h2D4: dout  = 8'b10000111; //  724 : 135 - 0x87
      12'h2D5: dout  = 8'b01001000; //  725 :  72 - 0x48
      12'h2D6: dout  = 8'b00111100; //  726 :  60 - 0x3c
      12'h2D7: dout  = 8'b11111100; //  727 : 252 - 0xfc
      12'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout  = 8'b11111111; //  729 : 255 - 0xff
      12'h2DA: dout  = 8'b11000011; //  730 : 195 - 0xc3
      12'h2DB: dout  = 8'b10000011; //  731 : 131 - 0x83
      12'h2DC: dout  = 8'b10000011; //  732 : 131 - 0x83
      12'h2DD: dout  = 8'b11111111; //  733 : 255 - 0xff
      12'h2DE: dout  = 8'b11111111; //  734 : 255 - 0xff
      12'h2DF: dout  = 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout  = 8'b00011111; //  736 :  31 - 0x1f -- Sprite 0x5c
      12'h2E1: dout  = 8'b00011111; //  737 :  31 - 0x1f
      12'h2E2: dout  = 8'b00001111; //  738 :  15 - 0xf
      12'h2E3: dout  = 8'b00000111; //  739 :   7 - 0x7
      12'h2E4: dout  = 8'b00000001; //  740 :   1 - 0x1
      12'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b11110000; //  744 : 240 - 0xf0 -- Sprite 0x5d
      12'h2E9: dout  = 8'b11111011; //  745 : 251 - 0xfb
      12'h2EA: dout  = 8'b11111111; //  746 : 255 - 0xff
      12'h2EB: dout  = 8'b11111111; //  747 : 255 - 0xff
      12'h2EC: dout  = 8'b11111110; //  748 : 254 - 0xfe
      12'h2ED: dout  = 8'b00111110; //  749 :  62 - 0x3e
      12'h2EE: dout  = 8'b00001100; //  750 :  12 - 0xc
      12'h2EF: dout  = 8'b00000100; //  751 :   4 - 0x4
      12'h2F0: dout  = 8'b00011111; //  752 :  31 - 0x1f -- Sprite 0x5e
      12'h2F1: dout  = 8'b00011111; //  753 :  31 - 0x1f
      12'h2F2: dout  = 8'b00001111; //  754 :  15 - 0xf
      12'h2F3: dout  = 8'b00001111; //  755 :  15 - 0xf
      12'h2F4: dout  = 8'b00000111; //  756 :   7 - 0x7
      12'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout  = 8'b11111011; //  760 : 251 - 0xfb -- Sprite 0x5f
      12'h2F9: dout  = 8'b11111111; //  761 : 255 - 0xff
      12'h2FA: dout  = 8'b11111111; //  762 : 255 - 0xff
      12'h2FB: dout  = 8'b11111111; //  763 : 255 - 0xff
      12'h2FC: dout  = 8'b11111111; //  764 : 255 - 0xff
      12'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout  = 8'b00011000; //  769 :  24 - 0x18
      12'h302: dout  = 8'b00111100; //  770 :  60 - 0x3c
      12'h303: dout  = 8'b01111110; //  771 : 126 - 0x7e
      12'h304: dout  = 8'b01101110; //  772 : 110 - 0x6e
      12'h305: dout  = 8'b11011111; //  773 : 223 - 0xdf
      12'h306: dout  = 8'b11011111; //  774 : 223 - 0xdf
      12'h307: dout  = 8'b11011111; //  775 : 223 - 0xdf
      12'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      12'h309: dout  = 8'b00011000; //  777 :  24 - 0x18
      12'h30A: dout  = 8'b00011000; //  778 :  24 - 0x18
      12'h30B: dout  = 8'b00111100; //  779 :  60 - 0x3c
      12'h30C: dout  = 8'b00111100; //  780 :  60 - 0x3c
      12'h30D: dout  = 8'b00111100; //  781 :  60 - 0x3c
      12'h30E: dout  = 8'b00111100; //  782 :  60 - 0x3c
      12'h30F: dout  = 8'b00011100; //  783 :  28 - 0x1c
      12'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      12'h311: dout  = 8'b00001000; //  785 :   8 - 0x8
      12'h312: dout  = 8'b00001000; //  786 :   8 - 0x8
      12'h313: dout  = 8'b00001000; //  787 :   8 - 0x8
      12'h314: dout  = 8'b00001000; //  788 :   8 - 0x8
      12'h315: dout  = 8'b00001000; //  789 :   8 - 0x8
      12'h316: dout  = 8'b00001000; //  790 :   8 - 0x8
      12'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      12'h319: dout  = 8'b00001000; //  793 :   8 - 0x8
      12'h31A: dout  = 8'b00001000; //  794 :   8 - 0x8
      12'h31B: dout  = 8'b00000100; //  795 :   4 - 0x4
      12'h31C: dout  = 8'b00000100; //  796 :   4 - 0x4
      12'h31D: dout  = 8'b00000100; //  797 :   4 - 0x4
      12'h31E: dout  = 8'b00000100; //  798 :   4 - 0x4
      12'h31F: dout  = 8'b00000100; //  799 :   4 - 0x4
      12'h320: dout  = 8'b00111100; //  800 :  60 - 0x3c -- Sprite 0x64
      12'h321: dout  = 8'b01111110; //  801 : 126 - 0x7e
      12'h322: dout  = 8'b01110111; //  802 : 119 - 0x77
      12'h323: dout  = 8'b11111011; //  803 : 251 - 0xfb
      12'h324: dout  = 8'b10011111; //  804 : 159 - 0x9f
      12'h325: dout  = 8'b01011111; //  805 :  95 - 0x5f
      12'h326: dout  = 8'b10001110; //  806 : 142 - 0x8e
      12'h327: dout  = 8'b00100000; //  807 :  32 - 0x20
      12'h328: dout  = 8'b01011100; //  808 :  92 - 0x5c -- Sprite 0x65
      12'h329: dout  = 8'b00101110; //  809 :  46 - 0x2e
      12'h32A: dout  = 8'b10001111; //  810 : 143 - 0x8f
      12'h32B: dout  = 8'b00111111; //  811 :  63 - 0x3f
      12'h32C: dout  = 8'b01111011; //  812 : 123 - 0x7b
      12'h32D: dout  = 8'b01110111; //  813 : 119 - 0x77
      12'h32E: dout  = 8'b01111110; //  814 : 126 - 0x7e
      12'h32F: dout  = 8'b00111100; //  815 :  60 - 0x3c
      12'h330: dout  = 8'b00010011; //  816 :  19 - 0x13 -- Sprite 0x66
      12'h331: dout  = 8'b01001111; //  817 :  79 - 0x4f
      12'h332: dout  = 8'b00111111; //  818 :  63 - 0x3f
      12'h333: dout  = 8'b10111111; //  819 : 191 - 0xbf
      12'h334: dout  = 8'b00111111; //  820 :  63 - 0x3f
      12'h335: dout  = 8'b01111010; //  821 : 122 - 0x7a
      12'h336: dout  = 8'b11111000; //  822 : 248 - 0xf8
      12'h337: dout  = 8'b11111000; //  823 : 248 - 0xf8
      12'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      12'h339: dout  = 8'b00001000; //  825 :   8 - 0x8
      12'h33A: dout  = 8'b00000101; //  826 :   5 - 0x5
      12'h33B: dout  = 8'b00001111; //  827 :  15 - 0xf
      12'h33C: dout  = 8'b00101111; //  828 :  47 - 0x2f
      12'h33D: dout  = 8'b00011101; //  829 :  29 - 0x1d
      12'h33E: dout  = 8'b00011100; //  830 :  28 - 0x1c
      12'h33F: dout  = 8'b00111100; //  831 :  60 - 0x3c
      12'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout  = 8'b00000010; //  836 :   2 - 0x2
      12'h345: dout  = 8'b00001011; //  837 :  11 - 0xb
      12'h346: dout  = 8'b00000111; //  838 :   7 - 0x7
      12'h347: dout  = 8'b00001111; //  839 :  15 - 0xf
      12'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout  = 8'b00001000; //  845 :   8 - 0x8
      12'h34E: dout  = 8'b00000100; //  846 :   4 - 0x4
      12'h34F: dout  = 8'b00000100; //  847 :   4 - 0x4
      12'h350: dout  = 8'b00000010; //  848 :   2 - 0x2 -- Sprite 0x6a
      12'h351: dout  = 8'b00000010; //  849 :   2 - 0x2
      12'h352: dout  = 8'b00000010; //  850 :   2 - 0x2
      12'h353: dout  = 8'b00000101; //  851 :   5 - 0x5
      12'h354: dout  = 8'b01110001; //  852 : 113 - 0x71
      12'h355: dout  = 8'b01111111; //  853 : 127 - 0x7f
      12'h356: dout  = 8'b01111111; //  854 : 127 - 0x7f
      12'h357: dout  = 8'b01111111; //  855 : 127 - 0x7f
      12'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout  = 8'b00000100; //  863 :   4 - 0x4
      12'h360: dout  = 8'b00000010; //  864 :   2 - 0x2 -- Sprite 0x6c
      12'h361: dout  = 8'b00000010; //  865 :   2 - 0x2
      12'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout  = 8'b00000001; //  867 :   1 - 0x1
      12'h364: dout  = 8'b00010011; //  868 :  19 - 0x13
      12'h365: dout  = 8'b00111111; //  869 :  63 - 0x3f
      12'h366: dout  = 8'b01111111; //  870 : 127 - 0x7f
      12'h367: dout  = 8'b01111111; //  871 : 127 - 0x7f
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout  = 8'b01000000; //  873 :  64 - 0x40
      12'h36A: dout  = 8'b01100000; //  874 :  96 - 0x60
      12'h36B: dout  = 8'b01110000; //  875 : 112 - 0x70
      12'h36C: dout  = 8'b01110011; //  876 : 115 - 0x73
      12'h36D: dout  = 8'b00100111; //  877 :  39 - 0x27
      12'h36E: dout  = 8'b00001111; //  878 :  15 - 0xf
      12'h36F: dout  = 8'b00011111; //  879 :  31 - 0x1f
      12'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout  = 8'b00000011; //  884 :   3 - 0x3
      12'h375: dout  = 8'b00000111; //  885 :   7 - 0x7
      12'h376: dout  = 8'b00001111; //  886 :  15 - 0xf
      12'h377: dout  = 8'b00011111; //  887 :  31 - 0x1f
      12'h378: dout  = 8'b01111111; //  888 : 127 - 0x7f -- Sprite 0x6f
      12'h379: dout  = 8'b01111111; //  889 : 127 - 0x7f
      12'h37A: dout  = 8'b00111111; //  890 :  63 - 0x3f
      12'h37B: dout  = 8'b00111111; //  891 :  63 - 0x3f
      12'h37C: dout  = 8'b00011111; //  892 :  31 - 0x1f
      12'h37D: dout  = 8'b00011111; //  893 :  31 - 0x1f
      12'h37E: dout  = 8'b00001111; //  894 :  15 - 0xf
      12'h37F: dout  = 8'b00000111; //  895 :   7 - 0x7
      12'h380: dout  = 8'b00000011; //  896 :   3 - 0x3 -- Sprite 0x70
      12'h381: dout  = 8'b00000111; //  897 :   7 - 0x7
      12'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      12'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      12'h384: dout  = 8'b00111111; //  900 :  63 - 0x3f
      12'h385: dout  = 8'b01110111; //  901 : 119 - 0x77
      12'h386: dout  = 8'b01110111; //  902 : 119 - 0x77
      12'h387: dout  = 8'b11110101; //  903 : 245 - 0xf5
      12'h388: dout  = 8'b11000000; //  904 : 192 - 0xc0 -- Sprite 0x71
      12'h389: dout  = 8'b11100000; //  905 : 224 - 0xe0
      12'h38A: dout  = 8'b11110000; //  906 : 240 - 0xf0
      12'h38B: dout  = 8'b11111000; //  907 : 248 - 0xf8
      12'h38C: dout  = 8'b11111100; //  908 : 252 - 0xfc
      12'h38D: dout  = 8'b11101110; //  909 : 238 - 0xee
      12'h38E: dout  = 8'b11101110; //  910 : 238 - 0xee
      12'h38F: dout  = 8'b10101111; //  911 : 175 - 0xaf
      12'h390: dout  = 8'b11110001; //  912 : 241 - 0xf1 -- Sprite 0x72
      12'h391: dout  = 8'b11111111; //  913 : 255 - 0xff
      12'h392: dout  = 8'b01111000; //  914 : 120 - 0x78
      12'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout  = 8'b00011000; //  917 :  24 - 0x18
      12'h396: dout  = 8'b00011100; //  918 :  28 - 0x1c
      12'h397: dout  = 8'b00001110; //  919 :  14 - 0xe
      12'h398: dout  = 8'b10001111; //  920 : 143 - 0x8f -- Sprite 0x73
      12'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout  = 8'b00011110; //  922 :  30 - 0x1e
      12'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout  = 8'b00001100; //  924 :  12 - 0xc
      12'h39D: dout  = 8'b00111110; //  925 :  62 - 0x3e
      12'h39E: dout  = 8'b01111110; //  926 : 126 - 0x7e
      12'h39F: dout  = 8'b01111100; //  927 : 124 - 0x7c
      12'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      12'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      12'h3A9: dout  = 8'b00000010; //  937 :   2 - 0x2
      12'h3AA: dout  = 8'b01000001; //  938 :  65 - 0x41
      12'h3AB: dout  = 8'b01000001; //  939 :  65 - 0x41
      12'h3AC: dout  = 8'b01100001; //  940 :  97 - 0x61
      12'h3AD: dout  = 8'b00110011; //  941 :  51 - 0x33
      12'h3AE: dout  = 8'b00000110; //  942 :   6 - 0x6
      12'h3AF: dout  = 8'b00111100; //  943 :  60 - 0x3c
      12'h3B0: dout  = 8'b00000011; //  944 :   3 - 0x3 -- Sprite 0x76
      12'h3B1: dout  = 8'b00000111; //  945 :   7 - 0x7
      12'h3B2: dout  = 8'b00001111; //  946 :  15 - 0xf
      12'h3B3: dout  = 8'b00011111; //  947 :  31 - 0x1f
      12'h3B4: dout  = 8'b00111111; //  948 :  63 - 0x3f
      12'h3B5: dout  = 8'b01111111; //  949 : 127 - 0x7f
      12'h3B6: dout  = 8'b01111111; //  950 : 127 - 0x7f
      12'h3B7: dout  = 8'b11111111; //  951 : 255 - 0xff
      12'h3B8: dout  = 8'b11000000; //  952 : 192 - 0xc0 -- Sprite 0x77
      12'h3B9: dout  = 8'b11100000; //  953 : 224 - 0xe0
      12'h3BA: dout  = 8'b11110000; //  954 : 240 - 0xf0
      12'h3BB: dout  = 8'b11111000; //  955 : 248 - 0xf8
      12'h3BC: dout  = 8'b11111100; //  956 : 252 - 0xfc
      12'h3BD: dout  = 8'b11111110; //  957 : 254 - 0xfe
      12'h3BE: dout  = 8'b11111110; //  958 : 254 - 0xfe
      12'h3BF: dout  = 8'b11111111; //  959 : 255 - 0xff
      12'h3C0: dout  = 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      12'h3C1: dout  = 8'b11111111; //  961 : 255 - 0xff
      12'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout  = 8'b01111000; //  963 : 120 - 0x78
      12'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      12'h3C9: dout  = 8'b11111111; //  969 : 255 - 0xff
      12'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      12'h3CB: dout  = 8'b00011110; //  971 :  30 - 0x1e
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b00100000; //  973 :  32 - 0x20
      12'h3CE: dout  = 8'b00100000; //  974 :  32 - 0x20
      12'h3CF: dout  = 8'b01000000; //  975 :  64 - 0x40
      12'h3D0: dout  = 8'b00010110; //  976 :  22 - 0x16 -- Sprite 0x7a
      12'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      12'h3D2: dout  = 8'b00111111; //  978 :  63 - 0x3f
      12'h3D3: dout  = 8'b01111111; //  979 : 127 - 0x7f
      12'h3D4: dout  = 8'b00111101; //  980 :  61 - 0x3d
      12'h3D5: dout  = 8'b00011101; //  981 :  29 - 0x1d
      12'h3D6: dout  = 8'b00111111; //  982 :  63 - 0x3f
      12'h3D7: dout  = 8'b00011111; //  983 :  31 - 0x1f
      12'h3D8: dout  = 8'b10000000; //  984 : 128 - 0x80 -- Sprite 0x7b
      12'h3D9: dout  = 8'b10000000; //  985 : 128 - 0x80
      12'h3DA: dout  = 8'b11000000; //  986 : 192 - 0xc0
      12'h3DB: dout  = 8'b11100000; //  987 : 224 - 0xe0
      12'h3DC: dout  = 8'b11110000; //  988 : 240 - 0xf0
      12'h3DD: dout  = 8'b11110000; //  989 : 240 - 0xf0
      12'h3DE: dout  = 8'b11110000; //  990 : 240 - 0xf0
      12'h3DF: dout  = 8'b11111000; //  991 : 248 - 0xf8
      12'h3E0: dout  = 8'b00111100; //  992 :  60 - 0x3c -- Sprite 0x7c
      12'h3E1: dout  = 8'b11111010; //  993 : 250 - 0xfa
      12'h3E2: dout  = 8'b10110001; //  994 : 177 - 0xb1
      12'h3E3: dout  = 8'b01110010; //  995 : 114 - 0x72
      12'h3E4: dout  = 8'b11110010; //  996 : 242 - 0xf2
      12'h3E5: dout  = 8'b11011011; //  997 : 219 - 0xdb
      12'h3E6: dout  = 8'b11011111; //  998 : 223 - 0xdf
      12'h3E7: dout  = 8'b01011111; //  999 :  95 - 0x5f
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000001; // 1003 :   1 - 0x1
      12'h3EC: dout  = 8'b00000001; // 1004 :   1 - 0x1
      12'h3ED: dout  = 8'b00000001; // 1005 :   1 - 0x1
      12'h3EE: dout  = 8'b00000110; // 1006 :   6 - 0x6
      12'h3EF: dout  = 8'b00011110; // 1007 :  30 - 0x1e
      12'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      12'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      12'h3F9: dout  = 8'b01111100; // 1017 : 124 - 0x7c
      12'h3FA: dout  = 8'b11010110; // 1018 : 214 - 0xd6
      12'h3FB: dout  = 8'b10010010; // 1019 : 146 - 0x92
      12'h3FC: dout  = 8'b10111010; // 1020 : 186 - 0xba
      12'h3FD: dout  = 8'b11101110; // 1021 : 238 - 0xee
      12'h3FE: dout  = 8'b11111110; // 1022 : 254 - 0xfe
      12'h3FF: dout  = 8'b00111000; // 1023 :  56 - 0x38
      12'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      12'h401: dout  = 8'b00010101; // 1025 :  21 - 0x15
      12'h402: dout  = 8'b00111111; // 1026 :  63 - 0x3f
      12'h403: dout  = 8'b01100010; // 1027 :  98 - 0x62
      12'h404: dout  = 8'b01011111; // 1028 :  95 - 0x5f
      12'h405: dout  = 8'b11111111; // 1029 : 255 - 0xff
      12'h406: dout  = 8'b10011111; // 1030 : 159 - 0x9f
      12'h407: dout  = 8'b01111101; // 1031 : 125 - 0x7d
      12'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      12'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout  = 8'b00101111; // 1040 :  47 - 0x2f -- Sprite 0x82
      12'h411: dout  = 8'b00011110; // 1041 :  30 - 0x1e
      12'h412: dout  = 8'b00101111; // 1042 :  47 - 0x2f
      12'h413: dout  = 8'b00101111; // 1043 :  47 - 0x2f
      12'h414: dout  = 8'b00101111; // 1044 :  47 - 0x2f
      12'h415: dout  = 8'b00010101; // 1045 :  21 - 0x15
      12'h416: dout  = 8'b00001101; // 1046 :  13 - 0xd
      12'h417: dout  = 8'b00001110; // 1047 :  14 - 0xe
      12'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      12'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout  = 8'b00011100; // 1056 :  28 - 0x1c -- Sprite 0x84
      12'h421: dout  = 8'b00111110; // 1057 :  62 - 0x3e
      12'h422: dout  = 8'b01111111; // 1058 : 127 - 0x7f
      12'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      12'h424: dout  = 8'b11111111; // 1060 : 255 - 0xff
      12'h425: dout  = 8'b11111110; // 1061 : 254 - 0xfe
      12'h426: dout  = 8'b01111100; // 1062 : 124 - 0x7c
      12'h427: dout  = 8'b00111000; // 1063 :  56 - 0x38
      12'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- Sprite 0x85
      12'h429: dout  = 8'b11111111; // 1065 : 255 - 0xff
      12'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout  = 8'b11111111; // 1067 : 255 - 0xff
      12'h42C: dout  = 8'b11111111; // 1068 : 255 - 0xff
      12'h42D: dout  = 8'b11111111; // 1069 : 255 - 0xff
      12'h42E: dout  = 8'b11111111; // 1070 : 255 - 0xff
      12'h42F: dout  = 8'b11111111; // 1071 : 255 - 0xff
      12'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      12'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      12'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      12'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      12'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      12'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      12'h436: dout  = 8'b11111111; // 1078 : 255 - 0xff
      12'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      12'h438: dout  = 8'b01111111; // 1080 : 127 - 0x7f -- Sprite 0x87
      12'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      12'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      12'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      12'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      12'h43D: dout  = 8'b11111111; // 1085 : 255 - 0xff
      12'h43E: dout  = 8'b11111111; // 1086 : 255 - 0xff
      12'h43F: dout  = 8'b11111111; // 1087 : 255 - 0xff
      12'h440: dout  = 8'b01101000; // 1088 : 104 - 0x68 -- Sprite 0x88
      12'h441: dout  = 8'b01001110; // 1089 :  78 - 0x4e
      12'h442: dout  = 8'b11100000; // 1090 : 224 - 0xe0
      12'h443: dout  = 8'b11100000; // 1091 : 224 - 0xe0
      12'h444: dout  = 8'b11100000; // 1092 : 224 - 0xe0
      12'h445: dout  = 8'b11110000; // 1093 : 240 - 0xf0
      12'h446: dout  = 8'b11111000; // 1094 : 248 - 0xf8
      12'h447: dout  = 8'b11111100; // 1095 : 252 - 0xfc
      12'h448: dout  = 8'b00111111; // 1096 :  63 - 0x3f -- Sprite 0x89
      12'h449: dout  = 8'b01011100; // 1097 :  92 - 0x5c
      12'h44A: dout  = 8'b00111001; // 1098 :  57 - 0x39
      12'h44B: dout  = 8'b00111011; // 1099 :  59 - 0x3b
      12'h44C: dout  = 8'b10111011; // 1100 : 187 - 0xbb
      12'h44D: dout  = 8'b11111001; // 1101 : 249 - 0xf9
      12'h44E: dout  = 8'b11111100; // 1102 : 252 - 0xfc
      12'h44F: dout  = 8'b11111110; // 1103 : 254 - 0xfe
      12'h450: dout  = 8'b11000000; // 1104 : 192 - 0xc0 -- Sprite 0x8a
      12'h451: dout  = 8'b11110000; // 1105 : 240 - 0xf0
      12'h452: dout  = 8'b11110000; // 1106 : 240 - 0xf0
      12'h453: dout  = 8'b11110000; // 1107 : 240 - 0xf0
      12'h454: dout  = 8'b11110000; // 1108 : 240 - 0xf0
      12'h455: dout  = 8'b11100000; // 1109 : 224 - 0xe0
      12'h456: dout  = 8'b11000000; // 1110 : 192 - 0xc0
      12'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe -- Sprite 0x8b
      12'h459: dout  = 8'b11111100; // 1113 : 252 - 0xfc
      12'h45A: dout  = 8'b01100001; // 1114 :  97 - 0x61
      12'h45B: dout  = 8'b00001111; // 1115 :  15 - 0xf
      12'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      12'h45D: dout  = 8'b11111110; // 1117 : 254 - 0xfe
      12'h45E: dout  = 8'b11110000; // 1118 : 240 - 0xf0
      12'h45F: dout  = 8'b11100000; // 1119 : 224 - 0xe0
      12'h460: dout  = 8'b01101110; // 1120 : 110 - 0x6e -- Sprite 0x8c
      12'h461: dout  = 8'b01000000; // 1121 :  64 - 0x40
      12'h462: dout  = 8'b11100000; // 1122 : 224 - 0xe0
      12'h463: dout  = 8'b11100000; // 1123 : 224 - 0xe0
      12'h464: dout  = 8'b11100000; // 1124 : 224 - 0xe0
      12'h465: dout  = 8'b11100000; // 1125 : 224 - 0xe0
      12'h466: dout  = 8'b11100000; // 1126 : 224 - 0xe0
      12'h467: dout  = 8'b11000000; // 1127 : 192 - 0xc0
      12'h468: dout  = 8'b00000001; // 1128 :   1 - 0x1 -- Sprite 0x8d
      12'h469: dout  = 8'b00000001; // 1129 :   1 - 0x1
      12'h46A: dout  = 8'b00000011; // 1130 :   3 - 0x3
      12'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      12'h46C: dout  = 8'b00000111; // 1132 :   7 - 0x7
      12'h46D: dout  = 8'b01111111; // 1133 : 127 - 0x7f
      12'h46E: dout  = 8'b01111111; // 1134 : 127 - 0x7f
      12'h46F: dout  = 8'b00111111; // 1135 :  63 - 0x3f
      12'h470: dout  = 8'b00000110; // 1136 :   6 - 0x6 -- Sprite 0x8e
      12'h471: dout  = 8'b00000111; // 1137 :   7 - 0x7
      12'h472: dout  = 8'b00111111; // 1138 :  63 - 0x3f
      12'h473: dout  = 8'b00111100; // 1139 :  60 - 0x3c
      12'h474: dout  = 8'b00011001; // 1140 :  25 - 0x19
      12'h475: dout  = 8'b01111011; // 1141 : 123 - 0x7b
      12'h476: dout  = 8'b01111111; // 1142 : 127 - 0x7f
      12'h477: dout  = 8'b00111111; // 1143 :  63 - 0x3f
      12'h478: dout  = 8'b00111111; // 1144 :  63 - 0x3f -- Sprite 0x8f
      12'h479: dout  = 8'b01111111; // 1145 : 127 - 0x7f
      12'h47A: dout  = 8'b01111111; // 1146 : 127 - 0x7f
      12'h47B: dout  = 8'b00011111; // 1147 :  31 - 0x1f
      12'h47C: dout  = 8'b00111111; // 1148 :  63 - 0x3f
      12'h47D: dout  = 8'b00111111; // 1149 :  63 - 0x3f
      12'h47E: dout  = 8'b00000111; // 1150 :   7 - 0x7
      12'h47F: dout  = 8'b00000110; // 1151 :   6 - 0x6
      12'h480: dout  = 8'b00000011; // 1152 :   3 - 0x3 -- Sprite 0x90
      12'h481: dout  = 8'b00000111; // 1153 :   7 - 0x7
      12'h482: dout  = 8'b00001111; // 1154 :  15 - 0xf
      12'h483: dout  = 8'b00001111; // 1155 :  15 - 0xf
      12'h484: dout  = 8'b00001111; // 1156 :  15 - 0xf
      12'h485: dout  = 8'b00001111; // 1157 :  15 - 0xf
      12'h486: dout  = 8'b00000111; // 1158 :   7 - 0x7
      12'h487: dout  = 8'b00000011; // 1159 :   3 - 0x3
      12'h488: dout  = 8'b11111000; // 1160 : 248 - 0xf8 -- Sprite 0x91
      12'h489: dout  = 8'b11111000; // 1161 : 248 - 0xf8
      12'h48A: dout  = 8'b11111000; // 1162 : 248 - 0xf8
      12'h48B: dout  = 8'b10100000; // 1163 : 160 - 0xa0
      12'h48C: dout  = 8'b11100001; // 1164 : 225 - 0xe1
      12'h48D: dout  = 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout  = 8'b11111111; // 1166 : 255 - 0xff
      12'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      12'h490: dout  = 8'b00001111; // 1168 :  15 - 0xf -- Sprite 0x92
      12'h491: dout  = 8'b00001111; // 1169 :  15 - 0xf
      12'h492: dout  = 8'b00001111; // 1170 :  15 - 0xf
      12'h493: dout  = 8'b00011111; // 1171 :  31 - 0x1f
      12'h494: dout  = 8'b00011111; // 1172 :  31 - 0x1f
      12'h495: dout  = 8'b00011111; // 1173 :  31 - 0x1f
      12'h496: dout  = 8'b00001111; // 1174 :  15 - 0xf
      12'h497: dout  = 8'b00000111; // 1175 :   7 - 0x7
      12'h498: dout  = 8'b11100000; // 1176 : 224 - 0xe0 -- Sprite 0x93
      12'h499: dout  = 8'b11111000; // 1177 : 248 - 0xf8
      12'h49A: dout  = 8'b11111000; // 1178 : 248 - 0xf8
      12'h49B: dout  = 8'b11111000; // 1179 : 248 - 0xf8
      12'h49C: dout  = 8'b11111111; // 1180 : 255 - 0xff
      12'h49D: dout  = 8'b11111110; // 1181 : 254 - 0xfe
      12'h49E: dout  = 8'b11110000; // 1182 : 240 - 0xf0
      12'h49F: dout  = 8'b11000000; // 1183 : 192 - 0xc0
      12'h4A0: dout  = 8'b00000001; // 1184 :   1 - 0x1 -- Sprite 0x94
      12'h4A1: dout  = 8'b00001111; // 1185 :  15 - 0xf
      12'h4A2: dout  = 8'b00001111; // 1186 :  15 - 0xf
      12'h4A3: dout  = 8'b00011111; // 1187 :  31 - 0x1f
      12'h4A4: dout  = 8'b00111001; // 1188 :  57 - 0x39
      12'h4A5: dout  = 8'b00110011; // 1189 :  51 - 0x33
      12'h4A6: dout  = 8'b00110111; // 1190 :  55 - 0x37
      12'h4A7: dout  = 8'b01111111; // 1191 : 127 - 0x7f
      12'h4A8: dout  = 8'b01111111; // 1192 : 127 - 0x7f -- Sprite 0x95
      12'h4A9: dout  = 8'b00111111; // 1193 :  63 - 0x3f
      12'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      12'h4AB: dout  = 8'b00111111; // 1195 :  63 - 0x3f
      12'h4AC: dout  = 8'b00011111; // 1196 :  31 - 0x1f
      12'h4AD: dout  = 8'b00001111; // 1197 :  15 - 0xf
      12'h4AE: dout  = 8'b00001111; // 1198 :  15 - 0xf
      12'h4AF: dout  = 8'b00000001; // 1199 :   1 - 0x1
      12'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      12'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout  = 8'b00000011; // 1202 :   3 - 0x3
      12'h4B3: dout  = 8'b00000011; // 1203 :   3 - 0x3
      12'h4B4: dout  = 8'b01000111; // 1204 :  71 - 0x47
      12'h4B5: dout  = 8'b01100111; // 1205 : 103 - 0x67
      12'h4B6: dout  = 8'b01110111; // 1206 : 119 - 0x77
      12'h4B7: dout  = 8'b01110111; // 1207 : 119 - 0x77
      12'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- Sprite 0x97
      12'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout  = 8'b10001000; // 1212 : 136 - 0x88
      12'h4BD: dout  = 8'b10011000; // 1213 : 152 - 0x98
      12'h4BE: dout  = 8'b11111000; // 1214 : 248 - 0xf8
      12'h4BF: dout  = 8'b11110000; // 1215 : 240 - 0xf0
      12'h4C0: dout  = 8'b01111110; // 1216 : 126 - 0x7e -- Sprite 0x98
      12'h4C1: dout  = 8'b01111111; // 1217 : 127 - 0x7f
      12'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout  = 8'b00011111; // 1219 :  31 - 0x1f
      12'h4C4: dout  = 8'b00000111; // 1220 :   7 - 0x7
      12'h4C5: dout  = 8'b00110000; // 1221 :  48 - 0x30
      12'h4C6: dout  = 8'b00011100; // 1222 :  28 - 0x1c
      12'h4C7: dout  = 8'b00001100; // 1223 :  12 - 0xc
      12'h4C8: dout  = 8'b01111110; // 1224 : 126 - 0x7e -- Sprite 0x99
      12'h4C9: dout  = 8'b00111000; // 1225 :  56 - 0x38
      12'h4CA: dout  = 8'b11110110; // 1226 : 246 - 0xf6
      12'h4CB: dout  = 8'b11101101; // 1227 : 237 - 0xed
      12'h4CC: dout  = 8'b11011111; // 1228 : 223 - 0xdf
      12'h4CD: dout  = 8'b00111000; // 1229 :  56 - 0x38
      12'h4CE: dout  = 8'b01110000; // 1230 : 112 - 0x70
      12'h4CF: dout  = 8'b01100000; // 1231 :  96 - 0x60
      12'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      12'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout  = 8'b00000011; // 1235 :   3 - 0x3
      12'h4D4: dout  = 8'b00000011; // 1236 :   3 - 0x3
      12'h4D5: dout  = 8'b01000111; // 1237 :  71 - 0x47
      12'h4D6: dout  = 8'b01100111; // 1238 : 103 - 0x67
      12'h4D7: dout  = 8'b01110111; // 1239 : 119 - 0x77
      12'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- Sprite 0x9b
      12'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout  = 8'b10001000; // 1245 : 136 - 0x88
      12'h4DE: dout  = 8'b10011000; // 1246 : 152 - 0x98
      12'h4DF: dout  = 8'b11111000; // 1247 : 248 - 0xf8
      12'h4E0: dout  = 8'b01110111; // 1248 : 119 - 0x77 -- Sprite 0x9c
      12'h4E1: dout  = 8'b01111110; // 1249 : 126 - 0x7e
      12'h4E2: dout  = 8'b01111111; // 1250 : 127 - 0x7f
      12'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      12'h4E4: dout  = 8'b00011111; // 1252 :  31 - 0x1f
      12'h4E5: dout  = 8'b00000111; // 1253 :   7 - 0x7
      12'h4E6: dout  = 8'b01110000; // 1254 : 112 - 0x70
      12'h4E7: dout  = 8'b11110000; // 1255 : 240 - 0xf0
      12'h4E8: dout  = 8'b11110000; // 1256 : 240 - 0xf0 -- Sprite 0x9d
      12'h4E9: dout  = 8'b01111110; // 1257 : 126 - 0x7e
      12'h4EA: dout  = 8'b00111000; // 1258 :  56 - 0x38
      12'h4EB: dout  = 8'b11110110; // 1259 : 246 - 0xf6
      12'h4EC: dout  = 8'b11101101; // 1260 : 237 - 0xed
      12'h4ED: dout  = 8'b11011111; // 1261 : 223 - 0xdf
      12'h4EE: dout  = 8'b00111000; // 1262 :  56 - 0x38
      12'h4EF: dout  = 8'b00111100; // 1263 :  60 - 0x3c
      12'h4F0: dout  = 8'b00000011; // 1264 :   3 - 0x3 -- Sprite 0x9e
      12'h4F1: dout  = 8'b00000111; // 1265 :   7 - 0x7
      12'h4F2: dout  = 8'b00001010; // 1266 :  10 - 0xa
      12'h4F3: dout  = 8'b00011010; // 1267 :  26 - 0x1a
      12'h4F4: dout  = 8'b00011100; // 1268 :  28 - 0x1c
      12'h4F5: dout  = 8'b00011110; // 1269 :  30 - 0x1e
      12'h4F6: dout  = 8'b00001011; // 1270 :  11 - 0xb
      12'h4F7: dout  = 8'b00001000; // 1271 :   8 - 0x8
      12'h4F8: dout  = 8'b00011100; // 1272 :  28 - 0x1c -- Sprite 0x9f
      12'h4F9: dout  = 8'b00111111; // 1273 :  63 - 0x3f
      12'h4FA: dout  = 8'b00111111; // 1274 :  63 - 0x3f
      12'h4FB: dout  = 8'b00111101; // 1275 :  61 - 0x3d
      12'h4FC: dout  = 8'b00111111; // 1276 :  63 - 0x3f
      12'h4FD: dout  = 8'b00011111; // 1277 :  31 - 0x1f
      12'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      12'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout  = 8'b00000100; // 1282 :   4 - 0x4
      12'h503: dout  = 8'b01001100; // 1283 :  76 - 0x4c
      12'h504: dout  = 8'b01001110; // 1284 :  78 - 0x4e
      12'h505: dout  = 8'b01001110; // 1285 :  78 - 0x4e
      12'h506: dout  = 8'b01000110; // 1286 :  70 - 0x46
      12'h507: dout  = 8'b01101111; // 1287 : 111 - 0x6f
      12'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      12'h509: dout  = 8'b00011111; // 1289 :  31 - 0x1f
      12'h50A: dout  = 8'b00111111; // 1290 :  63 - 0x3f
      12'h50B: dout  = 8'b00111111; // 1291 :  63 - 0x3f
      12'h50C: dout  = 8'b01001111; // 1292 :  79 - 0x4f
      12'h50D: dout  = 8'b01011111; // 1293 :  95 - 0x5f
      12'h50E: dout  = 8'b01111111; // 1294 : 127 - 0x7f
      12'h50F: dout  = 8'b01111111; // 1295 : 127 - 0x7f
      12'h510: dout  = 8'b01111111; // 1296 : 127 - 0x7f -- Sprite 0xa2
      12'h511: dout  = 8'b01100111; // 1297 : 103 - 0x67
      12'h512: dout  = 8'b10100011; // 1298 : 163 - 0xa3
      12'h513: dout  = 8'b10110000; // 1299 : 176 - 0xb0
      12'h514: dout  = 8'b11011000; // 1300 : 216 - 0xd8
      12'h515: dout  = 8'b11011110; // 1301 : 222 - 0xde
      12'h516: dout  = 8'b11011100; // 1302 : 220 - 0xdc
      12'h517: dout  = 8'b11001000; // 1303 : 200 - 0xc8
      12'h518: dout  = 8'b01111111; // 1304 : 127 - 0x7f -- Sprite 0xa3
      12'h519: dout  = 8'b01111111; // 1305 : 127 - 0x7f
      12'h51A: dout  = 8'b01111111; // 1306 : 127 - 0x7f
      12'h51B: dout  = 8'b00011111; // 1307 :  31 - 0x1f
      12'h51C: dout  = 8'b01000111; // 1308 :  71 - 0x47
      12'h51D: dout  = 8'b01110000; // 1309 : 112 - 0x70
      12'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      12'h51F: dout  = 8'b00111001; // 1311 :  57 - 0x39
      12'h520: dout  = 8'b11101000; // 1312 : 232 - 0xe8 -- Sprite 0xa4
      12'h521: dout  = 8'b11101000; // 1313 : 232 - 0xe8
      12'h522: dout  = 8'b11100000; // 1314 : 224 - 0xe0
      12'h523: dout  = 8'b11000000; // 1315 : 192 - 0xc0
      12'h524: dout  = 8'b00010000; // 1316 :  16 - 0x10
      12'h525: dout  = 8'b01110000; // 1317 : 112 - 0x70
      12'h526: dout  = 8'b11100000; // 1318 : 224 - 0xe0
      12'h527: dout  = 8'b11000000; // 1319 : 192 - 0xc0
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      12'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout  = 8'b00100000; // 1323 :  32 - 0x20
      12'h52C: dout  = 8'b01100110; // 1324 : 102 - 0x66
      12'h52D: dout  = 8'b01100110; // 1325 : 102 - 0x66
      12'h52E: dout  = 8'b01100110; // 1326 : 102 - 0x66
      12'h52F: dout  = 8'b01100010; // 1327 :  98 - 0x62
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout  = 8'b00011111; // 1330 :  31 - 0x1f
      12'h533: dout  = 8'b00111111; // 1331 :  63 - 0x3f
      12'h534: dout  = 8'b01111111; // 1332 : 127 - 0x7f
      12'h535: dout  = 8'b01001111; // 1333 :  79 - 0x4f
      12'h536: dout  = 8'b01011111; // 1334 :  95 - 0x5f
      12'h537: dout  = 8'b01111111; // 1335 : 127 - 0x7f
      12'h538: dout  = 8'b01110111; // 1336 : 119 - 0x77 -- Sprite 0xa7
      12'h539: dout  = 8'b01111111; // 1337 : 127 - 0x7f
      12'h53A: dout  = 8'b00111111; // 1338 :  63 - 0x3f
      12'h53B: dout  = 8'b10110111; // 1339 : 183 - 0xb7
      12'h53C: dout  = 8'b10110011; // 1340 : 179 - 0xb3
      12'h53D: dout  = 8'b11011011; // 1341 : 219 - 0xdb
      12'h53E: dout  = 8'b11011010; // 1342 : 218 - 0xda
      12'h53F: dout  = 8'b11011000; // 1343 : 216 - 0xd8
      12'h540: dout  = 8'b01111111; // 1344 : 127 - 0x7f -- Sprite 0xa8
      12'h541: dout  = 8'b01111111; // 1345 : 127 - 0x7f
      12'h542: dout  = 8'b01111111; // 1346 : 127 - 0x7f
      12'h543: dout  = 8'b01111111; // 1347 : 127 - 0x7f
      12'h544: dout  = 8'b00011111; // 1348 :  31 - 0x1f
      12'h545: dout  = 8'b00000111; // 1349 :   7 - 0x7
      12'h546: dout  = 8'b01110000; // 1350 : 112 - 0x70
      12'h547: dout  = 8'b11110000; // 1351 : 240 - 0xf0
      12'h548: dout  = 8'b11001100; // 1352 : 204 - 0xcc -- Sprite 0xa9
      12'h549: dout  = 8'b11101000; // 1353 : 232 - 0xe8
      12'h54A: dout  = 8'b11101000; // 1354 : 232 - 0xe8
      12'h54B: dout  = 8'b11100000; // 1355 : 224 - 0xe0
      12'h54C: dout  = 8'b11000000; // 1356 : 192 - 0xc0
      12'h54D: dout  = 8'b00011000; // 1357 :  24 - 0x18
      12'h54E: dout  = 8'b01111100; // 1358 : 124 - 0x7c
      12'h54F: dout  = 8'b00111110; // 1359 :  62 - 0x3e
      12'h550: dout  = 8'b00000011; // 1360 :   3 - 0x3 -- Sprite 0xaa
      12'h551: dout  = 8'b00001111; // 1361 :  15 - 0xf
      12'h552: dout  = 8'b00011111; // 1362 :  31 - 0x1f
      12'h553: dout  = 8'b00111111; // 1363 :  63 - 0x3f
      12'h554: dout  = 8'b00111011; // 1364 :  59 - 0x3b
      12'h555: dout  = 8'b00111111; // 1365 :  63 - 0x3f
      12'h556: dout  = 8'b01111111; // 1366 : 127 - 0x7f
      12'h557: dout  = 8'b01111111; // 1367 : 127 - 0x7f
      12'h558: dout  = 8'b10000000; // 1368 : 128 - 0x80 -- Sprite 0xab
      12'h559: dout  = 8'b11110000; // 1369 : 240 - 0xf0
      12'h55A: dout  = 8'b11111000; // 1370 : 248 - 0xf8
      12'h55B: dout  = 8'b11111100; // 1371 : 252 - 0xfc
      12'h55C: dout  = 8'b11111110; // 1372 : 254 - 0xfe
      12'h55D: dout  = 8'b11111110; // 1373 : 254 - 0xfe
      12'h55E: dout  = 8'b11111111; // 1374 : 255 - 0xff
      12'h55F: dout  = 8'b11111110; // 1375 : 254 - 0xfe
      12'h560: dout  = 8'b01111111; // 1376 : 127 - 0x7f -- Sprite 0xac
      12'h561: dout  = 8'b01111111; // 1377 : 127 - 0x7f
      12'h562: dout  = 8'b01111111; // 1378 : 127 - 0x7f
      12'h563: dout  = 8'b01111111; // 1379 : 127 - 0x7f
      12'h564: dout  = 8'b11111111; // 1380 : 255 - 0xff
      12'h565: dout  = 8'b00001111; // 1381 :  15 - 0xf
      12'h566: dout  = 8'b00000011; // 1382 :   3 - 0x3
      12'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout  = 8'b11111110; // 1384 : 254 - 0xfe -- Sprite 0xad
      12'h569: dout  = 8'b11111011; // 1385 : 251 - 0xfb
      12'h56A: dout  = 8'b11111111; // 1386 : 255 - 0xff
      12'h56B: dout  = 8'b11111111; // 1387 : 255 - 0xff
      12'h56C: dout  = 8'b11110110; // 1388 : 246 - 0xf6
      12'h56D: dout  = 8'b11100000; // 1389 : 224 - 0xe0
      12'h56E: dout  = 8'b11000000; // 1390 : 192 - 0xc0
      12'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout  = 8'b00000011; // 1393 :   3 - 0x3
      12'h572: dout  = 8'b00001111; // 1394 :  15 - 0xf
      12'h573: dout  = 8'b00011111; // 1395 :  31 - 0x1f
      12'h574: dout  = 8'b00111111; // 1396 :  63 - 0x3f
      12'h575: dout  = 8'b00111011; // 1397 :  59 - 0x3b
      12'h576: dout  = 8'b00111111; // 1398 :  63 - 0x3f
      12'h577: dout  = 8'b01111111; // 1399 : 127 - 0x7f
      12'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      12'h579: dout  = 8'b11000000; // 1401 : 192 - 0xc0
      12'h57A: dout  = 8'b11110000; // 1402 : 240 - 0xf0
      12'h57B: dout  = 8'b11111000; // 1403 : 248 - 0xf8
      12'h57C: dout  = 8'b11111100; // 1404 : 252 - 0xfc
      12'h57D: dout  = 8'b11111110; // 1405 : 254 - 0xfe
      12'h57E: dout  = 8'b11111110; // 1406 : 254 - 0xfe
      12'h57F: dout  = 8'b11111111; // 1407 : 255 - 0xff
      12'h580: dout  = 8'b01111111; // 1408 : 127 - 0x7f -- Sprite 0xb0
      12'h581: dout  = 8'b01111111; // 1409 : 127 - 0x7f
      12'h582: dout  = 8'b01111111; // 1410 : 127 - 0x7f
      12'h583: dout  = 8'b01111111; // 1411 : 127 - 0x7f
      12'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      12'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout  = 8'b00001111; // 1414 :  15 - 0xf
      12'h587: dout  = 8'b00000011; // 1415 :   3 - 0x3
      12'h588: dout  = 8'b11111110; // 1416 : 254 - 0xfe -- Sprite 0xb1
      12'h589: dout  = 8'b11111110; // 1417 : 254 - 0xfe
      12'h58A: dout  = 8'b11111011; // 1418 : 251 - 0xfb
      12'h58B: dout  = 8'b11111111; // 1419 : 255 - 0xff
      12'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      12'h58D: dout  = 8'b11110110; // 1421 : 246 - 0xf6
      12'h58E: dout  = 8'b11100000; // 1422 : 224 - 0xe0
      12'h58F: dout  = 8'b11000000; // 1423 : 192 - 0xc0
      12'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      12'h591: dout  = 8'b00000001; // 1425 :   1 - 0x1
      12'h592: dout  = 8'b00000001; // 1426 :   1 - 0x1
      12'h593: dout  = 8'b00000001; // 1427 :   1 - 0x1
      12'h594: dout  = 8'b00000001; // 1428 :   1 - 0x1
      12'h595: dout  = 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout  = 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout  = 8'b00001000; // 1431 :   8 - 0x8
      12'h598: dout  = 8'b01111000; // 1432 : 120 - 0x78 -- Sprite 0xb3
      12'h599: dout  = 8'b11110000; // 1433 : 240 - 0xf0
      12'h59A: dout  = 8'b11111000; // 1434 : 248 - 0xf8
      12'h59B: dout  = 8'b11100100; // 1435 : 228 - 0xe4
      12'h59C: dout  = 8'b11000000; // 1436 : 192 - 0xc0
      12'h59D: dout  = 8'b11001010; // 1437 : 202 - 0xca
      12'h59E: dout  = 8'b11001010; // 1438 : 202 - 0xca
      12'h59F: dout  = 8'b11000000; // 1439 : 192 - 0xc0
      12'h5A0: dout  = 8'b00001111; // 1440 :  15 - 0xf -- Sprite 0xb4
      12'h5A1: dout  = 8'b00011111; // 1441 :  31 - 0x1f
      12'h5A2: dout  = 8'b10011111; // 1442 : 159 - 0x9f
      12'h5A3: dout  = 8'b11111111; // 1443 : 255 - 0xff
      12'h5A4: dout  = 8'b11111111; // 1444 : 255 - 0xff
      12'h5A5: dout  = 8'b01111111; // 1445 : 127 - 0x7f
      12'h5A6: dout  = 8'b01110100; // 1446 : 116 - 0x74
      12'h5A7: dout  = 8'b00100000; // 1447 :  32 - 0x20
      12'h5A8: dout  = 8'b11100100; // 1448 : 228 - 0xe4 -- Sprite 0xb5
      12'h5A9: dout  = 8'b11111111; // 1449 : 255 - 0xff
      12'h5AA: dout  = 8'b11111110; // 1450 : 254 - 0xfe
      12'h5AB: dout  = 8'b11111100; // 1451 : 252 - 0xfc
      12'h5AC: dout  = 8'b10011100; // 1452 : 156 - 0x9c
      12'h5AD: dout  = 8'b00011110; // 1453 :  30 - 0x1e
      12'h5AE: dout  = 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout  = 8'b00000001; // 1457 :   1 - 0x1
      12'h5B2: dout  = 8'b00000011; // 1458 :   3 - 0x3
      12'h5B3: dout  = 8'b00000011; // 1459 :   3 - 0x3
      12'h5B4: dout  = 8'b00000111; // 1460 :   7 - 0x7
      12'h5B5: dout  = 8'b00000011; // 1461 :   3 - 0x3
      12'h5B6: dout  = 8'b00000001; // 1462 :   1 - 0x1
      12'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0 -- Sprite 0xb7
      12'h5B9: dout  = 8'b01011111; // 1465 :  95 - 0x5f
      12'h5BA: dout  = 8'b01111111; // 1466 : 127 - 0x7f
      12'h5BB: dout  = 8'b01111111; // 1467 : 127 - 0x7f
      12'h5BC: dout  = 8'b00111111; // 1468 :  63 - 0x3f
      12'h5BD: dout  = 8'b00111111; // 1469 :  63 - 0x3f
      12'h5BE: dout  = 8'b00010100; // 1470 :  20 - 0x14
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b11000000; // 1472 : 192 - 0xc0 -- Sprite 0xb8
      12'h5C1: dout  = 8'b11100000; // 1473 : 224 - 0xe0
      12'h5C2: dout  = 8'b11110000; // 1474 : 240 - 0xf0
      12'h5C3: dout  = 8'b00110000; // 1475 :  48 - 0x30
      12'h5C4: dout  = 8'b00111000; // 1476 :  56 - 0x38
      12'h5C5: dout  = 8'b00111100; // 1477 :  60 - 0x3c
      12'h5C6: dout  = 8'b00111100; // 1478 :  60 - 0x3c
      12'h5C7: dout  = 8'b11111100; // 1479 : 252 - 0xfc
      12'h5C8: dout  = 8'b00000111; // 1480 :   7 - 0x7 -- Sprite 0xb9
      12'h5C9: dout  = 8'b00001111; // 1481 :  15 - 0xf
      12'h5CA: dout  = 8'b00011111; // 1482 :  31 - 0x1f
      12'h5CB: dout  = 8'b00100010; // 1483 :  34 - 0x22
      12'h5CC: dout  = 8'b00100000; // 1484 :  32 - 0x20
      12'h5CD: dout  = 8'b00100101; // 1485 :  37 - 0x25
      12'h5CE: dout  = 8'b00100101; // 1486 :  37 - 0x25
      12'h5CF: dout  = 8'b00011111; // 1487 :  31 - 0x1f
      12'h5D0: dout  = 8'b11111110; // 1488 : 254 - 0xfe -- Sprite 0xba
      12'h5D1: dout  = 8'b11111110; // 1489 : 254 - 0xfe
      12'h5D2: dout  = 8'b01111110; // 1490 : 126 - 0x7e
      12'h5D3: dout  = 8'b00111010; // 1491 :  58 - 0x3a
      12'h5D4: dout  = 8'b00000010; // 1492 :   2 - 0x2
      12'h5D5: dout  = 8'b00000001; // 1493 :   1 - 0x1
      12'h5D6: dout  = 8'b01000001; // 1494 :  65 - 0x41
      12'h5D7: dout  = 8'b01000001; // 1495 :  65 - 0x41
      12'h5D8: dout  = 8'b00011111; // 1496 :  31 - 0x1f -- Sprite 0xbb
      12'h5D9: dout  = 8'b00111111; // 1497 :  63 - 0x3f
      12'h5DA: dout  = 8'b01111110; // 1498 : 126 - 0x7e
      12'h5DB: dout  = 8'b01011100; // 1499 :  92 - 0x5c
      12'h5DC: dout  = 8'b01000000; // 1500 :  64 - 0x40
      12'h5DD: dout  = 8'b10000000; // 1501 : 128 - 0x80
      12'h5DE: dout  = 8'b10000010; // 1502 : 130 - 0x82
      12'h5DF: dout  = 8'b10000010; // 1503 : 130 - 0x82
      12'h5E0: dout  = 8'b10000010; // 1504 : 130 - 0x82 -- Sprite 0xbc
      12'h5E1: dout  = 8'b10000000; // 1505 : 128 - 0x80
      12'h5E2: dout  = 8'b10100000; // 1506 : 160 - 0xa0
      12'h5E3: dout  = 8'b01000100; // 1507 :  68 - 0x44
      12'h5E4: dout  = 8'b01000011; // 1508 :  67 - 0x43
      12'h5E5: dout  = 8'b01000000; // 1509 :  64 - 0x40
      12'h5E6: dout  = 8'b00100001; // 1510 :  33 - 0x21
      12'h5E7: dout  = 8'b00011110; // 1511 :  30 - 0x1e
      12'h5E8: dout  = 8'b00011100; // 1512 :  28 - 0x1c -- Sprite 0xbd
      12'h5E9: dout  = 8'b00111111; // 1513 :  63 - 0x3f
      12'h5EA: dout  = 8'b00111110; // 1514 :  62 - 0x3e
      12'h5EB: dout  = 8'b00111100; // 1515 :  60 - 0x3c
      12'h5EC: dout  = 8'b01000000; // 1516 :  64 - 0x40
      12'h5ED: dout  = 8'b10000000; // 1517 : 128 - 0x80
      12'h5EE: dout  = 8'b10000010; // 1518 : 130 - 0x82
      12'h5EF: dout  = 8'b10000010; // 1519 : 130 - 0x82
      12'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout  = 8'b10000000; // 1522 : 128 - 0x80
      12'h5F3: dout  = 8'b10000000; // 1523 : 128 - 0x80
      12'h5F4: dout  = 8'b10010010; // 1524 : 146 - 0x92
      12'h5F5: dout  = 8'b10011101; // 1525 : 157 - 0x9d
      12'h5F6: dout  = 8'b11000111; // 1526 : 199 - 0xc7
      12'h5F7: dout  = 8'b11101111; // 1527 : 239 - 0xef
      12'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout  = 8'b00100011; // 1529 :  35 - 0x23
      12'h5FA: dout  = 8'b00110011; // 1530 :  51 - 0x33
      12'h5FB: dout  = 8'b00111111; // 1531 :  63 - 0x3f
      12'h5FC: dout  = 8'b00111111; // 1532 :  63 - 0x3f
      12'h5FD: dout  = 8'b01111111; // 1533 : 127 - 0x7f
      12'h5FE: dout  = 8'b01111111; // 1534 : 127 - 0x7f
      12'h5FF: dout  = 8'b01111111; // 1535 : 127 - 0x7f
      12'h600: dout  = 8'b11111110; // 1536 : 254 - 0xfe -- Sprite 0xc0
      12'h601: dout  = 8'b11111000; // 1537 : 248 - 0xf8
      12'h602: dout  = 8'b10100000; // 1538 : 160 - 0xa0
      12'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout  = 8'b10000000; // 1542 : 128 - 0x80
      12'h607: dout  = 8'b10000000; // 1543 : 128 - 0x80
      12'h608: dout  = 8'b01111110; // 1544 : 126 - 0x7e -- Sprite 0xc1
      12'h609: dout  = 8'b01111111; // 1545 : 127 - 0x7f
      12'h60A: dout  = 8'b01111101; // 1546 : 125 - 0x7d
      12'h60B: dout  = 8'b00111111; // 1547 :  63 - 0x3f
      12'h60C: dout  = 8'b00011110; // 1548 :  30 - 0x1e
      12'h60D: dout  = 8'b10001111; // 1549 : 143 - 0x8f
      12'h60E: dout  = 8'b10001111; // 1550 : 143 - 0x8f
      12'h60F: dout  = 8'b00011001; // 1551 :  25 - 0x19
      12'h610: dout  = 8'b11100000; // 1552 : 224 - 0xe0 -- Sprite 0xc2
      12'h611: dout  = 8'b00001110; // 1553 :  14 - 0xe
      12'h612: dout  = 8'b01110011; // 1554 : 115 - 0x73
      12'h613: dout  = 8'b11110011; // 1555 : 243 - 0xf3
      12'h614: dout  = 8'b11111001; // 1556 : 249 - 0xf9
      12'h615: dout  = 8'b11111001; // 1557 : 249 - 0xf9
      12'h616: dout  = 8'b11111000; // 1558 : 248 - 0xf8
      12'h617: dout  = 8'b01110000; // 1559 : 112 - 0x70
      12'h618: dout  = 8'b00001110; // 1560 :  14 - 0xe -- Sprite 0xc3
      12'h619: dout  = 8'b01100110; // 1561 : 102 - 0x66
      12'h61A: dout  = 8'b11100010; // 1562 : 226 - 0xe2
      12'h61B: dout  = 8'b11110110; // 1563 : 246 - 0xf6
      12'h61C: dout  = 8'b11111111; // 1564 : 255 - 0xff
      12'h61D: dout  = 8'b11111111; // 1565 : 255 - 0xff
      12'h61E: dout  = 8'b00011111; // 1566 :  31 - 0x1f
      12'h61F: dout  = 8'b10011000; // 1567 : 152 - 0x98
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout  = 8'b00000100; // 1571 :   4 - 0x4
      12'h624: dout  = 8'b00001111; // 1572 :  15 - 0xf
      12'h625: dout  = 8'b00001111; // 1573 :  15 - 0xf
      12'h626: dout  = 8'b00011111; // 1574 :  31 - 0x1f
      12'h627: dout  = 8'b00000111; // 1575 :   7 - 0x7
      12'h628: dout  = 8'b11110011; // 1576 : 243 - 0xf3 -- Sprite 0xc5
      12'h629: dout  = 8'b11100111; // 1577 : 231 - 0xe7
      12'h62A: dout  = 8'b11101110; // 1578 : 238 - 0xee
      12'h62B: dout  = 8'b11101100; // 1579 : 236 - 0xec
      12'h62C: dout  = 8'b11001101; // 1580 : 205 - 0xcd
      12'h62D: dout  = 8'b11001111; // 1581 : 207 - 0xcf
      12'h62E: dout  = 8'b11001111; // 1582 : 207 - 0xcf
      12'h62F: dout  = 8'b11011111; // 1583 : 223 - 0xdf
      12'h630: dout  = 8'b00100111; // 1584 :  39 - 0x27 -- Sprite 0xc6
      12'h631: dout  = 8'b00111111; // 1585 :  63 - 0x3f
      12'h632: dout  = 8'b00111111; // 1586 :  63 - 0x3f
      12'h633: dout  = 8'b01111000; // 1587 : 120 - 0x78
      12'h634: dout  = 8'b00111100; // 1588 :  60 - 0x3c
      12'h635: dout  = 8'b00011111; // 1589 :  31 - 0x1f
      12'h636: dout  = 8'b00011111; // 1590 :  31 - 0x1f
      12'h637: dout  = 8'b01110011; // 1591 : 115 - 0x73
      12'h638: dout  = 8'b10011111; // 1592 : 159 - 0x9f -- Sprite 0xc7
      12'h639: dout  = 8'b00111110; // 1593 :  62 - 0x3e
      12'h63A: dout  = 8'b01111100; // 1594 : 124 - 0x7c
      12'h63B: dout  = 8'b11111100; // 1595 : 252 - 0xfc
      12'h63C: dout  = 8'b11111000; // 1596 : 248 - 0xf8
      12'h63D: dout  = 8'b11111000; // 1597 : 248 - 0xf8
      12'h63E: dout  = 8'b11000000; // 1598 : 192 - 0xc0
      12'h63F: dout  = 8'b01000000; // 1599 :  64 - 0x40
      12'h640: dout  = 8'b01111111; // 1600 : 127 - 0x7f -- Sprite 0xc8
      12'h641: dout  = 8'b01111110; // 1601 : 126 - 0x7e
      12'h642: dout  = 8'b01111000; // 1602 : 120 - 0x78
      12'h643: dout  = 8'b00000001; // 1603 :   1 - 0x1
      12'h644: dout  = 8'b00000111; // 1604 :   7 - 0x7
      12'h645: dout  = 8'b00011111; // 1605 :  31 - 0x1f
      12'h646: dout  = 8'b00111100; // 1606 :  60 - 0x3c
      12'h647: dout  = 8'b01111100; // 1607 : 124 - 0x7c
      12'h648: dout  = 8'b11111100; // 1608 : 252 - 0xfc -- Sprite 0xc9
      12'h649: dout  = 8'b11111000; // 1609 : 248 - 0xf8
      12'h64A: dout  = 8'b10100000; // 1610 : 160 - 0xa0
      12'h64B: dout  = 8'b11111110; // 1611 : 254 - 0xfe
      12'h64C: dout  = 8'b11111100; // 1612 : 252 - 0xfc
      12'h64D: dout  = 8'b11110000; // 1613 : 240 - 0xf0
      12'h64E: dout  = 8'b10000000; // 1614 : 128 - 0x80
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b01111110; // 1616 : 126 - 0x7e -- Sprite 0xca
      12'h651: dout  = 8'b01111111; // 1617 : 127 - 0x7f
      12'h652: dout  = 8'b01111111; // 1618 : 127 - 0x7f
      12'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      12'h654: dout  = 8'b00011111; // 1620 :  31 - 0x1f
      12'h655: dout  = 8'b10001111; // 1621 : 143 - 0x8f
      12'h656: dout  = 8'b10001111; // 1622 : 143 - 0x8f
      12'h657: dout  = 8'b00011000; // 1623 :  24 - 0x18
      12'h658: dout  = 8'b10011111; // 1624 : 159 - 0x9f -- Sprite 0xcb
      12'h659: dout  = 8'b00111110; // 1625 :  62 - 0x3e
      12'h65A: dout  = 8'b01111100; // 1626 : 124 - 0x7c
      12'h65B: dout  = 8'b11111000; // 1627 : 248 - 0xf8
      12'h65C: dout  = 8'b11111000; // 1628 : 248 - 0xf8
      12'h65D: dout  = 8'b00111100; // 1629 :  60 - 0x3c
      12'h65E: dout  = 8'b00011000; // 1630 :  24 - 0x18
      12'h65F: dout  = 8'b11111000; // 1631 : 248 - 0xf8
      12'h660: dout  = 8'b01111111; // 1632 : 127 - 0x7f -- Sprite 0xcc
      12'h661: dout  = 8'b01111111; // 1633 : 127 - 0x7f
      12'h662: dout  = 8'b01111000; // 1634 : 120 - 0x78
      12'h663: dout  = 8'b00000001; // 1635 :   1 - 0x1
      12'h664: dout  = 8'b00000111; // 1636 :   7 - 0x7
      12'h665: dout  = 8'b00010011; // 1637 :  19 - 0x13
      12'h666: dout  = 8'b11110001; // 1638 : 241 - 0xf1
      12'h667: dout  = 8'b00000011; // 1639 :   3 - 0x3
      12'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout  = 8'b00011100; // 1642 :  28 - 0x1c
      12'h66B: dout  = 8'b00011101; // 1643 :  29 - 0x1d
      12'h66C: dout  = 8'b00011011; // 1644 :  27 - 0x1b
      12'h66D: dout  = 8'b11000011; // 1645 : 195 - 0xc3
      12'h66E: dout  = 8'b11100011; // 1646 : 227 - 0xe3
      12'h66F: dout  = 8'b11100001; // 1647 : 225 - 0xe1
      12'h670: dout  = 8'b11100000; // 1648 : 224 - 0xe0 -- Sprite 0xce
      12'h671: dout  = 8'b11001101; // 1649 : 205 - 0xcd
      12'h672: dout  = 8'b00011101; // 1650 :  29 - 0x1d
      12'h673: dout  = 8'b01001111; // 1651 :  79 - 0x4f
      12'h674: dout  = 8'b11101110; // 1652 : 238 - 0xee
      12'h675: dout  = 8'b11111111; // 1653 : 255 - 0xff
      12'h676: dout  = 8'b00111111; // 1654 :  63 - 0x3f
      12'h677: dout  = 8'b00111111; // 1655 :  63 - 0x3f
      12'h678: dout  = 8'b00111111; // 1656 :  63 - 0x3f -- Sprite 0xcf
      12'h679: dout  = 8'b00111111; // 1657 :  63 - 0x3f
      12'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout  = 8'b01110000; // 1660 : 112 - 0x70
      12'h67D: dout  = 8'b10111000; // 1661 : 184 - 0xb8
      12'h67E: dout  = 8'b11111100; // 1662 : 252 - 0xfc
      12'h67F: dout  = 8'b11111100; // 1663 : 252 - 0xfc
      12'h680: dout  = 8'b00000111; // 1664 :   7 - 0x7 -- Sprite 0xd0
      12'h681: dout  = 8'b00001111; // 1665 :  15 - 0xf
      12'h682: dout  = 8'b00011111; // 1666 :  31 - 0x1f
      12'h683: dout  = 8'b00111111; // 1667 :  63 - 0x3f
      12'h684: dout  = 8'b00111110; // 1668 :  62 - 0x3e
      12'h685: dout  = 8'b01111100; // 1669 : 124 - 0x7c
      12'h686: dout  = 8'b01111000; // 1670 : 120 - 0x78
      12'h687: dout  = 8'b01111000; // 1671 : 120 - 0x78
      12'h688: dout  = 8'b00111111; // 1672 :  63 - 0x3f -- Sprite 0xd1
      12'h689: dout  = 8'b01011100; // 1673 :  92 - 0x5c
      12'h68A: dout  = 8'b00111001; // 1674 :  57 - 0x39
      12'h68B: dout  = 8'b00111011; // 1675 :  59 - 0x3b
      12'h68C: dout  = 8'b10111111; // 1676 : 191 - 0xbf
      12'h68D: dout  = 8'b11111111; // 1677 : 255 - 0xff
      12'h68E: dout  = 8'b11111110; // 1678 : 254 - 0xfe
      12'h68F: dout  = 8'b11111110; // 1679 : 254 - 0xfe
      12'h690: dout  = 8'b11000000; // 1680 : 192 - 0xc0 -- Sprite 0xd2
      12'h691: dout  = 8'b11000000; // 1681 : 192 - 0xc0
      12'h692: dout  = 8'b10000000; // 1682 : 128 - 0x80
      12'h693: dout  = 8'b10000000; // 1683 : 128 - 0x80
      12'h694: dout  = 8'b10000000; // 1684 : 128 - 0x80
      12'h695: dout  = 8'b10000000; // 1685 : 128 - 0x80
      12'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout  = 8'b11111110; // 1688 : 254 - 0xfe -- Sprite 0xd3
      12'h699: dout  = 8'b11111100; // 1689 : 252 - 0xfc
      12'h69A: dout  = 8'b01100001; // 1690 :  97 - 0x61
      12'h69B: dout  = 8'b00001111; // 1691 :  15 - 0xf
      12'h69C: dout  = 8'b01111111; // 1692 : 127 - 0x7f
      12'h69D: dout  = 8'b00111111; // 1693 :  63 - 0x3f
      12'h69E: dout  = 8'b00011111; // 1694 :  31 - 0x1f
      12'h69F: dout  = 8'b00011110; // 1695 :  30 - 0x1e
      12'h6A0: dout  = 8'b11110000; // 1696 : 240 - 0xf0 -- Sprite 0xd4
      12'h6A1: dout  = 8'b01111000; // 1697 : 120 - 0x78
      12'h6A2: dout  = 8'b11100100; // 1698 : 228 - 0xe4
      12'h6A3: dout  = 8'b11001000; // 1699 : 200 - 0xc8
      12'h6A4: dout  = 8'b11001100; // 1700 : 204 - 0xcc
      12'h6A5: dout  = 8'b10111110; // 1701 : 190 - 0xbe
      12'h6A6: dout  = 8'b10111110; // 1702 : 190 - 0xbe
      12'h6A7: dout  = 8'b00111110; // 1703 :  62 - 0x3e
      12'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      12'h6A9: dout  = 8'b00000001; // 1705 :   1 - 0x1
      12'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout  = 8'b00000111; // 1707 :   7 - 0x7
      12'h6AC: dout  = 8'b00000111; // 1708 :   7 - 0x7
      12'h6AD: dout  = 8'b00000111; // 1709 :   7 - 0x7
      12'h6AE: dout  = 8'b00000111; // 1710 :   7 - 0x7
      12'h6AF: dout  = 8'b00011111; // 1711 :  31 - 0x1f
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout  = 8'b00001111; // 1714 :  15 - 0xf
      12'h6B3: dout  = 8'b00111111; // 1715 :  63 - 0x3f
      12'h6B4: dout  = 8'b00111111; // 1716 :  63 - 0x3f
      12'h6B5: dout  = 8'b00001111; // 1717 :  15 - 0xf
      12'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout  = 8'b01111000; // 1720 : 120 - 0x78 -- Sprite 0xd7
      12'h6B9: dout  = 8'b01111100; // 1721 : 124 - 0x7c
      12'h6BA: dout  = 8'b01111110; // 1722 : 126 - 0x7e
      12'h6BB: dout  = 8'b01111111; // 1723 : 127 - 0x7f
      12'h6BC: dout  = 8'b00111111; // 1724 :  63 - 0x3f
      12'h6BD: dout  = 8'b00111111; // 1725 :  63 - 0x3f
      12'h6BE: dout  = 8'b00011011; // 1726 :  27 - 0x1b
      12'h6BF: dout  = 8'b00001001; // 1727 :   9 - 0x9
      12'h6C0: dout  = 8'b00001100; // 1728 :  12 - 0xc -- Sprite 0xd8
      12'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout  = 8'b00000111; // 1732 :   7 - 0x7
      12'h6C5: dout  = 8'b01111111; // 1733 : 127 - 0x7f
      12'h6C6: dout  = 8'b01111100; // 1734 : 124 - 0x7c
      12'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout  = 8'b00000001; // 1736 :   1 - 0x1 -- Sprite 0xd9
      12'h6C9: dout  = 8'b11100001; // 1737 : 225 - 0xe1
      12'h6CA: dout  = 8'b01110001; // 1738 : 113 - 0x71
      12'h6CB: dout  = 8'b01111001; // 1739 : 121 - 0x79
      12'h6CC: dout  = 8'b00111101; // 1740 :  61 - 0x3d
      12'h6CD: dout  = 8'b00111101; // 1741 :  61 - 0x3d
      12'h6CE: dout  = 8'b00011111; // 1742 :  31 - 0x1f
      12'h6CF: dout  = 8'b00000011; // 1743 :   3 - 0x3
      12'h6D0: dout  = 8'b00111111; // 1744 :  63 - 0x3f -- Sprite 0xda
      12'h6D1: dout  = 8'b00111111; // 1745 :  63 - 0x3f
      12'h6D2: dout  = 8'b00011111; // 1746 :  31 - 0x1f
      12'h6D3: dout  = 8'b00011011; // 1747 :  27 - 0x1b
      12'h6D4: dout  = 8'b00110110; // 1748 :  54 - 0x36
      12'h6D5: dout  = 8'b00110000; // 1749 :  48 - 0x30
      12'h6D6: dout  = 8'b01111111; // 1750 : 127 - 0x7f
      12'h6D7: dout  = 8'b00111111; // 1751 :  63 - 0x3f
      12'h6D8: dout  = 8'b11111000; // 1752 : 248 - 0xf8 -- Sprite 0xdb
      12'h6D9: dout  = 8'b11111000; // 1753 : 248 - 0xf8
      12'h6DA: dout  = 8'b11111000; // 1754 : 248 - 0xf8
      12'h6DB: dout  = 8'b10111000; // 1755 : 184 - 0xb8
      12'h6DC: dout  = 8'b00011000; // 1756 :  24 - 0x18
      12'h6DD: dout  = 8'b11011000; // 1757 : 216 - 0xd8
      12'h6DE: dout  = 8'b11011000; // 1758 : 216 - 0xd8
      12'h6DF: dout  = 8'b10111000; // 1759 : 184 - 0xb8
      12'h6E0: dout  = 8'b00000001; // 1760 :   1 - 0x1 -- Sprite 0xdc
      12'h6E1: dout  = 8'b00000010; // 1761 :   2 - 0x2
      12'h6E2: dout  = 8'b00000100; // 1762 :   4 - 0x4
      12'h6E3: dout  = 8'b00000100; // 1763 :   4 - 0x4
      12'h6E4: dout  = 8'b00001000; // 1764 :   8 - 0x8
      12'h6E5: dout  = 8'b00001000; // 1765 :   8 - 0x8
      12'h6E6: dout  = 8'b00010000; // 1766 :  16 - 0x10
      12'h6E7: dout  = 8'b00010000; // 1767 :  16 - 0x10
      12'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      12'h6E9: dout  = 8'b00001111; // 1769 :  15 - 0xf
      12'h6EA: dout  = 8'b00010011; // 1770 :  19 - 0x13
      12'h6EB: dout  = 8'b00001101; // 1771 :  13 - 0xd
      12'h6EC: dout  = 8'b00001101; // 1772 :  13 - 0xd
      12'h6ED: dout  = 8'b00010011; // 1773 :  19 - 0x13
      12'h6EE: dout  = 8'b00001100; // 1774 :  12 - 0xc
      12'h6EF: dout  = 8'b00100000; // 1775 :  32 - 0x20
      12'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0xde
      12'h6F1: dout  = 8'b00100100; // 1777 :  36 - 0x24
      12'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout  = 8'b00100100; // 1779 :  36 - 0x24
      12'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout  = 8'b00000100; // 1781 :   4 - 0x4
      12'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout  = 8'b00001111; // 1784 :  15 - 0xf -- Sprite 0xdf
      12'h6F9: dout  = 8'b01000001; // 1785 :  65 - 0x41
      12'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout  = 8'b10001000; // 1787 : 136 - 0x88
      12'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout  = 8'b01000100; // 1789 :  68 - 0x44
      12'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout  = 8'b00111000; // 1792 :  56 - 0x38 -- Sprite 0xe0
      12'h701: dout  = 8'b01111100; // 1793 : 124 - 0x7c
      12'h702: dout  = 8'b11111110; // 1794 : 254 - 0xfe
      12'h703: dout  = 8'b11111110; // 1795 : 254 - 0xfe
      12'h704: dout  = 8'b00111011; // 1796 :  59 - 0x3b
      12'h705: dout  = 8'b00000011; // 1797 :   3 - 0x3
      12'h706: dout  = 8'b00000011; // 1798 :   3 - 0x3
      12'h707: dout  = 8'b00000011; // 1799 :   3 - 0x3
      12'h708: dout  = 8'b00000011; // 1800 :   3 - 0x3 -- Sprite 0xe1
      12'h709: dout  = 8'b00110011; // 1801 :  51 - 0x33
      12'h70A: dout  = 8'b01111011; // 1802 : 123 - 0x7b
      12'h70B: dout  = 8'b01111111; // 1803 : 127 - 0x7f
      12'h70C: dout  = 8'b11111111; // 1804 : 255 - 0xff
      12'h70D: dout  = 8'b11111011; // 1805 : 251 - 0xfb
      12'h70E: dout  = 8'b00000011; // 1806 :   3 - 0x3
      12'h70F: dout  = 8'b00000011; // 1807 :   3 - 0x3
      12'h710: dout  = 8'b11011100; // 1808 : 220 - 0xdc -- Sprite 0xe2
      12'h711: dout  = 8'b11000000; // 1809 : 192 - 0xc0
      12'h712: dout  = 8'b11100000; // 1810 : 224 - 0xe0
      12'h713: dout  = 8'b11100000; // 1811 : 224 - 0xe0
      12'h714: dout  = 8'b11100000; // 1812 : 224 - 0xe0
      12'h715: dout  = 8'b11100000; // 1813 : 224 - 0xe0
      12'h716: dout  = 8'b11100000; // 1814 : 224 - 0xe0
      12'h717: dout  = 8'b11000000; // 1815 : 192 - 0xc0
      12'h718: dout  = 8'b00111111; // 1816 :  63 - 0x3f -- Sprite 0xe3
      12'h719: dout  = 8'b01011111; // 1817 :  95 - 0x5f
      12'h71A: dout  = 8'b00111111; // 1818 :  63 - 0x3f
      12'h71B: dout  = 8'b00111111; // 1819 :  63 - 0x3f
      12'h71C: dout  = 8'b10111011; // 1820 : 187 - 0xbb
      12'h71D: dout  = 8'b11111000; // 1821 : 248 - 0xf8
      12'h71E: dout  = 8'b11111110; // 1822 : 254 - 0xfe
      12'h71F: dout  = 8'b11111110; // 1823 : 254 - 0xfe
      12'h720: dout  = 8'b00011111; // 1824 :  31 - 0x1f -- Sprite 0xe4
      12'h721: dout  = 8'b00001111; // 1825 :  15 - 0xf
      12'h722: dout  = 8'b00001111; // 1826 :  15 - 0xf
      12'h723: dout  = 8'b00011111; // 1827 :  31 - 0x1f
      12'h724: dout  = 8'b00011111; // 1828 :  31 - 0x1f
      12'h725: dout  = 8'b00011110; // 1829 :  30 - 0x1e
      12'h726: dout  = 8'b00111000; // 1830 :  56 - 0x38
      12'h727: dout  = 8'b00110000; // 1831 :  48 - 0x30
      12'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      12'h729: dout  = 8'b00100000; // 1833 :  32 - 0x20
      12'h72A: dout  = 8'b01100000; // 1834 :  96 - 0x60
      12'h72B: dout  = 8'b01100000; // 1835 :  96 - 0x60
      12'h72C: dout  = 8'b01110000; // 1836 : 112 - 0x70
      12'h72D: dout  = 8'b11110000; // 1837 : 240 - 0xf0
      12'h72E: dout  = 8'b11111000; // 1838 : 248 - 0xf8
      12'h72F: dout  = 8'b11111000; // 1839 : 248 - 0xf8
      12'h730: dout  = 8'b11111000; // 1840 : 248 - 0xf8 -- Sprite 0xe6
      12'h731: dout  = 8'b11111100; // 1841 : 252 - 0xfc
      12'h732: dout  = 8'b11111100; // 1842 : 252 - 0xfc
      12'h733: dout  = 8'b01111110; // 1843 : 126 - 0x7e
      12'h734: dout  = 8'b01111110; // 1844 : 126 - 0x7e
      12'h735: dout  = 8'b00111110; // 1845 :  62 - 0x3e
      12'h736: dout  = 8'b00011111; // 1846 :  31 - 0x1f
      12'h737: dout  = 8'b00000111; // 1847 :   7 - 0x7
      12'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      12'h739: dout  = 8'b11000000; // 1849 : 192 - 0xc0
      12'h73A: dout  = 8'b01110000; // 1850 : 112 - 0x70
      12'h73B: dout  = 8'b10111000; // 1851 : 184 - 0xb8
      12'h73C: dout  = 8'b11110100; // 1852 : 244 - 0xf4
      12'h73D: dout  = 8'b11110010; // 1853 : 242 - 0xf2
      12'h73E: dout  = 8'b11110101; // 1854 : 245 - 0xf5
      12'h73F: dout  = 8'b01111011; // 1855 : 123 - 0x7b
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout  = 8'b11011111; // 1857 : 223 - 0xdf
      12'h742: dout  = 8'b00010000; // 1858 :  16 - 0x10
      12'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout  = 8'b11011111; // 1860 : 223 - 0xdf
      12'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout  = 8'b11111001; // 1863 : 249 - 0xf9
      12'h748: dout  = 8'b00011111; // 1864 :  31 - 0x1f -- Sprite 0xe9
      12'h749: dout  = 8'b00011111; // 1865 :  31 - 0x1f
      12'h74A: dout  = 8'b00111110; // 1866 :  62 - 0x3e
      12'h74B: dout  = 8'b11111100; // 1867 : 252 - 0xfc
      12'h74C: dout  = 8'b11111000; // 1868 : 248 - 0xf8
      12'h74D: dout  = 8'b11110000; // 1869 : 240 - 0xf0
      12'h74E: dout  = 8'b11000000; // 1870 : 192 - 0xc0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b11111000; // 1872 : 248 - 0xf8 -- Sprite 0xea
      12'h751: dout  = 8'b11111100; // 1873 : 252 - 0xfc
      12'h752: dout  = 8'b11111110; // 1874 : 254 - 0xfe
      12'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout  = 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout  = 8'b11011111; // 1877 : 223 - 0xdf
      12'h756: dout  = 8'b11011111; // 1878 : 223 - 0xdf
      12'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout  = 8'b11000001; // 1880 : 193 - 0xc1 -- Sprite 0xeb
      12'h759: dout  = 8'b11110001; // 1881 : 241 - 0xf1
      12'h75A: dout  = 8'b01111001; // 1882 : 121 - 0x79
      12'h75B: dout  = 8'b01111101; // 1883 : 125 - 0x7d
      12'h75C: dout  = 8'b00111101; // 1884 :  61 - 0x3d
      12'h75D: dout  = 8'b00111111; // 1885 :  63 - 0x3f
      12'h75E: dout  = 8'b00011111; // 1886 :  31 - 0x1f
      12'h75F: dout  = 8'b00000011; // 1887 :   3 - 0x3
      12'h760: dout  = 8'b00000010; // 1888 :   2 - 0x2 -- Sprite 0xec
      12'h761: dout  = 8'b00000110; // 1889 :   6 - 0x6
      12'h762: dout  = 8'b00001110; // 1890 :  14 - 0xe
      12'h763: dout  = 8'b00001110; // 1891 :  14 - 0xe
      12'h764: dout  = 8'b00011110; // 1892 :  30 - 0x1e
      12'h765: dout  = 8'b00011110; // 1893 :  30 - 0x1e
      12'h766: dout  = 8'b00111110; // 1894 :  62 - 0x3e
      12'h767: dout  = 8'b00111110; // 1895 :  62 - 0x3e
      12'h768: dout  = 8'b00111110; // 1896 :  62 - 0x3e -- Sprite 0xed
      12'h769: dout  = 8'b00111110; // 1897 :  62 - 0x3e
      12'h76A: dout  = 8'b00111110; // 1898 :  62 - 0x3e
      12'h76B: dout  = 8'b00111110; // 1899 :  62 - 0x3e
      12'h76C: dout  = 8'b00011110; // 1900 :  30 - 0x1e
      12'h76D: dout  = 8'b00011110; // 1901 :  30 - 0x1e
      12'h76E: dout  = 8'b00001110; // 1902 :  14 - 0xe
      12'h76F: dout  = 8'b00000010; // 1903 :   2 - 0x2
      12'h770: dout  = 8'b11000001; // 1904 : 193 - 0xc1 -- Sprite 0xee
      12'h771: dout  = 8'b11110001; // 1905 : 241 - 0xf1
      12'h772: dout  = 8'b01111001; // 1906 : 121 - 0x79
      12'h773: dout  = 8'b01111101; // 1907 : 125 - 0x7d
      12'h774: dout  = 8'b00111101; // 1908 :  61 - 0x3d
      12'h775: dout  = 8'b00111111; // 1909 :  63 - 0x3f
      12'h776: dout  = 8'b00011111; // 1910 :  31 - 0x1f
      12'h777: dout  = 8'b00000011; // 1911 :   3 - 0x3
      12'h778: dout  = 8'b01111100; // 1912 : 124 - 0x7c -- Sprite 0xef
      12'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout  = 8'b11000011; // 1916 : 195 - 0xc3
      12'h77D: dout  = 8'b01111111; // 1917 : 127 - 0x7f
      12'h77E: dout  = 8'b00011111; // 1918 :  31 - 0x1f
      12'h77F: dout  = 8'b00000011; // 1919 :   3 - 0x3
      12'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0xf0
      12'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout  = 8'b01111100; // 1922 : 124 - 0x7c
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b01111100; // 1925 : 124 - 0x7c
      12'h786: dout  = 8'b11111111; // 1926 : 255 - 0xff
      12'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      12'h789: dout  = 8'b11111111; // 1929 : 255 - 0xff
      12'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout  = 8'b00000100; // 1931 :   4 - 0x4
      12'h78C: dout  = 8'b00001100; // 1932 :  12 - 0xc
      12'h78D: dout  = 8'b00011000; // 1933 :  24 - 0x18
      12'h78E: dout  = 8'b00110000; // 1934 :  48 - 0x30
      12'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0xf2
      12'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout  = 8'b00000100; // 1939 :   4 - 0x4
      12'h794: dout  = 8'b00000100; // 1940 :   4 - 0x4
      12'h795: dout  = 8'b00000100; // 1941 :   4 - 0x4
      12'h796: dout  = 8'b00001000; // 1942 :   8 - 0x8
      12'h797: dout  = 8'b00001000; // 1943 :   8 - 0x8
      12'h798: dout  = 8'b00001000; // 1944 :   8 - 0x8 -- Sprite 0xf3
      12'h799: dout  = 8'b00010000; // 1945 :  16 - 0x10
      12'h79A: dout  = 8'b00010000; // 1946 :  16 - 0x10
      12'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout  = 8'b00010000; // 1949 :  16 - 0x10
      12'h79E: dout  = 8'b00010000; // 1950 :  16 - 0x10
      12'h79F: dout  = 8'b00001000; // 1951 :   8 - 0x8
      12'h7A0: dout  = 8'b01111111; // 1952 : 127 - 0x7f -- Sprite 0xf4
      12'h7A1: dout  = 8'b00111111; // 1953 :  63 - 0x3f
      12'h7A2: dout  = 8'b00111111; // 1954 :  63 - 0x3f
      12'h7A3: dout  = 8'b00111110; // 1955 :  62 - 0x3e
      12'h7A4: dout  = 8'b00011111; // 1956 :  31 - 0x1f
      12'h7A5: dout  = 8'b00001111; // 1957 :  15 - 0xf
      12'h7A6: dout  = 8'b00000011; // 1958 :   3 - 0x3
      12'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout  = 8'b00000011; // 1960 :   3 - 0x3 -- Sprite 0xf5
      12'h7A9: dout  = 8'b00001111; // 1961 :  15 - 0xf
      12'h7AA: dout  = 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout  = 8'b01111111; // 1963 : 127 - 0x7f
      12'h7AC: dout  = 8'b01111111; // 1964 : 127 - 0x7f
      12'h7AD: dout  = 8'b01111111; // 1965 : 127 - 0x7f
      12'h7AE: dout  = 8'b01111111; // 1966 : 127 - 0x7f
      12'h7AF: dout  = 8'b01111111; // 1967 : 127 - 0x7f
      12'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      12'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      12'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      12'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      12'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      12'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      12'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      12'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout  = 8'b01111100; // 2045 : 124 - 0x7c
      12'h7FE: dout  = 8'b00111000; // 2046 :  56 - 0x38
      12'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
          // Background pattern Table
      12'h800: dout  = 8'b00111000; // 2048 :  56 - 0x38 -- Background 0x0
      12'h801: dout  = 8'b01001100; // 2049 :  76 - 0x4c
      12'h802: dout  = 8'b11000110; // 2050 : 198 - 0xc6
      12'h803: dout  = 8'b11000110; // 2051 : 198 - 0xc6
      12'h804: dout  = 8'b11000110; // 2052 : 198 - 0xc6
      12'h805: dout  = 8'b01100100; // 2053 : 100 - 0x64
      12'h806: dout  = 8'b00111000; // 2054 :  56 - 0x38
      12'h807: dout  = 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout  = 8'b00011000; // 2056 :  24 - 0x18 -- Background 0x1
      12'h809: dout  = 8'b00111000; // 2057 :  56 - 0x38
      12'h80A: dout  = 8'b00011000; // 2058 :  24 - 0x18
      12'h80B: dout  = 8'b00011000; // 2059 :  24 - 0x18
      12'h80C: dout  = 8'b00011000; // 2060 :  24 - 0x18
      12'h80D: dout  = 8'b00011000; // 2061 :  24 - 0x18
      12'h80E: dout  = 8'b01111110; // 2062 : 126 - 0x7e
      12'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout  = 8'b01111100; // 2064 : 124 - 0x7c -- Background 0x2
      12'h811: dout  = 8'b11000110; // 2065 : 198 - 0xc6
      12'h812: dout  = 8'b00001110; // 2066 :  14 - 0xe
      12'h813: dout  = 8'b00111100; // 2067 :  60 - 0x3c
      12'h814: dout  = 8'b01111000; // 2068 : 120 - 0x78
      12'h815: dout  = 8'b11100000; // 2069 : 224 - 0xe0
      12'h816: dout  = 8'b11111110; // 2070 : 254 - 0xfe
      12'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout  = 8'b01111110; // 2072 : 126 - 0x7e -- Background 0x3
      12'h819: dout  = 8'b00001100; // 2073 :  12 - 0xc
      12'h81A: dout  = 8'b00011000; // 2074 :  24 - 0x18
      12'h81B: dout  = 8'b00111100; // 2075 :  60 - 0x3c
      12'h81C: dout  = 8'b00000110; // 2076 :   6 - 0x6
      12'h81D: dout  = 8'b11000110; // 2077 : 198 - 0xc6
      12'h81E: dout  = 8'b01111100; // 2078 : 124 - 0x7c
      12'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout  = 8'b00011100; // 2080 :  28 - 0x1c -- Background 0x4
      12'h821: dout  = 8'b00111100; // 2081 :  60 - 0x3c
      12'h822: dout  = 8'b01101100; // 2082 : 108 - 0x6c
      12'h823: dout  = 8'b11001100; // 2083 : 204 - 0xcc
      12'h824: dout  = 8'b11111110; // 2084 : 254 - 0xfe
      12'h825: dout  = 8'b00001100; // 2085 :  12 - 0xc
      12'h826: dout  = 8'b00001100; // 2086 :  12 - 0xc
      12'h827: dout  = 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout  = 8'b11111100; // 2088 : 252 - 0xfc -- Background 0x5
      12'h829: dout  = 8'b11000000; // 2089 : 192 - 0xc0
      12'h82A: dout  = 8'b11111100; // 2090 : 252 - 0xfc
      12'h82B: dout  = 8'b00000110; // 2091 :   6 - 0x6
      12'h82C: dout  = 8'b00000110; // 2092 :   6 - 0x6
      12'h82D: dout  = 8'b11000110; // 2093 : 198 - 0xc6
      12'h82E: dout  = 8'b01111100; // 2094 : 124 - 0x7c
      12'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout  = 8'b00111100; // 2096 :  60 - 0x3c -- Background 0x6
      12'h831: dout  = 8'b01100000; // 2097 :  96 - 0x60
      12'h832: dout  = 8'b11000000; // 2098 : 192 - 0xc0
      12'h833: dout  = 8'b11111100; // 2099 : 252 - 0xfc
      12'h834: dout  = 8'b11000110; // 2100 : 198 - 0xc6
      12'h835: dout  = 8'b11000110; // 2101 : 198 - 0xc6
      12'h836: dout  = 8'b01111100; // 2102 : 124 - 0x7c
      12'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout  = 8'b11111110; // 2104 : 254 - 0xfe -- Background 0x7
      12'h839: dout  = 8'b11000110; // 2105 : 198 - 0xc6
      12'h83A: dout  = 8'b00001100; // 2106 :  12 - 0xc
      12'h83B: dout  = 8'b00011000; // 2107 :  24 - 0x18
      12'h83C: dout  = 8'b00110000; // 2108 :  48 - 0x30
      12'h83D: dout  = 8'b00110000; // 2109 :  48 - 0x30
      12'h83E: dout  = 8'b00110000; // 2110 :  48 - 0x30
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b01111100; // 2112 : 124 - 0x7c -- Background 0x8
      12'h841: dout  = 8'b11000110; // 2113 : 198 - 0xc6
      12'h842: dout  = 8'b11000110; // 2114 : 198 - 0xc6
      12'h843: dout  = 8'b01111100; // 2115 : 124 - 0x7c
      12'h844: dout  = 8'b11000110; // 2116 : 198 - 0xc6
      12'h845: dout  = 8'b11000110; // 2117 : 198 - 0xc6
      12'h846: dout  = 8'b01111100; // 2118 : 124 - 0x7c
      12'h847: dout  = 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout  = 8'b01111100; // 2120 : 124 - 0x7c -- Background 0x9
      12'h849: dout  = 8'b11000110; // 2121 : 198 - 0xc6
      12'h84A: dout  = 8'b11000110; // 2122 : 198 - 0xc6
      12'h84B: dout  = 8'b01111110; // 2123 : 126 - 0x7e
      12'h84C: dout  = 8'b00000110; // 2124 :   6 - 0x6
      12'h84D: dout  = 8'b00001100; // 2125 :  12 - 0xc
      12'h84E: dout  = 8'b01111000; // 2126 : 120 - 0x78
      12'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout  = 8'b00111000; // 2128 :  56 - 0x38 -- Background 0xa
      12'h851: dout  = 8'b01101100; // 2129 : 108 - 0x6c
      12'h852: dout  = 8'b11000110; // 2130 : 198 - 0xc6
      12'h853: dout  = 8'b11000110; // 2131 : 198 - 0xc6
      12'h854: dout  = 8'b11111110; // 2132 : 254 - 0xfe
      12'h855: dout  = 8'b11000110; // 2133 : 198 - 0xc6
      12'h856: dout  = 8'b11000110; // 2134 : 198 - 0xc6
      12'h857: dout  = 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout  = 8'b11111100; // 2136 : 252 - 0xfc -- Background 0xb
      12'h859: dout  = 8'b11000110; // 2137 : 198 - 0xc6
      12'h85A: dout  = 8'b11000110; // 2138 : 198 - 0xc6
      12'h85B: dout  = 8'b11111100; // 2139 : 252 - 0xfc
      12'h85C: dout  = 8'b11000110; // 2140 : 198 - 0xc6
      12'h85D: dout  = 8'b11000110; // 2141 : 198 - 0xc6
      12'h85E: dout  = 8'b11111100; // 2142 : 252 - 0xfc
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b00111100; // 2144 :  60 - 0x3c -- Background 0xc
      12'h861: dout  = 8'b01100110; // 2145 : 102 - 0x66
      12'h862: dout  = 8'b11000000; // 2146 : 192 - 0xc0
      12'h863: dout  = 8'b11000000; // 2147 : 192 - 0xc0
      12'h864: dout  = 8'b11000000; // 2148 : 192 - 0xc0
      12'h865: dout  = 8'b01100110; // 2149 : 102 - 0x66
      12'h866: dout  = 8'b00111100; // 2150 :  60 - 0x3c
      12'h867: dout  = 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout  = 8'b11111000; // 2152 : 248 - 0xf8 -- Background 0xd
      12'h869: dout  = 8'b11001100; // 2153 : 204 - 0xcc
      12'h86A: dout  = 8'b11000110; // 2154 : 198 - 0xc6
      12'h86B: dout  = 8'b11000110; // 2155 : 198 - 0xc6
      12'h86C: dout  = 8'b11000110; // 2156 : 198 - 0xc6
      12'h86D: dout  = 8'b11001100; // 2157 : 204 - 0xcc
      12'h86E: dout  = 8'b11111000; // 2158 : 248 - 0xf8
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b11111110; // 2160 : 254 - 0xfe -- Background 0xe
      12'h871: dout  = 8'b11000000; // 2161 : 192 - 0xc0
      12'h872: dout  = 8'b11000000; // 2162 : 192 - 0xc0
      12'h873: dout  = 8'b11111100; // 2163 : 252 - 0xfc
      12'h874: dout  = 8'b11000000; // 2164 : 192 - 0xc0
      12'h875: dout  = 8'b11000000; // 2165 : 192 - 0xc0
      12'h876: dout  = 8'b11111110; // 2166 : 254 - 0xfe
      12'h877: dout  = 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout  = 8'b11111110; // 2168 : 254 - 0xfe -- Background 0xf
      12'h879: dout  = 8'b11000000; // 2169 : 192 - 0xc0
      12'h87A: dout  = 8'b11000000; // 2170 : 192 - 0xc0
      12'h87B: dout  = 8'b11111100; // 2171 : 252 - 0xfc
      12'h87C: dout  = 8'b11000000; // 2172 : 192 - 0xc0
      12'h87D: dout  = 8'b11000000; // 2173 : 192 - 0xc0
      12'h87E: dout  = 8'b11000000; // 2174 : 192 - 0xc0
      12'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout  = 8'b00111110; // 2176 :  62 - 0x3e -- Background 0x10
      12'h881: dout  = 8'b01100000; // 2177 :  96 - 0x60
      12'h882: dout  = 8'b11000000; // 2178 : 192 - 0xc0
      12'h883: dout  = 8'b11001110; // 2179 : 206 - 0xce
      12'h884: dout  = 8'b11000110; // 2180 : 198 - 0xc6
      12'h885: dout  = 8'b01100110; // 2181 : 102 - 0x66
      12'h886: dout  = 8'b00111110; // 2182 :  62 - 0x3e
      12'h887: dout  = 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout  = 8'b11000110; // 2184 : 198 - 0xc6 -- Background 0x11
      12'h889: dout  = 8'b11000110; // 2185 : 198 - 0xc6
      12'h88A: dout  = 8'b11000110; // 2186 : 198 - 0xc6
      12'h88B: dout  = 8'b11111110; // 2187 : 254 - 0xfe
      12'h88C: dout  = 8'b11000110; // 2188 : 198 - 0xc6
      12'h88D: dout  = 8'b11000110; // 2189 : 198 - 0xc6
      12'h88E: dout  = 8'b11000110; // 2190 : 198 - 0xc6
      12'h88F: dout  = 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout  = 8'b01111110; // 2192 : 126 - 0x7e -- Background 0x12
      12'h891: dout  = 8'b00011000; // 2193 :  24 - 0x18
      12'h892: dout  = 8'b00011000; // 2194 :  24 - 0x18
      12'h893: dout  = 8'b00011000; // 2195 :  24 - 0x18
      12'h894: dout  = 8'b00011000; // 2196 :  24 - 0x18
      12'h895: dout  = 8'b00011000; // 2197 :  24 - 0x18
      12'h896: dout  = 8'b01111110; // 2198 : 126 - 0x7e
      12'h897: dout  = 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout  = 8'b00011110; // 2200 :  30 - 0x1e -- Background 0x13
      12'h899: dout  = 8'b00000110; // 2201 :   6 - 0x6
      12'h89A: dout  = 8'b00000110; // 2202 :   6 - 0x6
      12'h89B: dout  = 8'b00000110; // 2203 :   6 - 0x6
      12'h89C: dout  = 8'b11000110; // 2204 : 198 - 0xc6
      12'h89D: dout  = 8'b11000110; // 2205 : 198 - 0xc6
      12'h89E: dout  = 8'b01111100; // 2206 : 124 - 0x7c
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b11000110; // 2208 : 198 - 0xc6 -- Background 0x14
      12'h8A1: dout  = 8'b11001100; // 2209 : 204 - 0xcc
      12'h8A2: dout  = 8'b11011000; // 2210 : 216 - 0xd8
      12'h8A3: dout  = 8'b11110000; // 2211 : 240 - 0xf0
      12'h8A4: dout  = 8'b11111000; // 2212 : 248 - 0xf8
      12'h8A5: dout  = 8'b11011100; // 2213 : 220 - 0xdc
      12'h8A6: dout  = 8'b11001110; // 2214 : 206 - 0xce
      12'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout  = 8'b01100000; // 2216 :  96 - 0x60 -- Background 0x15
      12'h8A9: dout  = 8'b01100000; // 2217 :  96 - 0x60
      12'h8AA: dout  = 8'b01100000; // 2218 :  96 - 0x60
      12'h8AB: dout  = 8'b01100000; // 2219 :  96 - 0x60
      12'h8AC: dout  = 8'b01100000; // 2220 :  96 - 0x60
      12'h8AD: dout  = 8'b01100000; // 2221 :  96 - 0x60
      12'h8AE: dout  = 8'b01111110; // 2222 : 126 - 0x7e
      12'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout  = 8'b11000110; // 2224 : 198 - 0xc6 -- Background 0x16
      12'h8B1: dout  = 8'b11101110; // 2225 : 238 - 0xee
      12'h8B2: dout  = 8'b11111110; // 2226 : 254 - 0xfe
      12'h8B3: dout  = 8'b11111110; // 2227 : 254 - 0xfe
      12'h8B4: dout  = 8'b11010110; // 2228 : 214 - 0xd6
      12'h8B5: dout  = 8'b11000110; // 2229 : 198 - 0xc6
      12'h8B6: dout  = 8'b11000110; // 2230 : 198 - 0xc6
      12'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout  = 8'b11000110; // 2232 : 198 - 0xc6 -- Background 0x17
      12'h8B9: dout  = 8'b11100110; // 2233 : 230 - 0xe6
      12'h8BA: dout  = 8'b11110110; // 2234 : 246 - 0xf6
      12'h8BB: dout  = 8'b11111110; // 2235 : 254 - 0xfe
      12'h8BC: dout  = 8'b11011110; // 2236 : 222 - 0xde
      12'h8BD: dout  = 8'b11001110; // 2237 : 206 - 0xce
      12'h8BE: dout  = 8'b11000110; // 2238 : 198 - 0xc6
      12'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout  = 8'b01111100; // 2240 : 124 - 0x7c -- Background 0x18
      12'h8C1: dout  = 8'b11000110; // 2241 : 198 - 0xc6
      12'h8C2: dout  = 8'b11000110; // 2242 : 198 - 0xc6
      12'h8C3: dout  = 8'b11000110; // 2243 : 198 - 0xc6
      12'h8C4: dout  = 8'b11000110; // 2244 : 198 - 0xc6
      12'h8C5: dout  = 8'b11000110; // 2245 : 198 - 0xc6
      12'h8C6: dout  = 8'b01111100; // 2246 : 124 - 0x7c
      12'h8C7: dout  = 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout  = 8'b11111100; // 2248 : 252 - 0xfc -- Background 0x19
      12'h8C9: dout  = 8'b11000110; // 2249 : 198 - 0xc6
      12'h8CA: dout  = 8'b11000110; // 2250 : 198 - 0xc6
      12'h8CB: dout  = 8'b11000110; // 2251 : 198 - 0xc6
      12'h8CC: dout  = 8'b11111100; // 2252 : 252 - 0xfc
      12'h8CD: dout  = 8'b11000000; // 2253 : 192 - 0xc0
      12'h8CE: dout  = 8'b11000000; // 2254 : 192 - 0xc0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b01111100; // 2256 : 124 - 0x7c -- Background 0x1a
      12'h8D1: dout  = 8'b11000110; // 2257 : 198 - 0xc6
      12'h8D2: dout  = 8'b11000110; // 2258 : 198 - 0xc6
      12'h8D3: dout  = 8'b11000110; // 2259 : 198 - 0xc6
      12'h8D4: dout  = 8'b11011110; // 2260 : 222 - 0xde
      12'h8D5: dout  = 8'b11001100; // 2261 : 204 - 0xcc
      12'h8D6: dout  = 8'b01111010; // 2262 : 122 - 0x7a
      12'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout  = 8'b11111100; // 2264 : 252 - 0xfc -- Background 0x1b
      12'h8D9: dout  = 8'b11000110; // 2265 : 198 - 0xc6
      12'h8DA: dout  = 8'b11000110; // 2266 : 198 - 0xc6
      12'h8DB: dout  = 8'b11001110; // 2267 : 206 - 0xce
      12'h8DC: dout  = 8'b11111000; // 2268 : 248 - 0xf8
      12'h8DD: dout  = 8'b11011100; // 2269 : 220 - 0xdc
      12'h8DE: dout  = 8'b11001110; // 2270 : 206 - 0xce
      12'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout  = 8'b01111000; // 2272 : 120 - 0x78 -- Background 0x1c
      12'h8E1: dout  = 8'b11001100; // 2273 : 204 - 0xcc
      12'h8E2: dout  = 8'b11000000; // 2274 : 192 - 0xc0
      12'h8E3: dout  = 8'b01111100; // 2275 : 124 - 0x7c
      12'h8E4: dout  = 8'b00000110; // 2276 :   6 - 0x6
      12'h8E5: dout  = 8'b11000110; // 2277 : 198 - 0xc6
      12'h8E6: dout  = 8'b01111100; // 2278 : 124 - 0x7c
      12'h8E7: dout  = 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout  = 8'b01111110; // 2280 : 126 - 0x7e -- Background 0x1d
      12'h8E9: dout  = 8'b00011000; // 2281 :  24 - 0x18
      12'h8EA: dout  = 8'b00011000; // 2282 :  24 - 0x18
      12'h8EB: dout  = 8'b00011000; // 2283 :  24 - 0x18
      12'h8EC: dout  = 8'b00011000; // 2284 :  24 - 0x18
      12'h8ED: dout  = 8'b00011000; // 2285 :  24 - 0x18
      12'h8EE: dout  = 8'b00011000; // 2286 :  24 - 0x18
      12'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout  = 8'b11000110; // 2288 : 198 - 0xc6 -- Background 0x1e
      12'h8F1: dout  = 8'b11000110; // 2289 : 198 - 0xc6
      12'h8F2: dout  = 8'b11000110; // 2290 : 198 - 0xc6
      12'h8F3: dout  = 8'b11000110; // 2291 : 198 - 0xc6
      12'h8F4: dout  = 8'b11000110; // 2292 : 198 - 0xc6
      12'h8F5: dout  = 8'b11000110; // 2293 : 198 - 0xc6
      12'h8F6: dout  = 8'b01111100; // 2294 : 124 - 0x7c
      12'h8F7: dout  = 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout  = 8'b11000110; // 2296 : 198 - 0xc6 -- Background 0x1f
      12'h8F9: dout  = 8'b11000110; // 2297 : 198 - 0xc6
      12'h8FA: dout  = 8'b11000110; // 2298 : 198 - 0xc6
      12'h8FB: dout  = 8'b11101110; // 2299 : 238 - 0xee
      12'h8FC: dout  = 8'b01111100; // 2300 : 124 - 0x7c
      12'h8FD: dout  = 8'b00111000; // 2301 :  56 - 0x38
      12'h8FE: dout  = 8'b00010000; // 2302 :  16 - 0x10
      12'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout  = 8'b11000110; // 2304 : 198 - 0xc6 -- Background 0x20
      12'h901: dout  = 8'b11000110; // 2305 : 198 - 0xc6
      12'h902: dout  = 8'b11010110; // 2306 : 214 - 0xd6
      12'h903: dout  = 8'b11111110; // 2307 : 254 - 0xfe
      12'h904: dout  = 8'b11111110; // 2308 : 254 - 0xfe
      12'h905: dout  = 8'b11101110; // 2309 : 238 - 0xee
      12'h906: dout  = 8'b11000110; // 2310 : 198 - 0xc6
      12'h907: dout  = 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout  = 8'b11000110; // 2312 : 198 - 0xc6 -- Background 0x21
      12'h909: dout  = 8'b11101110; // 2313 : 238 - 0xee
      12'h90A: dout  = 8'b01111100; // 2314 : 124 - 0x7c
      12'h90B: dout  = 8'b00111000; // 2315 :  56 - 0x38
      12'h90C: dout  = 8'b01111100; // 2316 : 124 - 0x7c
      12'h90D: dout  = 8'b11101110; // 2317 : 238 - 0xee
      12'h90E: dout  = 8'b11000110; // 2318 : 198 - 0xc6
      12'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout  = 8'b01100110; // 2320 : 102 - 0x66 -- Background 0x22
      12'h911: dout  = 8'b01100110; // 2321 : 102 - 0x66
      12'h912: dout  = 8'b01100110; // 2322 : 102 - 0x66
      12'h913: dout  = 8'b00111100; // 2323 :  60 - 0x3c
      12'h914: dout  = 8'b00011000; // 2324 :  24 - 0x18
      12'h915: dout  = 8'b00011000; // 2325 :  24 - 0x18
      12'h916: dout  = 8'b00011000; // 2326 :  24 - 0x18
      12'h917: dout  = 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout  = 8'b11111110; // 2328 : 254 - 0xfe -- Background 0x23
      12'h919: dout  = 8'b00001110; // 2329 :  14 - 0xe
      12'h91A: dout  = 8'b00011100; // 2330 :  28 - 0x1c
      12'h91B: dout  = 8'b00111000; // 2331 :  56 - 0x38
      12'h91C: dout  = 8'b01110000; // 2332 : 112 - 0x70
      12'h91D: dout  = 8'b11100000; // 2333 : 224 - 0xe0
      12'h91E: dout  = 8'b11111110; // 2334 : 254 - 0xfe
      12'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout  = 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout  = 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout  = 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout  = 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout  = 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout  = 8'b11111111; // 2344 : 255 - 0xff -- Background 0x25
      12'h929: dout  = 8'b11111111; // 2345 : 255 - 0xff
      12'h92A: dout  = 8'b11111111; // 2346 : 255 - 0xff
      12'h92B: dout  = 8'b11111111; // 2347 : 255 - 0xff
      12'h92C: dout  = 8'b11111111; // 2348 : 255 - 0xff
      12'h92D: dout  = 8'b11111111; // 2349 : 255 - 0xff
      12'h92E: dout  = 8'b11111111; // 2350 : 255 - 0xff
      12'h92F: dout  = 8'b11111111; // 2351 : 255 - 0xff
      12'h930: dout  = 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout  = 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout  = 8'b00000000; // 2354 :   0 - 0x0
      12'h933: dout  = 8'b00000000; // 2355 :   0 - 0x0
      12'h934: dout  = 8'b00000000; // 2356 :   0 - 0x0
      12'h935: dout  = 8'b00000000; // 2357 :   0 - 0x0
      12'h936: dout  = 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout  = 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout  = 8'b11111111; // 2360 : 255 - 0xff -- Background 0x27
      12'h939: dout  = 8'b11111111; // 2361 : 255 - 0xff
      12'h93A: dout  = 8'b11111111; // 2362 : 255 - 0xff
      12'h93B: dout  = 8'b11111111; // 2363 : 255 - 0xff
      12'h93C: dout  = 8'b11111111; // 2364 : 255 - 0xff
      12'h93D: dout  = 8'b11111111; // 2365 : 255 - 0xff
      12'h93E: dout  = 8'b11111111; // 2366 : 255 - 0xff
      12'h93F: dout  = 8'b11111111; // 2367 : 255 - 0xff
      12'h940: dout  = 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout  = 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout  = 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout  = 8'b01111110; // 2371 : 126 - 0x7e
      12'h944: dout  = 8'b01111110; // 2372 : 126 - 0x7e
      12'h945: dout  = 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout  = 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout  = 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0 -- Background 0x29
      12'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout  = 8'b01000100; // 2378 :  68 - 0x44
      12'h94B: dout  = 8'b00101000; // 2379 :  40 - 0x28
      12'h94C: dout  = 8'b00010000; // 2380 :  16 - 0x10
      12'h94D: dout  = 8'b00101000; // 2381 :  40 - 0x28
      12'h94E: dout  = 8'b01000100; // 2382 :  68 - 0x44
      12'h94F: dout  = 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout  = 8'b11111111; // 2384 : 255 - 0xff -- Background 0x2a
      12'h951: dout  = 8'b11111111; // 2385 : 255 - 0xff
      12'h952: dout  = 8'b11111111; // 2386 : 255 - 0xff
      12'h953: dout  = 8'b11111111; // 2387 : 255 - 0xff
      12'h954: dout  = 8'b11111111; // 2388 : 255 - 0xff
      12'h955: dout  = 8'b11111111; // 2389 : 255 - 0xff
      12'h956: dout  = 8'b11111111; // 2390 : 255 - 0xff
      12'h957: dout  = 8'b11111111; // 2391 : 255 - 0xff
      12'h958: dout  = 8'b00011000; // 2392 :  24 - 0x18 -- Background 0x2b
      12'h959: dout  = 8'b00111100; // 2393 :  60 - 0x3c
      12'h95A: dout  = 8'b00111100; // 2394 :  60 - 0x3c
      12'h95B: dout  = 8'b00111100; // 2395 :  60 - 0x3c
      12'h95C: dout  = 8'b00011000; // 2396 :  24 - 0x18
      12'h95D: dout  = 8'b00011000; // 2397 :  24 - 0x18
      12'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout  = 8'b00011000; // 2399 :  24 - 0x18
      12'h960: dout  = 8'b11111111; // 2400 : 255 - 0xff -- Background 0x2c
      12'h961: dout  = 8'b01111111; // 2401 : 127 - 0x7f
      12'h962: dout  = 8'b01111111; // 2402 : 127 - 0x7f
      12'h963: dout  = 8'b01111111; // 2403 : 127 - 0x7f
      12'h964: dout  = 8'b01111111; // 2404 : 127 - 0x7f
      12'h965: dout  = 8'b11111111; // 2405 : 255 - 0xff
      12'h966: dout  = 8'b11100011; // 2406 : 227 - 0xe3
      12'h967: dout  = 8'b11000001; // 2407 : 193 - 0xc1
      12'h968: dout  = 8'b10000000; // 2408 : 128 - 0x80 -- Background 0x2d
      12'h969: dout  = 8'b10000000; // 2409 : 128 - 0x80
      12'h96A: dout  = 8'b10000000; // 2410 : 128 - 0x80
      12'h96B: dout  = 8'b11000001; // 2411 : 193 - 0xc1
      12'h96C: dout  = 8'b11100011; // 2412 : 227 - 0xe3
      12'h96D: dout  = 8'b11111111; // 2413 : 255 - 0xff
      12'h96E: dout  = 8'b11111111; // 2414 : 255 - 0xff
      12'h96F: dout  = 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout  = 8'b00111000; // 2416 :  56 - 0x38 -- Background 0x2e
      12'h971: dout  = 8'b01111100; // 2417 : 124 - 0x7c
      12'h972: dout  = 8'b01111100; // 2418 : 124 - 0x7c
      12'h973: dout  = 8'b01111100; // 2419 : 124 - 0x7c
      12'h974: dout  = 8'b01111100; // 2420 : 124 - 0x7c
      12'h975: dout  = 8'b01111100; // 2421 : 124 - 0x7c
      12'h976: dout  = 8'b00111000; // 2422 :  56 - 0x38
      12'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout  = 8'b00000011; // 2424 :   3 - 0x3 -- Background 0x2f
      12'h979: dout  = 8'b00000110; // 2425 :   6 - 0x6
      12'h97A: dout  = 8'b00001100; // 2426 :  12 - 0xc
      12'h97B: dout  = 8'b00001100; // 2427 :  12 - 0xc
      12'h97C: dout  = 8'b00001000; // 2428 :   8 - 0x8
      12'h97D: dout  = 8'b00001000; // 2429 :   8 - 0x8
      12'h97E: dout  = 8'b00000100; // 2430 :   4 - 0x4
      12'h97F: dout  = 8'b00000011; // 2431 :   3 - 0x3
      12'h980: dout  = 8'b00000001; // 2432 :   1 - 0x1 -- Background 0x30
      12'h981: dout  = 8'b00000010; // 2433 :   2 - 0x2
      12'h982: dout  = 8'b00000100; // 2434 :   4 - 0x4
      12'h983: dout  = 8'b00001000; // 2435 :   8 - 0x8
      12'h984: dout  = 8'b00010000; // 2436 :  16 - 0x10
      12'h985: dout  = 8'b00100000; // 2437 :  32 - 0x20
      12'h986: dout  = 8'b01000000; // 2438 :  64 - 0x40
      12'h987: dout  = 8'b10000000; // 2439 : 128 - 0x80
      12'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0 -- Background 0x31
      12'h989: dout  = 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout  = 8'b00000111; // 2445 :   7 - 0x7
      12'h98E: dout  = 8'b00111000; // 2446 :  56 - 0x38
      12'h98F: dout  = 8'b11000000; // 2447 : 192 - 0xc0
      12'h990: dout  = 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x32
      12'h991: dout  = 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout  = 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout  = 8'b00000000; // 2452 :   0 - 0x0
      12'h995: dout  = 8'b11100000; // 2453 : 224 - 0xe0
      12'h996: dout  = 8'b00011100; // 2454 :  28 - 0x1c
      12'h997: dout  = 8'b00000011; // 2455 :   3 - 0x3
      12'h998: dout  = 8'b10000000; // 2456 : 128 - 0x80 -- Background 0x33
      12'h999: dout  = 8'b01000000; // 2457 :  64 - 0x40
      12'h99A: dout  = 8'b00100000; // 2458 :  32 - 0x20
      12'h99B: dout  = 8'b00010000; // 2459 :  16 - 0x10
      12'h99C: dout  = 8'b00001000; // 2460 :   8 - 0x8
      12'h99D: dout  = 8'b00000100; // 2461 :   4 - 0x4
      12'h99E: dout  = 8'b00000010; // 2462 :   2 - 0x2
      12'h99F: dout  = 8'b00000001; // 2463 :   1 - 0x1
      12'h9A0: dout  = 8'b00000100; // 2464 :   4 - 0x4 -- Background 0x34
      12'h9A1: dout  = 8'b00001110; // 2465 :  14 - 0xe
      12'h9A2: dout  = 8'b00001110; // 2466 :  14 - 0xe
      12'h9A3: dout  = 8'b00001110; // 2467 :  14 - 0xe
      12'h9A4: dout  = 8'b01101110; // 2468 : 110 - 0x6e
      12'h9A5: dout  = 8'b01100100; // 2469 : 100 - 0x64
      12'h9A6: dout  = 8'b01100000; // 2470 :  96 - 0x60
      12'h9A7: dout  = 8'b01100000; // 2471 :  96 - 0x60
      12'h9A8: dout  = 8'b00000111; // 2472 :   7 - 0x7 -- Background 0x35
      12'h9A9: dout  = 8'b00001111; // 2473 :  15 - 0xf
      12'h9AA: dout  = 8'b00011111; // 2474 :  31 - 0x1f
      12'h9AB: dout  = 8'b00011111; // 2475 :  31 - 0x1f
      12'h9AC: dout  = 8'b01111111; // 2476 : 127 - 0x7f
      12'h9AD: dout  = 8'b11111111; // 2477 : 255 - 0xff
      12'h9AE: dout  = 8'b11111111; // 2478 : 255 - 0xff
      12'h9AF: dout  = 8'b01111111; // 2479 : 127 - 0x7f
      12'h9B0: dout  = 8'b00000011; // 2480 :   3 - 0x3 -- Background 0x36
      12'h9B1: dout  = 8'b00000111; // 2481 :   7 - 0x7
      12'h9B2: dout  = 8'b00011111; // 2482 :  31 - 0x1f
      12'h9B3: dout  = 8'b00111111; // 2483 :  63 - 0x3f
      12'h9B4: dout  = 8'b00111111; // 2484 :  63 - 0x3f
      12'h9B5: dout  = 8'b00111111; // 2485 :  63 - 0x3f
      12'h9B6: dout  = 8'b01111001; // 2486 : 121 - 0x79
      12'h9B7: dout  = 8'b11110111; // 2487 : 247 - 0xf7
      12'h9B8: dout  = 8'b11000000; // 2488 : 192 - 0xc0 -- Background 0x37
      12'h9B9: dout  = 8'b11100000; // 2489 : 224 - 0xe0
      12'h9BA: dout  = 8'b11110000; // 2490 : 240 - 0xf0
      12'h9BB: dout  = 8'b11110100; // 2491 : 244 - 0xf4
      12'h9BC: dout  = 8'b11111110; // 2492 : 254 - 0xfe
      12'h9BD: dout  = 8'b10111111; // 2493 : 191 - 0xbf
      12'h9BE: dout  = 8'b11011111; // 2494 : 223 - 0xdf
      12'h9BF: dout  = 8'b11111111; // 2495 : 255 - 0xff
      12'h9C0: dout  = 8'b10010000; // 2496 : 144 - 0x90 -- Background 0x38
      12'h9C1: dout  = 8'b10111000; // 2497 : 184 - 0xb8
      12'h9C2: dout  = 8'b11111000; // 2498 : 248 - 0xf8
      12'h9C3: dout  = 8'b11111010; // 2499 : 250 - 0xfa
      12'h9C4: dout  = 8'b11111111; // 2500 : 255 - 0xff
      12'h9C5: dout  = 8'b11111111; // 2501 : 255 - 0xff
      12'h9C6: dout  = 8'b11111111; // 2502 : 255 - 0xff
      12'h9C7: dout  = 8'b11111110; // 2503 : 254 - 0xfe
      12'h9C8: dout  = 8'b00111011; // 2504 :  59 - 0x3b -- Background 0x39
      12'h9C9: dout  = 8'b00011101; // 2505 :  29 - 0x1d
      12'h9CA: dout  = 8'b00001110; // 2506 :  14 - 0xe
      12'h9CB: dout  = 8'b00001111; // 2507 :  15 - 0xf
      12'h9CC: dout  = 8'b00000111; // 2508 :   7 - 0x7
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b11111111; // 2512 : 255 - 0xff -- Background 0x3a
      12'h9D1: dout  = 8'b10111111; // 2513 : 191 - 0xbf
      12'h9D2: dout  = 8'b00011100; // 2514 :  28 - 0x1c
      12'h9D3: dout  = 8'b11000000; // 2515 : 192 - 0xc0
      12'h9D4: dout  = 8'b11110011; // 2516 : 243 - 0xf3
      12'h9D5: dout  = 8'b11111111; // 2517 : 255 - 0xff
      12'h9D6: dout  = 8'b01111110; // 2518 : 126 - 0x7e
      12'h9D7: dout  = 8'b00011100; // 2519 :  28 - 0x1c
      12'h9D8: dout  = 8'b10111111; // 2520 : 191 - 0xbf -- Background 0x3b
      12'h9D9: dout  = 8'b01111111; // 2521 : 127 - 0x7f
      12'h9DA: dout  = 8'b00111101; // 2522 :  61 - 0x3d
      12'h9DB: dout  = 8'b10000011; // 2523 : 131 - 0x83
      12'h9DC: dout  = 8'b11000111; // 2524 : 199 - 0xc7
      12'h9DD: dout  = 8'b11111111; // 2525 : 255 - 0xff
      12'h9DE: dout  = 8'b11111111; // 2526 : 255 - 0xff
      12'h9DF: dout  = 8'b00111100; // 2527 :  60 - 0x3c
      12'h9E0: dout  = 8'b11111100; // 2528 : 252 - 0xfc -- Background 0x3c
      12'h9E1: dout  = 8'b11111110; // 2529 : 254 - 0xfe
      12'h9E2: dout  = 8'b11111111; // 2530 : 255 - 0xff
      12'h9E3: dout  = 8'b11111110; // 2531 : 254 - 0xfe
      12'h9E4: dout  = 8'b11111110; // 2532 : 254 - 0xfe
      12'h9E5: dout  = 8'b11111000; // 2533 : 248 - 0xf8
      12'h9E6: dout  = 8'b01100000; // 2534 :  96 - 0x60
      12'h9E7: dout  = 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout  = 8'b11000000; // 2536 : 192 - 0xc0 -- Background 0x3d
      12'h9E9: dout  = 8'b00100000; // 2537 :  32 - 0x20
      12'h9EA: dout  = 8'b00010000; // 2538 :  16 - 0x10
      12'h9EB: dout  = 8'b00010000; // 2539 :  16 - 0x10
      12'h9EC: dout  = 8'b00010000; // 2540 :  16 - 0x10
      12'h9ED: dout  = 8'b00010000; // 2541 :  16 - 0x10
      12'h9EE: dout  = 8'b00100000; // 2542 :  32 - 0x20
      12'h9EF: dout  = 8'b11000000; // 2543 : 192 - 0xc0
      12'h9F0: dout  = 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout  = 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout  = 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout  = 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout  = 8'b00111111; // 2548 :  63 - 0x3f
      12'h9F5: dout  = 8'b01111111; // 2549 : 127 - 0x7f
      12'h9F6: dout  = 8'b11100000; // 2550 : 224 - 0xe0
      12'h9F7: dout  = 8'b11000000; // 2551 : 192 - 0xc0
      12'h9F8: dout  = 8'b10001000; // 2552 : 136 - 0x88 -- Background 0x3f
      12'h9F9: dout  = 8'b10011100; // 2553 : 156 - 0x9c
      12'h9FA: dout  = 8'b10001000; // 2554 : 136 - 0x88
      12'h9FB: dout  = 8'b10000000; // 2555 : 128 - 0x80
      12'h9FC: dout  = 8'b10000000; // 2556 : 128 - 0x80
      12'h9FD: dout  = 8'b10000000; // 2557 : 128 - 0x80
      12'h9FE: dout  = 8'b10000000; // 2558 : 128 - 0x80
      12'h9FF: dout  = 8'b10000000; // 2559 : 128 - 0x80
      12'hA00: dout  = 8'b11111110; // 2560 : 254 - 0xfe -- Background 0x40
      12'hA01: dout  = 8'b11111110; // 2561 : 254 - 0xfe
      12'hA02: dout  = 8'b11111110; // 2562 : 254 - 0xfe
      12'hA03: dout  = 8'b11111110; // 2563 : 254 - 0xfe
      12'hA04: dout  = 8'b11111110; // 2564 : 254 - 0xfe
      12'hA05: dout  = 8'b11111110; // 2565 : 254 - 0xfe
      12'hA06: dout  = 8'b11111110; // 2566 : 254 - 0xfe
      12'hA07: dout  = 8'b11111110; // 2567 : 254 - 0xfe
      12'hA08: dout  = 8'b00001000; // 2568 :   8 - 0x8 -- Background 0x41
      12'hA09: dout  = 8'b00010100; // 2569 :  20 - 0x14
      12'hA0A: dout  = 8'b00100100; // 2570 :  36 - 0x24
      12'hA0B: dout  = 8'b11000100; // 2571 : 196 - 0xc4
      12'hA0C: dout  = 8'b00000011; // 2572 :   3 - 0x3
      12'hA0D: dout  = 8'b01000000; // 2573 :  64 - 0x40
      12'hA0E: dout  = 8'b10100001; // 2574 : 161 - 0xa1
      12'hA0F: dout  = 8'b00100110; // 2575 :  38 - 0x26
      12'hA10: dout  = 8'b11111111; // 2576 : 255 - 0xff -- Background 0x42
      12'hA11: dout  = 8'b11111111; // 2577 : 255 - 0xff
      12'hA12: dout  = 8'b11111111; // 2578 : 255 - 0xff
      12'hA13: dout  = 8'b11111111; // 2579 : 255 - 0xff
      12'hA14: dout  = 8'b01111111; // 2580 : 127 - 0x7f
      12'hA15: dout  = 8'b01111111; // 2581 : 127 - 0x7f
      12'hA16: dout  = 8'b01111111; // 2582 : 127 - 0x7f
      12'hA17: dout  = 8'b01111111; // 2583 : 127 - 0x7f
      12'hA18: dout  = 8'b11111111; // 2584 : 255 - 0xff -- Background 0x43
      12'hA19: dout  = 8'b11111111; // 2585 : 255 - 0xff
      12'hA1A: dout  = 8'b11111111; // 2586 : 255 - 0xff
      12'hA1B: dout  = 8'b11111111; // 2587 : 255 - 0xff
      12'hA1C: dout  = 8'b11111111; // 2588 : 255 - 0xff
      12'hA1D: dout  = 8'b11111111; // 2589 : 255 - 0xff
      12'hA1E: dout  = 8'b11111111; // 2590 : 255 - 0xff
      12'hA1F: dout  = 8'b11111111; // 2591 : 255 - 0xff
      12'hA20: dout  = 8'b01111111; // 2592 : 127 - 0x7f -- Background 0x44
      12'hA21: dout  = 8'b10000000; // 2593 : 128 - 0x80
      12'hA22: dout  = 8'b10000000; // 2594 : 128 - 0x80
      12'hA23: dout  = 8'b10011000; // 2595 : 152 - 0x98
      12'hA24: dout  = 8'b10011100; // 2596 : 156 - 0x9c
      12'hA25: dout  = 8'b10001100; // 2597 : 140 - 0x8c
      12'hA26: dout  = 8'b10000000; // 2598 : 128 - 0x80
      12'hA27: dout  = 8'b10000000; // 2599 : 128 - 0x80
      12'hA28: dout  = 8'b11111111; // 2600 : 255 - 0xff -- Background 0x45
      12'hA29: dout  = 8'b00000001; // 2601 :   1 - 0x1
      12'hA2A: dout  = 8'b00000001; // 2602 :   1 - 0x1
      12'hA2B: dout  = 8'b11111111; // 2603 : 255 - 0xff
      12'hA2C: dout  = 8'b00010000; // 2604 :  16 - 0x10
      12'hA2D: dout  = 8'b00010000; // 2605 :  16 - 0x10
      12'hA2E: dout  = 8'b00010000; // 2606 :  16 - 0x10
      12'hA2F: dout  = 8'b11111111; // 2607 : 255 - 0xff
      12'hA30: dout  = 8'b10000000; // 2608 : 128 - 0x80 -- Background 0x46
      12'hA31: dout  = 8'b10000000; // 2609 : 128 - 0x80
      12'hA32: dout  = 8'b10000000; // 2610 : 128 - 0x80
      12'hA33: dout  = 8'b10000000; // 2611 : 128 - 0x80
      12'hA34: dout  = 8'b10000000; // 2612 : 128 - 0x80
      12'hA35: dout  = 8'b10000000; // 2613 : 128 - 0x80
      12'hA36: dout  = 8'b10000000; // 2614 : 128 - 0x80
      12'hA37: dout  = 8'b10000000; // 2615 : 128 - 0x80
      12'hA38: dout  = 8'b00000001; // 2616 :   1 - 0x1 -- Background 0x47
      12'hA39: dout  = 8'b00000001; // 2617 :   1 - 0x1
      12'hA3A: dout  = 8'b00000001; // 2618 :   1 - 0x1
      12'hA3B: dout  = 8'b11111111; // 2619 : 255 - 0xff
      12'hA3C: dout  = 8'b00010000; // 2620 :  16 - 0x10
      12'hA3D: dout  = 8'b00010000; // 2621 :  16 - 0x10
      12'hA3E: dout  = 8'b00010000; // 2622 :  16 - 0x10
      12'hA3F: dout  = 8'b11111111; // 2623 : 255 - 0xff
      12'hA40: dout  = 8'b11111111; // 2624 : 255 - 0xff -- Background 0x48
      12'hA41: dout  = 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout  = 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout  = 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout  = 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout  = 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout  = 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout  = 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout  = 8'b11111110; // 2632 : 254 - 0xfe -- Background 0x49
      12'hA49: dout  = 8'b00000001; // 2633 :   1 - 0x1
      12'hA4A: dout  = 8'b00000001; // 2634 :   1 - 0x1
      12'hA4B: dout  = 8'b00011001; // 2635 :  25 - 0x19
      12'hA4C: dout  = 8'b00011101; // 2636 :  29 - 0x1d
      12'hA4D: dout  = 8'b00001101; // 2637 :  13 - 0xd
      12'hA4E: dout  = 8'b00000001; // 2638 :   1 - 0x1
      12'hA4F: dout  = 8'b00000001; // 2639 :   1 - 0x1
      12'hA50: dout  = 8'b00000001; // 2640 :   1 - 0x1 -- Background 0x4a
      12'hA51: dout  = 8'b00000001; // 2641 :   1 - 0x1
      12'hA52: dout  = 8'b00000001; // 2642 :   1 - 0x1
      12'hA53: dout  = 8'b00000001; // 2643 :   1 - 0x1
      12'hA54: dout  = 8'b00000001; // 2644 :   1 - 0x1
      12'hA55: dout  = 8'b00000001; // 2645 :   1 - 0x1
      12'hA56: dout  = 8'b00000001; // 2646 :   1 - 0x1
      12'hA57: dout  = 8'b00000001; // 2647 :   1 - 0x1
      12'hA58: dout  = 8'b00111111; // 2648 :  63 - 0x3f -- Background 0x4b
      12'hA59: dout  = 8'b01111111; // 2649 : 127 - 0x7f
      12'hA5A: dout  = 8'b01111111; // 2650 : 127 - 0x7f
      12'hA5B: dout  = 8'b11111111; // 2651 : 255 - 0xff
      12'hA5C: dout  = 8'b11111111; // 2652 : 255 - 0xff
      12'hA5D: dout  = 8'b11111111; // 2653 : 255 - 0xff
      12'hA5E: dout  = 8'b11111111; // 2654 : 255 - 0xff
      12'hA5F: dout  = 8'b11111111; // 2655 : 255 - 0xff
      12'hA60: dout  = 8'b11111111; // 2656 : 255 - 0xff -- Background 0x4c
      12'hA61: dout  = 8'b11111111; // 2657 : 255 - 0xff
      12'hA62: dout  = 8'b11111111; // 2658 : 255 - 0xff
      12'hA63: dout  = 8'b11111111; // 2659 : 255 - 0xff
      12'hA64: dout  = 8'b11111111; // 2660 : 255 - 0xff
      12'hA65: dout  = 8'b11111111; // 2661 : 255 - 0xff
      12'hA66: dout  = 8'b01111110; // 2662 : 126 - 0x7e
      12'hA67: dout  = 8'b00111100; // 2663 :  60 - 0x3c
      12'hA68: dout  = 8'b11111111; // 2664 : 255 - 0xff -- Background 0x4d
      12'hA69: dout  = 8'b11111111; // 2665 : 255 - 0xff
      12'hA6A: dout  = 8'b11111111; // 2666 : 255 - 0xff
      12'hA6B: dout  = 8'b11111111; // 2667 : 255 - 0xff
      12'hA6C: dout  = 8'b11111111; // 2668 : 255 - 0xff
      12'hA6D: dout  = 8'b11111111; // 2669 : 255 - 0xff
      12'hA6E: dout  = 8'b11111111; // 2670 : 255 - 0xff
      12'hA6F: dout  = 8'b11111111; // 2671 : 255 - 0xff
      12'hA70: dout  = 8'b11111111; // 2672 : 255 - 0xff -- Background 0x4e
      12'hA71: dout  = 8'b11111111; // 2673 : 255 - 0xff
      12'hA72: dout  = 8'b11111111; // 2674 : 255 - 0xff
      12'hA73: dout  = 8'b11111111; // 2675 : 255 - 0xff
      12'hA74: dout  = 8'b11111111; // 2676 : 255 - 0xff
      12'hA75: dout  = 8'b11111111; // 2677 : 255 - 0xff
      12'hA76: dout  = 8'b11111110; // 2678 : 254 - 0xfe
      12'hA77: dout  = 8'b01111100; // 2679 : 124 - 0x7c
      12'hA78: dout  = 8'b11111111; // 2680 : 255 - 0xff -- Background 0x4f
      12'hA79: dout  = 8'b11111111; // 2681 : 255 - 0xff
      12'hA7A: dout  = 8'b11111111; // 2682 : 255 - 0xff
      12'hA7B: dout  = 8'b11111111; // 2683 : 255 - 0xff
      12'hA7C: dout  = 8'b11111111; // 2684 : 255 - 0xff
      12'hA7D: dout  = 8'b11111111; // 2685 : 255 - 0xff
      12'hA7E: dout  = 8'b11111110; // 2686 : 254 - 0xfe
      12'hA7F: dout  = 8'b01111100; // 2687 : 124 - 0x7c
      12'hA80: dout  = 8'b11111000; // 2688 : 248 - 0xf8 -- Background 0x50
      12'hA81: dout  = 8'b11111100; // 2689 : 252 - 0xfc
      12'hA82: dout  = 8'b11111110; // 2690 : 254 - 0xfe
      12'hA83: dout  = 8'b11111110; // 2691 : 254 - 0xfe
      12'hA84: dout  = 8'b11111111; // 2692 : 255 - 0xff
      12'hA85: dout  = 8'b11111111; // 2693 : 255 - 0xff
      12'hA86: dout  = 8'b11111111; // 2694 : 255 - 0xff
      12'hA87: dout  = 8'b11111111; // 2695 : 255 - 0xff
      12'hA88: dout  = 8'b11111111; // 2696 : 255 - 0xff -- Background 0x51
      12'hA89: dout  = 8'b11111111; // 2697 : 255 - 0xff
      12'hA8A: dout  = 8'b11111111; // 2698 : 255 - 0xff
      12'hA8B: dout  = 8'b11111111; // 2699 : 255 - 0xff
      12'hA8C: dout  = 8'b11111111; // 2700 : 255 - 0xff
      12'hA8D: dout  = 8'b11111111; // 2701 : 255 - 0xff
      12'hA8E: dout  = 8'b01111110; // 2702 : 126 - 0x7e
      12'hA8F: dout  = 8'b00111100; // 2703 :  60 - 0x3c
      12'hA90: dout  = 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout  = 8'b00001000; // 2705 :   8 - 0x8
      12'hA92: dout  = 8'b00001000; // 2706 :   8 - 0x8
      12'hA93: dout  = 8'b00001000; // 2707 :   8 - 0x8
      12'hA94: dout  = 8'b00010000; // 2708 :  16 - 0x10
      12'hA95: dout  = 8'b00010000; // 2709 :  16 - 0x10
      12'hA96: dout  = 8'b00010000; // 2710 :  16 - 0x10
      12'hA97: dout  = 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout  = 8'b01111111; // 2713 : 127 - 0x7f
      12'hA9A: dout  = 8'b01111111; // 2714 : 127 - 0x7f
      12'hA9B: dout  = 8'b01111000; // 2715 : 120 - 0x78
      12'hA9C: dout  = 8'b01110011; // 2716 : 115 - 0x73
      12'hA9D: dout  = 8'b01110011; // 2717 : 115 - 0x73
      12'hA9E: dout  = 8'b01110011; // 2718 : 115 - 0x73
      12'hA9F: dout  = 8'b01111111; // 2719 : 127 - 0x7f
      12'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout  = 8'b11111111; // 2721 : 255 - 0xff
      12'hAA2: dout  = 8'b11111111; // 2722 : 255 - 0xff
      12'hAA3: dout  = 8'b00111111; // 2723 :  63 - 0x3f
      12'hAA4: dout  = 8'b10011111; // 2724 : 159 - 0x9f
      12'hAA5: dout  = 8'b10011111; // 2725 : 159 - 0x9f
      12'hAA6: dout  = 8'b10011111; // 2726 : 159 - 0x9f
      12'hAA7: dout  = 8'b00011111; // 2727 :  31 - 0x1f
      12'hAA8: dout  = 8'b01111110; // 2728 : 126 - 0x7e -- Background 0x55
      12'hAA9: dout  = 8'b01111110; // 2729 : 126 - 0x7e
      12'hAAA: dout  = 8'b01111111; // 2730 : 127 - 0x7f
      12'hAAB: dout  = 8'b01111110; // 2731 : 126 - 0x7e
      12'hAAC: dout  = 8'b01111110; // 2732 : 126 - 0x7e
      12'hAAD: dout  = 8'b01111111; // 2733 : 127 - 0x7f
      12'hAAE: dout  = 8'b01111111; // 2734 : 127 - 0x7f
      12'hAAF: dout  = 8'b11111111; // 2735 : 255 - 0xff
      12'hAB0: dout  = 8'b01111111; // 2736 : 127 - 0x7f -- Background 0x56
      12'hAB1: dout  = 8'b01111111; // 2737 : 127 - 0x7f
      12'hAB2: dout  = 8'b11111111; // 2738 : 255 - 0xff
      12'hAB3: dout  = 8'b01111111; // 2739 : 127 - 0x7f
      12'hAB4: dout  = 8'b01111111; // 2740 : 127 - 0x7f
      12'hAB5: dout  = 8'b11111111; // 2741 : 255 - 0xff
      12'hAB6: dout  = 8'b11111111; // 2742 : 255 - 0xff
      12'hAB7: dout  = 8'b11111111; // 2743 : 255 - 0xff
      12'hAB8: dout  = 8'b01111111; // 2744 : 127 - 0x7f -- Background 0x57
      12'hAB9: dout  = 8'b10000000; // 2745 : 128 - 0x80
      12'hABA: dout  = 8'b10100000; // 2746 : 160 - 0xa0
      12'hABB: dout  = 8'b10000000; // 2747 : 128 - 0x80
      12'hABC: dout  = 8'b10000000; // 2748 : 128 - 0x80
      12'hABD: dout  = 8'b10000000; // 2749 : 128 - 0x80
      12'hABE: dout  = 8'b10000000; // 2750 : 128 - 0x80
      12'hABF: dout  = 8'b10000000; // 2751 : 128 - 0x80
      12'hAC0: dout  = 8'b11111110; // 2752 : 254 - 0xfe -- Background 0x58
      12'hAC1: dout  = 8'b00000001; // 2753 :   1 - 0x1
      12'hAC2: dout  = 8'b00000101; // 2754 :   5 - 0x5
      12'hAC3: dout  = 8'b00000001; // 2755 :   1 - 0x1
      12'hAC4: dout  = 8'b00000001; // 2756 :   1 - 0x1
      12'hAC5: dout  = 8'b00000001; // 2757 :   1 - 0x1
      12'hAC6: dout  = 8'b00000001; // 2758 :   1 - 0x1
      12'hAC7: dout  = 8'b00000001; // 2759 :   1 - 0x1
      12'hAC8: dout  = 8'b10000000; // 2760 : 128 - 0x80 -- Background 0x59
      12'hAC9: dout  = 8'b10000000; // 2761 : 128 - 0x80
      12'hACA: dout  = 8'b10000000; // 2762 : 128 - 0x80
      12'hACB: dout  = 8'b10000000; // 2763 : 128 - 0x80
      12'hACC: dout  = 8'b10000000; // 2764 : 128 - 0x80
      12'hACD: dout  = 8'b10100000; // 2765 : 160 - 0xa0
      12'hACE: dout  = 8'b10000000; // 2766 : 128 - 0x80
      12'hACF: dout  = 8'b01111111; // 2767 : 127 - 0x7f
      12'hAD0: dout  = 8'b00000001; // 2768 :   1 - 0x1 -- Background 0x5a
      12'hAD1: dout  = 8'b00000001; // 2769 :   1 - 0x1
      12'hAD2: dout  = 8'b00000001; // 2770 :   1 - 0x1
      12'hAD3: dout  = 8'b00000001; // 2771 :   1 - 0x1
      12'hAD4: dout  = 8'b00000001; // 2772 :   1 - 0x1
      12'hAD5: dout  = 8'b00000101; // 2773 :   5 - 0x5
      12'hAD6: dout  = 8'b00000001; // 2774 :   1 - 0x1
      12'hAD7: dout  = 8'b11111110; // 2775 : 254 - 0xfe
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout  = 8'b11111100; // 2780 : 252 - 0xfc
      12'hADD: dout  = 8'b11111110; // 2781 : 254 - 0xfe
      12'hADE: dout  = 8'b00000111; // 2782 :   7 - 0x7
      12'hADF: dout  = 8'b00000011; // 2783 :   3 - 0x3
      12'hAE0: dout  = 8'b00010001; // 2784 :  17 - 0x11 -- Background 0x5c
      12'hAE1: dout  = 8'b00111001; // 2785 :  57 - 0x39
      12'hAE2: dout  = 8'b00010001; // 2786 :  17 - 0x11
      12'hAE3: dout  = 8'b00000001; // 2787 :   1 - 0x1
      12'hAE4: dout  = 8'b00000001; // 2788 :   1 - 0x1
      12'hAE5: dout  = 8'b00000001; // 2789 :   1 - 0x1
      12'hAE6: dout  = 8'b00000001; // 2790 :   1 - 0x1
      12'hAE7: dout  = 8'b00000001; // 2791 :   1 - 0x1
      12'hAE8: dout  = 8'b11101111; // 2792 : 239 - 0xef -- Background 0x5d
      12'hAE9: dout  = 8'b00101000; // 2793 :  40 - 0x28
      12'hAEA: dout  = 8'b00101000; // 2794 :  40 - 0x28
      12'hAEB: dout  = 8'b00101000; // 2795 :  40 - 0x28
      12'hAEC: dout  = 8'b00101000; // 2796 :  40 - 0x28
      12'hAED: dout  = 8'b00101000; // 2797 :  40 - 0x28
      12'hAEE: dout  = 8'b11101111; // 2798 : 239 - 0xef
      12'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout  = 8'b11111110; // 2800 : 254 - 0xfe -- Background 0x5e
      12'hAF1: dout  = 8'b10000010; // 2801 : 130 - 0x82
      12'hAF2: dout  = 8'b10000010; // 2802 : 130 - 0x82
      12'hAF3: dout  = 8'b10000010; // 2803 : 130 - 0x82
      12'hAF4: dout  = 8'b10000010; // 2804 : 130 - 0x82
      12'hAF5: dout  = 8'b10000010; // 2805 : 130 - 0x82
      12'hAF6: dout  = 8'b11111110; // 2806 : 254 - 0xfe
      12'hAF7: dout  = 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout  = 8'b10000000; // 2808 : 128 - 0x80 -- Background 0x5f
      12'hAF9: dout  = 8'b10000000; // 2809 : 128 - 0x80
      12'hAFA: dout  = 8'b10000000; // 2810 : 128 - 0x80
      12'hAFB: dout  = 8'b10011000; // 2811 : 152 - 0x98
      12'hAFC: dout  = 8'b10011100; // 2812 : 156 - 0x9c
      12'hAFD: dout  = 8'b10001100; // 2813 : 140 - 0x8c
      12'hAFE: dout  = 8'b10000000; // 2814 : 128 - 0x80
      12'hAFF: dout  = 8'b01111111; // 2815 : 127 - 0x7f
      12'hB00: dout  = 8'b11111111; // 2816 : 255 - 0xff -- Background 0x60
      12'hB01: dout  = 8'b11111111; // 2817 : 255 - 0xff
      12'hB02: dout  = 8'b10000011; // 2818 : 131 - 0x83
      12'hB03: dout  = 8'b11110011; // 2819 : 243 - 0xf3
      12'hB04: dout  = 8'b11110011; // 2820 : 243 - 0xf3
      12'hB05: dout  = 8'b11110011; // 2821 : 243 - 0xf3
      12'hB06: dout  = 8'b11110011; // 2822 : 243 - 0xf3
      12'hB07: dout  = 8'b11110011; // 2823 : 243 - 0xf3
      12'hB08: dout  = 8'b11111111; // 2824 : 255 - 0xff -- Background 0x61
      12'hB09: dout  = 8'b11111111; // 2825 : 255 - 0xff
      12'hB0A: dout  = 8'b11110000; // 2826 : 240 - 0xf0
      12'hB0B: dout  = 8'b11110110; // 2827 : 246 - 0xf6
      12'hB0C: dout  = 8'b11110110; // 2828 : 246 - 0xf6
      12'hB0D: dout  = 8'b11110110; // 2829 : 246 - 0xf6
      12'hB0E: dout  = 8'b11110110; // 2830 : 246 - 0xf6
      12'hB0F: dout  = 8'b11110110; // 2831 : 246 - 0xf6
      12'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Background 0x62
      12'hB11: dout  = 8'b11111111; // 2833 : 255 - 0xff
      12'hB12: dout  = 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout  = 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout  = 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout  = 8'b00000000; // 2837 :   0 - 0x0
      12'hB16: dout  = 8'b00000000; // 2838 :   0 - 0x0
      12'hB17: dout  = 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout  = 8'b11111111; // 2840 : 255 - 0xff -- Background 0x63
      12'hB19: dout  = 8'b11111111; // 2841 : 255 - 0xff
      12'hB1A: dout  = 8'b00000001; // 2842 :   1 - 0x1
      12'hB1B: dout  = 8'b01010111; // 2843 :  87 - 0x57
      12'hB1C: dout  = 8'b00101111; // 2844 :  47 - 0x2f
      12'hB1D: dout  = 8'b01010111; // 2845 :  87 - 0x57
      12'hB1E: dout  = 8'b00101111; // 2846 :  47 - 0x2f
      12'hB1F: dout  = 8'b01010111; // 2847 :  87 - 0x57
      12'hB20: dout  = 8'b11110011; // 2848 : 243 - 0xf3 -- Background 0x64
      12'hB21: dout  = 8'b11110011; // 2849 : 243 - 0xf3
      12'hB22: dout  = 8'b11110011; // 2850 : 243 - 0xf3
      12'hB23: dout  = 8'b11110011; // 2851 : 243 - 0xf3
      12'hB24: dout  = 8'b11110011; // 2852 : 243 - 0xf3
      12'hB25: dout  = 8'b11110011; // 2853 : 243 - 0xf3
      12'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      12'hB27: dout  = 8'b00111111; // 2855 :  63 - 0x3f
      12'hB28: dout  = 8'b11110110; // 2856 : 246 - 0xf6 -- Background 0x65
      12'hB29: dout  = 8'b11110110; // 2857 : 246 - 0xf6
      12'hB2A: dout  = 8'b11110110; // 2858 : 246 - 0xf6
      12'hB2B: dout  = 8'b11110110; // 2859 : 246 - 0xf6
      12'hB2C: dout  = 8'b11110110; // 2860 : 246 - 0xf6
      12'hB2D: dout  = 8'b11110110; // 2861 : 246 - 0xf6
      12'hB2E: dout  = 8'b11111111; // 2862 : 255 - 0xff
      12'hB2F: dout  = 8'b11111111; // 2863 : 255 - 0xff
      12'hB30: dout  = 8'b00000000; // 2864 :   0 - 0x0 -- Background 0x66
      12'hB31: dout  = 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout  = 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout  = 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout  = 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout  = 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout  = 8'b11111111; // 2870 : 255 - 0xff
      12'hB37: dout  = 8'b11111111; // 2871 : 255 - 0xff
      12'hB38: dout  = 8'b00101111; // 2872 :  47 - 0x2f -- Background 0x67
      12'hB39: dout  = 8'b01010111; // 2873 :  87 - 0x57
      12'hB3A: dout  = 8'b00101111; // 2874 :  47 - 0x2f
      12'hB3B: dout  = 8'b01010111; // 2875 :  87 - 0x57
      12'hB3C: dout  = 8'b00101111; // 2876 :  47 - 0x2f
      12'hB3D: dout  = 8'b01010111; // 2877 :  87 - 0x57
      12'hB3E: dout  = 8'b11111111; // 2878 : 255 - 0xff
      12'hB3F: dout  = 8'b11111100; // 2879 : 252 - 0xfc
      12'hB40: dout  = 8'b00111100; // 2880 :  60 - 0x3c -- Background 0x68
      12'hB41: dout  = 8'b00111100; // 2881 :  60 - 0x3c
      12'hB42: dout  = 8'b00111100; // 2882 :  60 - 0x3c
      12'hB43: dout  = 8'b00111100; // 2883 :  60 - 0x3c
      12'hB44: dout  = 8'b00111100; // 2884 :  60 - 0x3c
      12'hB45: dout  = 8'b00111100; // 2885 :  60 - 0x3c
      12'hB46: dout  = 8'b00111100; // 2886 :  60 - 0x3c
      12'hB47: dout  = 8'b00111100; // 2887 :  60 - 0x3c
      12'hB48: dout  = 8'b11111011; // 2888 : 251 - 0xfb -- Background 0x69
      12'hB49: dout  = 8'b11111011; // 2889 : 251 - 0xfb
      12'hB4A: dout  = 8'b11111011; // 2890 : 251 - 0xfb
      12'hB4B: dout  = 8'b11111011; // 2891 : 251 - 0xfb
      12'hB4C: dout  = 8'b11111011; // 2892 : 251 - 0xfb
      12'hB4D: dout  = 8'b11111011; // 2893 : 251 - 0xfb
      12'hB4E: dout  = 8'b11111011; // 2894 : 251 - 0xfb
      12'hB4F: dout  = 8'b11111011; // 2895 : 251 - 0xfb
      12'hB50: dout  = 8'b10111100; // 2896 : 188 - 0xbc -- Background 0x6a
      12'hB51: dout  = 8'b01011100; // 2897 :  92 - 0x5c
      12'hB52: dout  = 8'b10111100; // 2898 : 188 - 0xbc
      12'hB53: dout  = 8'b01011100; // 2899 :  92 - 0x5c
      12'hB54: dout  = 8'b10111100; // 2900 : 188 - 0xbc
      12'hB55: dout  = 8'b01011100; // 2901 :  92 - 0x5c
      12'hB56: dout  = 8'b10111100; // 2902 : 188 - 0xbc
      12'hB57: dout  = 8'b01011100; // 2903 :  92 - 0x5c
      12'hB58: dout  = 8'b00011111; // 2904 :  31 - 0x1f -- Background 0x6b
      12'hB59: dout  = 8'b00100000; // 2905 :  32 - 0x20
      12'hB5A: dout  = 8'b01000000; // 2906 :  64 - 0x40
      12'hB5B: dout  = 8'b01000000; // 2907 :  64 - 0x40
      12'hB5C: dout  = 8'b10000000; // 2908 : 128 - 0x80
      12'hB5D: dout  = 8'b10000000; // 2909 : 128 - 0x80
      12'hB5E: dout  = 8'b10000000; // 2910 : 128 - 0x80
      12'hB5F: dout  = 8'b10000001; // 2911 : 129 - 0x81
      12'hB60: dout  = 8'b11111111; // 2912 : 255 - 0xff -- Background 0x6c
      12'hB61: dout  = 8'b10000000; // 2913 : 128 - 0x80
      12'hB62: dout  = 8'b10000000; // 2914 : 128 - 0x80
      12'hB63: dout  = 8'b11000000; // 2915 : 192 - 0xc0
      12'hB64: dout  = 8'b11111111; // 2916 : 255 - 0xff
      12'hB65: dout  = 8'b11111111; // 2917 : 255 - 0xff
      12'hB66: dout  = 8'b11111110; // 2918 : 254 - 0xfe
      12'hB67: dout  = 8'b11111110; // 2919 : 254 - 0xfe
      12'hB68: dout  = 8'b11111111; // 2920 : 255 - 0xff -- Background 0x6d
      12'hB69: dout  = 8'b01111111; // 2921 : 127 - 0x7f
      12'hB6A: dout  = 8'b01111111; // 2922 : 127 - 0x7f
      12'hB6B: dout  = 8'b11111111; // 2923 : 255 - 0xff
      12'hB6C: dout  = 8'b11111111; // 2924 : 255 - 0xff
      12'hB6D: dout  = 8'b00000111; // 2925 :   7 - 0x7
      12'hB6E: dout  = 8'b00000011; // 2926 :   3 - 0x3
      12'hB6F: dout  = 8'b00000011; // 2927 :   3 - 0x3
      12'hB70: dout  = 8'b11111111; // 2928 : 255 - 0xff -- Background 0x6e
      12'hB71: dout  = 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout  = 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout  = 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout  = 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout  = 8'b10000001; // 2933 : 129 - 0x81
      12'hB76: dout  = 8'b11000011; // 2934 : 195 - 0xc3
      12'hB77: dout  = 8'b11111111; // 2935 : 255 - 0xff
      12'hB78: dout  = 8'b11111000; // 2936 : 248 - 0xf8 -- Background 0x6f
      12'hB79: dout  = 8'b11111100; // 2937 : 252 - 0xfc
      12'hB7A: dout  = 8'b11111110; // 2938 : 254 - 0xfe
      12'hB7B: dout  = 8'b11111110; // 2939 : 254 - 0xfe
      12'hB7C: dout  = 8'b11100011; // 2940 : 227 - 0xe3
      12'hB7D: dout  = 8'b11000001; // 2941 : 193 - 0xc1
      12'hB7E: dout  = 8'b10000001; // 2942 : 129 - 0x81
      12'hB7F: dout  = 8'b10000001; // 2943 : 129 - 0x81
      12'hB80: dout  = 8'b10000011; // 2944 : 131 - 0x83 -- Background 0x70
      12'hB81: dout  = 8'b11111111; // 2945 : 255 - 0xff
      12'hB82: dout  = 8'b11111111; // 2946 : 255 - 0xff
      12'hB83: dout  = 8'b11111111; // 2947 : 255 - 0xff
      12'hB84: dout  = 8'b11111111; // 2948 : 255 - 0xff
      12'hB85: dout  = 8'b11111111; // 2949 : 255 - 0xff
      12'hB86: dout  = 8'b01111111; // 2950 : 127 - 0x7f
      12'hB87: dout  = 8'b00011111; // 2951 :  31 - 0x1f
      12'hB88: dout  = 8'b11111100; // 2952 : 252 - 0xfc -- Background 0x71
      12'hB89: dout  = 8'b11111100; // 2953 : 252 - 0xfc
      12'hB8A: dout  = 8'b11111100; // 2954 : 252 - 0xfc
      12'hB8B: dout  = 8'b11111100; // 2955 : 252 - 0xfc
      12'hB8C: dout  = 8'b11111110; // 2956 : 254 - 0xfe
      12'hB8D: dout  = 8'b11111110; // 2957 : 254 - 0xfe
      12'hB8E: dout  = 8'b11111111; // 2958 : 255 - 0xff
      12'hB8F: dout  = 8'b11111111; // 2959 : 255 - 0xff
      12'hB90: dout  = 8'b00000001; // 2960 :   1 - 0x1 -- Background 0x72
      12'hB91: dout  = 8'b00000001; // 2961 :   1 - 0x1
      12'hB92: dout  = 8'b00000001; // 2962 :   1 - 0x1
      12'hB93: dout  = 8'b00000001; // 2963 :   1 - 0x1
      12'hB94: dout  = 8'b00000011; // 2964 :   3 - 0x3
      12'hB95: dout  = 8'b00000011; // 2965 :   3 - 0x3
      12'hB96: dout  = 8'b00000111; // 2966 :   7 - 0x7
      12'hB97: dout  = 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout  = 8'b11111111; // 2968 : 255 - 0xff -- Background 0x73
      12'hB99: dout  = 8'b11111111; // 2969 : 255 - 0xff
      12'hB9A: dout  = 8'b11111111; // 2970 : 255 - 0xff
      12'hB9B: dout  = 8'b11111111; // 2971 : 255 - 0xff
      12'hB9C: dout  = 8'b11111111; // 2972 : 255 - 0xff
      12'hB9D: dout  = 8'b11111111; // 2973 : 255 - 0xff
      12'hB9E: dout  = 8'b11111111; // 2974 : 255 - 0xff
      12'hB9F: dout  = 8'b11111111; // 2975 : 255 - 0xff
      12'hBA0: dout  = 8'b10000001; // 2976 : 129 - 0x81 -- Background 0x74
      12'hBA1: dout  = 8'b11000001; // 2977 : 193 - 0xc1
      12'hBA2: dout  = 8'b11100011; // 2978 : 227 - 0xe3
      12'hBA3: dout  = 8'b11111111; // 2979 : 255 - 0xff
      12'hBA4: dout  = 8'b11111111; // 2980 : 255 - 0xff
      12'hBA5: dout  = 8'b11111111; // 2981 : 255 - 0xff
      12'hBA6: dout  = 8'b11111111; // 2982 : 255 - 0xff
      12'hBA7: dout  = 8'b11111110; // 2983 : 254 - 0xfe
      12'hBA8: dout  = 8'b11111111; // 2984 : 255 - 0xff -- Background 0x75
      12'hBA9: dout  = 8'b11111111; // 2985 : 255 - 0xff
      12'hBAA: dout  = 8'b11111111; // 2986 : 255 - 0xff
      12'hBAB: dout  = 8'b11111111; // 2987 : 255 - 0xff
      12'hBAC: dout  = 8'b11111111; // 2988 : 255 - 0xff
      12'hBAD: dout  = 8'b11111011; // 2989 : 251 - 0xfb
      12'hBAE: dout  = 8'b10110101; // 2990 : 181 - 0xb5
      12'hBAF: dout  = 8'b11001110; // 2991 : 206 - 0xce
      12'hBB0: dout  = 8'b11111111; // 2992 : 255 - 0xff -- Background 0x76
      12'hBB1: dout  = 8'b11111111; // 2993 : 255 - 0xff
      12'hBB2: dout  = 8'b11111111; // 2994 : 255 - 0xff
      12'hBB3: dout  = 8'b11111111; // 2995 : 255 - 0xff
      12'hBB4: dout  = 8'b11111111; // 2996 : 255 - 0xff
      12'hBB5: dout  = 8'b11011111; // 2997 : 223 - 0xdf
      12'hBB6: dout  = 8'b10101101; // 2998 : 173 - 0xad
      12'hBB7: dout  = 8'b01110011; // 2999 : 115 - 0x73
      12'hBB8: dout  = 8'b01110111; // 3000 : 119 - 0x77 -- Background 0x77
      12'hBB9: dout  = 8'b01110111; // 3001 : 119 - 0x77
      12'hBBA: dout  = 8'b01110111; // 3002 : 119 - 0x77
      12'hBBB: dout  = 8'b01110111; // 3003 : 119 - 0x77
      12'hBBC: dout  = 8'b01110111; // 3004 : 119 - 0x77
      12'hBBD: dout  = 8'b01110111; // 3005 : 119 - 0x77
      12'hBBE: dout  = 8'b01110111; // 3006 : 119 - 0x77
      12'hBBF: dout  = 8'b01110111; // 3007 : 119 - 0x77
      12'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout  = 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout  = 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout  = 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout  = 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout  = 8'b11111111; // 3015 : 255 - 0xff
      12'hBC8: dout  = 8'b01110111; // 3016 : 119 - 0x77 -- Background 0x79
      12'hBC9: dout  = 8'b01110111; // 3017 : 119 - 0x77
      12'hBCA: dout  = 8'b01110111; // 3018 : 119 - 0x77
      12'hBCB: dout  = 8'b01110111; // 3019 : 119 - 0x77
      12'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout  = 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout  = 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout  = 8'b00000001; // 3024 :   1 - 0x1 -- Background 0x7a
      12'hBD1: dout  = 8'b00000001; // 3025 :   1 - 0x1
      12'hBD2: dout  = 8'b00000001; // 3026 :   1 - 0x1
      12'hBD3: dout  = 8'b00011001; // 3027 :  25 - 0x19
      12'hBD4: dout  = 8'b00011101; // 3028 :  29 - 0x1d
      12'hBD5: dout  = 8'b00001101; // 3029 :  13 - 0xd
      12'hBD6: dout  = 8'b00000001; // 3030 :   1 - 0x1
      12'hBD7: dout  = 8'b11111110; // 3031 : 254 - 0xfe
      12'hBD8: dout  = 8'b00100000; // 3032 :  32 - 0x20 -- Background 0x7b
      12'hBD9: dout  = 8'b01111000; // 3033 : 120 - 0x78
      12'hBDA: dout  = 8'b01111111; // 3034 : 127 - 0x7f
      12'hBDB: dout  = 8'b11111110; // 3035 : 254 - 0xfe
      12'hBDC: dout  = 8'b11111110; // 3036 : 254 - 0xfe
      12'hBDD: dout  = 8'b11111110; // 3037 : 254 - 0xfe
      12'hBDE: dout  = 8'b11111110; // 3038 : 254 - 0xfe
      12'hBDF: dout  = 8'b11111110; // 3039 : 254 - 0xfe
      12'hBE0: dout  = 8'b00000100; // 3040 :   4 - 0x4 -- Background 0x7c
      12'hBE1: dout  = 8'b10011010; // 3041 : 154 - 0x9a
      12'hBE2: dout  = 8'b11111010; // 3042 : 250 - 0xfa
      12'hBE3: dout  = 8'b11111101; // 3043 : 253 - 0xfd
      12'hBE4: dout  = 8'b11111101; // 3044 : 253 - 0xfd
      12'hBE5: dout  = 8'b11111101; // 3045 : 253 - 0xfd
      12'hBE6: dout  = 8'b11111101; // 3046 : 253 - 0xfd
      12'hBE7: dout  = 8'b11111101; // 3047 : 253 - 0xfd
      12'hBE8: dout  = 8'b01111110; // 3048 : 126 - 0x7e -- Background 0x7d
      12'hBE9: dout  = 8'b00111000; // 3049 :  56 - 0x38
      12'hBEA: dout  = 8'b00100001; // 3050 :  33 - 0x21
      12'hBEB: dout  = 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout  = 8'b00000001; // 3052 :   1 - 0x1
      12'hBED: dout  = 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout  = 8'b00000001; // 3054 :   1 - 0x1
      12'hBEF: dout  = 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout  = 8'b11111010; // 3056 : 250 - 0xfa -- Background 0x7e
      12'hBF1: dout  = 8'b10001010; // 3057 : 138 - 0x8a
      12'hBF2: dout  = 8'b10000100; // 3058 : 132 - 0x84
      12'hBF3: dout  = 8'b10000000; // 3059 : 128 - 0x80
      12'hBF4: dout  = 8'b10000000; // 3060 : 128 - 0x80
      12'hBF5: dout  = 8'b10000000; // 3061 : 128 - 0x80
      12'hBF6: dout  = 8'b10000000; // 3062 : 128 - 0x80
      12'hBF7: dout  = 8'b10000000; // 3063 : 128 - 0x80
      12'hBF8: dout  = 8'b00000010; // 3064 :   2 - 0x2 -- Background 0x7f
      12'hBF9: dout  = 8'b00000100; // 3065 :   4 - 0x4
      12'hBFA: dout  = 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout  = 8'b00010000; // 3067 :  16 - 0x10
      12'hBFC: dout  = 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout  = 8'b01000000; // 3069 :  64 - 0x40
      12'hBFE: dout  = 8'b10000000; // 3070 : 128 - 0x80
      12'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout  = 8'b00001011; // 3072 :  11 - 0xb -- Background 0x80
      12'hC01: dout  = 8'b00001011; // 3073 :  11 - 0xb
      12'hC02: dout  = 8'b00111011; // 3074 :  59 - 0x3b
      12'hC03: dout  = 8'b00001011; // 3075 :  11 - 0xb
      12'hC04: dout  = 8'b11111011; // 3076 : 251 - 0xfb
      12'hC05: dout  = 8'b00001011; // 3077 :  11 - 0xb
      12'hC06: dout  = 8'b00001011; // 3078 :  11 - 0xb
      12'hC07: dout  = 8'b00001010; // 3079 :  10 - 0xa
      12'hC08: dout  = 8'b10010000; // 3080 : 144 - 0x90 -- Background 0x81
      12'hC09: dout  = 8'b00010000; // 3081 :  16 - 0x10
      12'hC0A: dout  = 8'b00011111; // 3082 :  31 - 0x1f
      12'hC0B: dout  = 8'b00010000; // 3083 :  16 - 0x10
      12'hC0C: dout  = 8'b00011111; // 3084 :  31 - 0x1f
      12'hC0D: dout  = 8'b00010000; // 3085 :  16 - 0x10
      12'hC0E: dout  = 8'b00010000; // 3086 :  16 - 0x10
      12'hC0F: dout  = 8'b10010000; // 3087 : 144 - 0x90
      12'hC10: dout  = 8'b00111111; // 3088 :  63 - 0x3f -- Background 0x82
      12'hC11: dout  = 8'b01111000; // 3089 : 120 - 0x78
      12'hC12: dout  = 8'b11100111; // 3090 : 231 - 0xe7
      12'hC13: dout  = 8'b11001111; // 3091 : 207 - 0xcf
      12'hC14: dout  = 8'b01011000; // 3092 :  88 - 0x58
      12'hC15: dout  = 8'b01011000; // 3093 :  88 - 0x58
      12'hC16: dout  = 8'b01010000; // 3094 :  80 - 0x50
      12'hC17: dout  = 8'b10010000; // 3095 : 144 - 0x90
      12'hC18: dout  = 8'b10110000; // 3096 : 176 - 0xb0 -- Background 0x83
      12'hC19: dout  = 8'b11111100; // 3097 : 252 - 0xfc
      12'hC1A: dout  = 8'b11100010; // 3098 : 226 - 0xe2
      12'hC1B: dout  = 8'b11000001; // 3099 : 193 - 0xc1
      12'hC1C: dout  = 8'b11000001; // 3100 : 193 - 0xc1
      12'hC1D: dout  = 8'b10000011; // 3101 : 131 - 0x83
      12'hC1E: dout  = 8'b10001111; // 3102 : 143 - 0x8f
      12'hC1F: dout  = 8'b01111110; // 3103 : 126 - 0x7e
      12'hC20: dout  = 8'b11111110; // 3104 : 254 - 0xfe -- Background 0x84
      12'hC21: dout  = 8'b00000011; // 3105 :   3 - 0x3
      12'hC22: dout  = 8'b00001111; // 3106 :  15 - 0xf
      12'hC23: dout  = 8'b10010001; // 3107 : 145 - 0x91
      12'hC24: dout  = 8'b01110000; // 3108 : 112 - 0x70
      12'hC25: dout  = 8'b01100000; // 3109 :  96 - 0x60
      12'hC26: dout  = 8'b00100000; // 3110 :  32 - 0x20
      12'hC27: dout  = 8'b00110001; // 3111 :  49 - 0x31
      12'hC28: dout  = 8'b00111111; // 3112 :  63 - 0x3f -- Background 0x85
      12'hC29: dout  = 8'b00111111; // 3113 :  63 - 0x3f
      12'hC2A: dout  = 8'b00011101; // 3114 :  29 - 0x1d
      12'hC2B: dout  = 8'b00111001; // 3115 :  57 - 0x39
      12'hC2C: dout  = 8'b01111011; // 3116 : 123 - 0x7b
      12'hC2D: dout  = 8'b11110011; // 3117 : 243 - 0xf3
      12'hC2E: dout  = 8'b10000110; // 3118 : 134 - 0x86
      12'hC2F: dout  = 8'b11111110; // 3119 : 254 - 0xfe
      12'hC30: dout  = 8'b11111111; // 3120 : 255 - 0xff -- Background 0x86
      12'hC31: dout  = 8'b11111111; // 3121 : 255 - 0xff
      12'hC32: dout  = 8'b11111111; // 3122 : 255 - 0xff
      12'hC33: dout  = 8'b11111111; // 3123 : 255 - 0xff
      12'hC34: dout  = 8'b11111111; // 3124 : 255 - 0xff
      12'hC35: dout  = 8'b10000000; // 3125 : 128 - 0x80
      12'hC36: dout  = 8'b10000000; // 3126 : 128 - 0x80
      12'hC37: dout  = 8'b11111111; // 3127 : 255 - 0xff
      12'hC38: dout  = 8'b11111110; // 3128 : 254 - 0xfe -- Background 0x87
      12'hC39: dout  = 8'b11111111; // 3129 : 255 - 0xff
      12'hC3A: dout  = 8'b11111111; // 3130 : 255 - 0xff
      12'hC3B: dout  = 8'b11111111; // 3131 : 255 - 0xff
      12'hC3C: dout  = 8'b11111111; // 3132 : 255 - 0xff
      12'hC3D: dout  = 8'b00000011; // 3133 :   3 - 0x3
      12'hC3E: dout  = 8'b00000011; // 3134 :   3 - 0x3
      12'hC3F: dout  = 8'b11111111; // 3135 : 255 - 0xff
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Background 0x88
      12'hC41: dout  = 8'b11111111; // 3137 : 255 - 0xff
      12'hC42: dout  = 8'b11111111; // 3138 : 255 - 0xff
      12'hC43: dout  = 8'b11111111; // 3139 : 255 - 0xff
      12'hC44: dout  = 8'b11111111; // 3140 : 255 - 0xff
      12'hC45: dout  = 8'b11111111; // 3141 : 255 - 0xff
      12'hC46: dout  = 8'b00000000; // 3142 :   0 - 0x0
      12'hC47: dout  = 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout  = 8'b00111100; // 3144 :  60 - 0x3c -- Background 0x89
      12'hC49: dout  = 8'b11111100; // 3145 : 252 - 0xfc
      12'hC4A: dout  = 8'b11111100; // 3146 : 252 - 0xfc
      12'hC4B: dout  = 8'b11111100; // 3147 : 252 - 0xfc
      12'hC4C: dout  = 8'b11111100; // 3148 : 252 - 0xfc
      12'hC4D: dout  = 8'b11111100; // 3149 : 252 - 0xfc
      12'hC4E: dout  = 8'b00000100; // 3150 :   4 - 0x4
      12'hC4F: dout  = 8'b00000100; // 3151 :   4 - 0x4
      12'hC50: dout  = 8'b11111111; // 3152 : 255 - 0xff -- Background 0x8a
      12'hC51: dout  = 8'b11111111; // 3153 : 255 - 0xff
      12'hC52: dout  = 8'b11111111; // 3154 : 255 - 0xff
      12'hC53: dout  = 8'b11111111; // 3155 : 255 - 0xff
      12'hC54: dout  = 8'b10000000; // 3156 : 128 - 0x80
      12'hC55: dout  = 8'b11111111; // 3157 : 255 - 0xff
      12'hC56: dout  = 8'b11111111; // 3158 : 255 - 0xff
      12'hC57: dout  = 8'b11111111; // 3159 : 255 - 0xff
      12'hC58: dout  = 8'b11111111; // 3160 : 255 - 0xff -- Background 0x8b
      12'hC59: dout  = 8'b11111111; // 3161 : 255 - 0xff
      12'hC5A: dout  = 8'b11111111; // 3162 : 255 - 0xff
      12'hC5B: dout  = 8'b11111111; // 3163 : 255 - 0xff
      12'hC5C: dout  = 8'b00000011; // 3164 :   3 - 0x3
      12'hC5D: dout  = 8'b11111111; // 3165 : 255 - 0xff
      12'hC5E: dout  = 8'b11111111; // 3166 : 255 - 0xff
      12'hC5F: dout  = 8'b11111111; // 3167 : 255 - 0xff
      12'hC60: dout  = 8'b11111111; // 3168 : 255 - 0xff -- Background 0x8c
      12'hC61: dout  = 8'b11111111; // 3169 : 255 - 0xff
      12'hC62: dout  = 8'b11111111; // 3170 : 255 - 0xff
      12'hC63: dout  = 8'b11111111; // 3171 : 255 - 0xff
      12'hC64: dout  = 8'b11111111; // 3172 : 255 - 0xff
      12'hC65: dout  = 8'b00000000; // 3173 :   0 - 0x0
      12'hC66: dout  = 8'b11111111; // 3174 : 255 - 0xff
      12'hC67: dout  = 8'b11111111; // 3175 : 255 - 0xff
      12'hC68: dout  = 8'b11111100; // 3176 : 252 - 0xfc -- Background 0x8d
      12'hC69: dout  = 8'b11111100; // 3177 : 252 - 0xfc
      12'hC6A: dout  = 8'b11111110; // 3178 : 254 - 0xfe
      12'hC6B: dout  = 8'b11111110; // 3179 : 254 - 0xfe
      12'hC6C: dout  = 8'b11111110; // 3180 : 254 - 0xfe
      12'hC6D: dout  = 8'b00000010; // 3181 :   2 - 0x2
      12'hC6E: dout  = 8'b11111110; // 3182 : 254 - 0xfe
      12'hC6F: dout  = 8'b11111110; // 3183 : 254 - 0xfe
      12'hC70: dout  = 8'b11111111; // 3184 : 255 - 0xff -- Background 0x8e
      12'hC71: dout  = 8'b10000000; // 3185 : 128 - 0x80
      12'hC72: dout  = 8'b10000000; // 3186 : 128 - 0x80
      12'hC73: dout  = 8'b10000000; // 3187 : 128 - 0x80
      12'hC74: dout  = 8'b10000000; // 3188 : 128 - 0x80
      12'hC75: dout  = 8'b10000000; // 3189 : 128 - 0x80
      12'hC76: dout  = 8'b10000000; // 3190 : 128 - 0x80
      12'hC77: dout  = 8'b10000000; // 3191 : 128 - 0x80
      12'hC78: dout  = 8'b11111111; // 3192 : 255 - 0xff -- Background 0x8f
      12'hC79: dout  = 8'b00000011; // 3193 :   3 - 0x3
      12'hC7A: dout  = 8'b00000011; // 3194 :   3 - 0x3
      12'hC7B: dout  = 8'b00000011; // 3195 :   3 - 0x3
      12'hC7C: dout  = 8'b00000011; // 3196 :   3 - 0x3
      12'hC7D: dout  = 8'b00000011; // 3197 :   3 - 0x3
      12'hC7E: dout  = 8'b00000011; // 3198 :   3 - 0x3
      12'hC7F: dout  = 8'b00000011; // 3199 :   3 - 0x3
      12'hC80: dout  = 8'b00000010; // 3200 :   2 - 0x2 -- Background 0x90
      12'hC81: dout  = 8'b00000010; // 3201 :   2 - 0x2
      12'hC82: dout  = 8'b00000010; // 3202 :   2 - 0x2
      12'hC83: dout  = 8'b00000010; // 3203 :   2 - 0x2
      12'hC84: dout  = 8'b00000010; // 3204 :   2 - 0x2
      12'hC85: dout  = 8'b00000010; // 3205 :   2 - 0x2
      12'hC86: dout  = 8'b00000100; // 3206 :   4 - 0x4
      12'hC87: dout  = 8'b00000100; // 3207 :   4 - 0x4
      12'hC88: dout  = 8'b10000000; // 3208 : 128 - 0x80 -- Background 0x91
      12'hC89: dout  = 8'b10000000; // 3209 : 128 - 0x80
      12'hC8A: dout  = 8'b10101010; // 3210 : 170 - 0xaa
      12'hC8B: dout  = 8'b11010101; // 3211 : 213 - 0xd5
      12'hC8C: dout  = 8'b10101010; // 3212 : 170 - 0xaa
      12'hC8D: dout  = 8'b11111111; // 3213 : 255 - 0xff
      12'hC8E: dout  = 8'b11111111; // 3214 : 255 - 0xff
      12'hC8F: dout  = 8'b11111111; // 3215 : 255 - 0xff
      12'hC90: dout  = 8'b00000011; // 3216 :   3 - 0x3 -- Background 0x92
      12'hC91: dout  = 8'b00000011; // 3217 :   3 - 0x3
      12'hC92: dout  = 8'b10101011; // 3218 : 171 - 0xab
      12'hC93: dout  = 8'b01010111; // 3219 :  87 - 0x57
      12'hC94: dout  = 8'b10101011; // 3220 : 171 - 0xab
      12'hC95: dout  = 8'b11111111; // 3221 : 255 - 0xff
      12'hC96: dout  = 8'b11111111; // 3222 : 255 - 0xff
      12'hC97: dout  = 8'b11111110; // 3223 : 254 - 0xfe
      12'hC98: dout  = 8'b00000000; // 3224 :   0 - 0x0 -- Background 0x93
      12'hC99: dout  = 8'b01010101; // 3225 :  85 - 0x55
      12'hC9A: dout  = 8'b10101010; // 3226 : 170 - 0xaa
      12'hC9B: dout  = 8'b01010101; // 3227 :  85 - 0x55
      12'hC9C: dout  = 8'b11111111; // 3228 : 255 - 0xff
      12'hC9D: dout  = 8'b11111111; // 3229 : 255 - 0xff
      12'hC9E: dout  = 8'b11111111; // 3230 : 255 - 0xff
      12'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout  = 8'b00000100; // 3232 :   4 - 0x4 -- Background 0x94
      12'hCA1: dout  = 8'b01010100; // 3233 :  84 - 0x54
      12'hCA2: dout  = 8'b10101100; // 3234 : 172 - 0xac
      12'hCA3: dout  = 8'b01011100; // 3235 :  92 - 0x5c
      12'hCA4: dout  = 8'b11111100; // 3236 : 252 - 0xfc
      12'hCA5: dout  = 8'b11111100; // 3237 : 252 - 0xfc
      12'hCA6: dout  = 8'b11111100; // 3238 : 252 - 0xfc
      12'hCA7: dout  = 8'b00111100; // 3239 :  60 - 0x3c
      12'hCA8: dout  = 8'b00111111; // 3240 :  63 - 0x3f -- Background 0x95
      12'hCA9: dout  = 8'b00111111; // 3241 :  63 - 0x3f
      12'hCAA: dout  = 8'b00111111; // 3242 :  63 - 0x3f
      12'hCAB: dout  = 8'b00111111; // 3243 :  63 - 0x3f
      12'hCAC: dout  = 8'b00000000; // 3244 :   0 - 0x0
      12'hCAD: dout  = 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout  = 8'b00000000; // 3246 :   0 - 0x0
      12'hCAF: dout  = 8'b11111111; // 3247 : 255 - 0xff
      12'hCB0: dout  = 8'b01111110; // 3248 : 126 - 0x7e -- Background 0x96
      12'hCB1: dout  = 8'b01111100; // 3249 : 124 - 0x7c
      12'hCB2: dout  = 8'b01111100; // 3250 : 124 - 0x7c
      12'hCB3: dout  = 8'b01111000; // 3251 : 120 - 0x78
      12'hCB4: dout  = 8'b00000000; // 3252 :   0 - 0x0
      12'hCB5: dout  = 8'b00000000; // 3253 :   0 - 0x0
      12'hCB6: dout  = 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout  = 8'b11111111; // 3255 : 255 - 0xff
      12'hCB8: dout  = 8'b00011111; // 3256 :  31 - 0x1f -- Background 0x97
      12'hCB9: dout  = 8'b00001111; // 3257 :  15 - 0xf
      12'hCBA: dout  = 8'b00001111; // 3258 :  15 - 0xf
      12'hCBB: dout  = 8'b00000111; // 3259 :   7 - 0x7
      12'hCBC: dout  = 8'b00000000; // 3260 :   0 - 0x0
      12'hCBD: dout  = 8'b00000000; // 3261 :   0 - 0x0
      12'hCBE: dout  = 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout  = 8'b11111111; // 3263 : 255 - 0xff
      12'hCC0: dout  = 8'b11111110; // 3264 : 254 - 0xfe -- Background 0x98
      12'hCC1: dout  = 8'b11111100; // 3265 : 252 - 0xfc
      12'hCC2: dout  = 8'b11111100; // 3266 : 252 - 0xfc
      12'hCC3: dout  = 8'b11111000; // 3267 : 248 - 0xf8
      12'hCC4: dout  = 8'b00000000; // 3268 :   0 - 0x0
      12'hCC5: dout  = 8'b00000000; // 3269 :   0 - 0x0
      12'hCC6: dout  = 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout  = 8'b00000000; // 3272 :   0 - 0x0 -- Background 0x99
      12'hCC9: dout  = 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout  = 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout  = 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      12'hCCD: dout  = 8'b11111111; // 3277 : 255 - 0xff
      12'hCCE: dout  = 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout  = 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout  = 8'b00011000; // 3280 :  24 - 0x18 -- Background 0x9a
      12'hCD1: dout  = 8'b00011000; // 3281 :  24 - 0x18
      12'hCD2: dout  = 8'b00011000; // 3282 :  24 - 0x18
      12'hCD3: dout  = 8'b00011000; // 3283 :  24 - 0x18
      12'hCD4: dout  = 8'b00011000; // 3284 :  24 - 0x18
      12'hCD5: dout  = 8'b00011000; // 3285 :  24 - 0x18
      12'hCD6: dout  = 8'b00011000; // 3286 :  24 - 0x18
      12'hCD7: dout  = 8'b00011000; // 3287 :  24 - 0x18
      12'hCD8: dout  = 8'b00000111; // 3288 :   7 - 0x7 -- Background 0x9b
      12'hCD9: dout  = 8'b00011111; // 3289 :  31 - 0x1f
      12'hCDA: dout  = 8'b00111111; // 3290 :  63 - 0x3f
      12'hCDB: dout  = 8'b11111111; // 3291 : 255 - 0xff
      12'hCDC: dout  = 8'b01111111; // 3292 : 127 - 0x7f
      12'hCDD: dout  = 8'b01111111; // 3293 : 127 - 0x7f
      12'hCDE: dout  = 8'b11111111; // 3294 : 255 - 0xff
      12'hCDF: dout  = 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout  = 8'b11100001; // 3296 : 225 - 0xe1 -- Background 0x9c
      12'hCE1: dout  = 8'b11111001; // 3297 : 249 - 0xf9
      12'hCE2: dout  = 8'b11111101; // 3298 : 253 - 0xfd
      12'hCE3: dout  = 8'b11111111; // 3299 : 255 - 0xff
      12'hCE4: dout  = 8'b11111110; // 3300 : 254 - 0xfe
      12'hCE5: dout  = 8'b11111110; // 3301 : 254 - 0xfe
      12'hCE6: dout  = 8'b11111111; // 3302 : 255 - 0xff
      12'hCE7: dout  = 8'b11111111; // 3303 : 255 - 0xff
      12'hCE8: dout  = 8'b11110000; // 3304 : 240 - 0xf0 -- Background 0x9d
      12'hCE9: dout  = 8'b00010000; // 3305 :  16 - 0x10
      12'hCEA: dout  = 8'b00010000; // 3306 :  16 - 0x10
      12'hCEB: dout  = 8'b00010000; // 3307 :  16 - 0x10
      12'hCEC: dout  = 8'b00010000; // 3308 :  16 - 0x10
      12'hCED: dout  = 8'b00010000; // 3309 :  16 - 0x10
      12'hCEE: dout  = 8'b00010000; // 3310 :  16 - 0x10
      12'hCEF: dout  = 8'b11111111; // 3311 : 255 - 0xff
      12'hCF0: dout  = 8'b00011111; // 3312 :  31 - 0x1f -- Background 0x9e
      12'hCF1: dout  = 8'b00010000; // 3313 :  16 - 0x10
      12'hCF2: dout  = 8'b00010000; // 3314 :  16 - 0x10
      12'hCF3: dout  = 8'b00010000; // 3315 :  16 - 0x10
      12'hCF4: dout  = 8'b00010000; // 3316 :  16 - 0x10
      12'hCF5: dout  = 8'b00010000; // 3317 :  16 - 0x10
      12'hCF6: dout  = 8'b00010000; // 3318 :  16 - 0x10
      12'hCF7: dout  = 8'b11111111; // 3319 : 255 - 0xff
      12'hCF8: dout  = 8'b10010010; // 3320 : 146 - 0x92 -- Background 0x9f
      12'hCF9: dout  = 8'b10010010; // 3321 : 146 - 0x92
      12'hCFA: dout  = 8'b10010010; // 3322 : 146 - 0x92
      12'hCFB: dout  = 8'b11111110; // 3323 : 254 - 0xfe
      12'hCFC: dout  = 8'b11111110; // 3324 : 254 - 0xfe
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00001010; // 3328 :  10 - 0xa -- Background 0xa0
      12'hD01: dout  = 8'b00001010; // 3329 :  10 - 0xa
      12'hD02: dout  = 8'b00111010; // 3330 :  58 - 0x3a
      12'hD03: dout  = 8'b00001010; // 3331 :  10 - 0xa
      12'hD04: dout  = 8'b11111011; // 3332 : 251 - 0xfb
      12'hD05: dout  = 8'b00001011; // 3333 :  11 - 0xb
      12'hD06: dout  = 8'b00001011; // 3334 :  11 - 0xb
      12'hD07: dout  = 8'b00001011; // 3335 :  11 - 0xb
      12'hD08: dout  = 8'b10010000; // 3336 : 144 - 0x90 -- Background 0xa1
      12'hD09: dout  = 8'b10010000; // 3337 : 144 - 0x90
      12'hD0A: dout  = 8'b10011111; // 3338 : 159 - 0x9f
      12'hD0B: dout  = 8'b10010000; // 3339 : 144 - 0x90
      12'hD0C: dout  = 8'b10011111; // 3340 : 159 - 0x9f
      12'hD0D: dout  = 8'b10010000; // 3341 : 144 - 0x90
      12'hD0E: dout  = 8'b10010000; // 3342 : 144 - 0x90
      12'hD0F: dout  = 8'b10010000; // 3343 : 144 - 0x90
      12'hD10: dout  = 8'b00000001; // 3344 :   1 - 0x1 -- Background 0xa2
      12'hD11: dout  = 8'b00000001; // 3345 :   1 - 0x1
      12'hD12: dout  = 8'b00000001; // 3346 :   1 - 0x1
      12'hD13: dout  = 8'b00000001; // 3347 :   1 - 0x1
      12'hD14: dout  = 8'b00000001; // 3348 :   1 - 0x1
      12'hD15: dout  = 8'b00000001; // 3349 :   1 - 0x1
      12'hD16: dout  = 8'b00000001; // 3350 :   1 - 0x1
      12'hD17: dout  = 8'b00000001; // 3351 :   1 - 0x1
      12'hD18: dout  = 8'b10000000; // 3352 : 128 - 0x80 -- Background 0xa3
      12'hD19: dout  = 8'b10000000; // 3353 : 128 - 0x80
      12'hD1A: dout  = 8'b10000000; // 3354 : 128 - 0x80
      12'hD1B: dout  = 8'b10000000; // 3355 : 128 - 0x80
      12'hD1C: dout  = 8'b10000000; // 3356 : 128 - 0x80
      12'hD1D: dout  = 8'b10000000; // 3357 : 128 - 0x80
      12'hD1E: dout  = 8'b10000000; // 3358 : 128 - 0x80
      12'hD1F: dout  = 8'b10000000; // 3359 : 128 - 0x80
      12'hD20: dout  = 8'b00001000; // 3360 :   8 - 0x8 -- Background 0xa4
      12'hD21: dout  = 8'b10001000; // 3361 : 136 - 0x88
      12'hD22: dout  = 8'b10010001; // 3362 : 145 - 0x91
      12'hD23: dout  = 8'b11010001; // 3363 : 209 - 0xd1
      12'hD24: dout  = 8'b01010011; // 3364 :  83 - 0x53
      12'hD25: dout  = 8'b01010011; // 3365 :  83 - 0x53
      12'hD26: dout  = 8'b01110011; // 3366 : 115 - 0x73
      12'hD27: dout  = 8'b00111111; // 3367 :  63 - 0x3f
      12'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0 -- Background 0xa5
      12'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout  = 8'b00000111; // 3370 :   7 - 0x7
      12'hD2B: dout  = 8'b00001111; // 3371 :  15 - 0xf
      12'hD2C: dout  = 8'b00001100; // 3372 :  12 - 0xc
      12'hD2D: dout  = 8'b00011011; // 3373 :  27 - 0x1b
      12'hD2E: dout  = 8'b00011011; // 3374 :  27 - 0x1b
      12'hD2F: dout  = 8'b00011011; // 3375 :  27 - 0x1b
      12'hD30: dout  = 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xa6
      12'hD31: dout  = 8'b00000000; // 3377 :   0 - 0x0
      12'hD32: dout  = 8'b11100000; // 3378 : 224 - 0xe0
      12'hD33: dout  = 8'b11110000; // 3379 : 240 - 0xf0
      12'hD34: dout  = 8'b11110000; // 3380 : 240 - 0xf0
      12'hD35: dout  = 8'b11111000; // 3381 : 248 - 0xf8
      12'hD36: dout  = 8'b11111000; // 3382 : 248 - 0xf8
      12'hD37: dout  = 8'b11111000; // 3383 : 248 - 0xf8
      12'hD38: dout  = 8'b00011011; // 3384 :  27 - 0x1b -- Background 0xa7
      12'hD39: dout  = 8'b00011011; // 3385 :  27 - 0x1b
      12'hD3A: dout  = 8'b00011011; // 3386 :  27 - 0x1b
      12'hD3B: dout  = 8'b00011011; // 3387 :  27 - 0x1b
      12'hD3C: dout  = 8'b00011011; // 3388 :  27 - 0x1b
      12'hD3D: dout  = 8'b00001111; // 3389 :  15 - 0xf
      12'hD3E: dout  = 8'b00001111; // 3390 :  15 - 0xf
      12'hD3F: dout  = 8'b00000111; // 3391 :   7 - 0x7
      12'hD40: dout  = 8'b11111000; // 3392 : 248 - 0xf8 -- Background 0xa8
      12'hD41: dout  = 8'b11111000; // 3393 : 248 - 0xf8
      12'hD42: dout  = 8'b11111000; // 3394 : 248 - 0xf8
      12'hD43: dout  = 8'b11111000; // 3395 : 248 - 0xf8
      12'hD44: dout  = 8'b11111000; // 3396 : 248 - 0xf8
      12'hD45: dout  = 8'b11110000; // 3397 : 240 - 0xf0
      12'hD46: dout  = 8'b11110000; // 3398 : 240 - 0xf0
      12'hD47: dout  = 8'b11100000; // 3399 : 224 - 0xe0
      12'hD48: dout  = 8'b11110001; // 3400 : 241 - 0xf1 -- Background 0xa9
      12'hD49: dout  = 8'b00010001; // 3401 :  17 - 0x11
      12'hD4A: dout  = 8'b00010001; // 3402 :  17 - 0x11
      12'hD4B: dout  = 8'b00011111; // 3403 :  31 - 0x1f
      12'hD4C: dout  = 8'b00010000; // 3404 :  16 - 0x10
      12'hD4D: dout  = 8'b00010000; // 3405 :  16 - 0x10
      12'hD4E: dout  = 8'b00010000; // 3406 :  16 - 0x10
      12'hD4F: dout  = 8'b11111111; // 3407 : 255 - 0xff
      12'hD50: dout  = 8'b00011111; // 3408 :  31 - 0x1f -- Background 0xaa
      12'hD51: dout  = 8'b00010000; // 3409 :  16 - 0x10
      12'hD52: dout  = 8'b00010000; // 3410 :  16 - 0x10
      12'hD53: dout  = 8'b11110000; // 3411 : 240 - 0xf0
      12'hD54: dout  = 8'b00010000; // 3412 :  16 - 0x10
      12'hD55: dout  = 8'b00010000; // 3413 :  16 - 0x10
      12'hD56: dout  = 8'b00010000; // 3414 :  16 - 0x10
      12'hD57: dout  = 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout  = 8'b01111111; // 3416 : 127 - 0x7f -- Background 0xab
      12'hD59: dout  = 8'b10111111; // 3417 : 191 - 0xbf
      12'hD5A: dout  = 8'b11011111; // 3418 : 223 - 0xdf
      12'hD5B: dout  = 8'b11101111; // 3419 : 239 - 0xef
      12'hD5C: dout  = 8'b11110000; // 3420 : 240 - 0xf0
      12'hD5D: dout  = 8'b11110000; // 3421 : 240 - 0xf0
      12'hD5E: dout  = 8'b11110000; // 3422 : 240 - 0xf0
      12'hD5F: dout  = 8'b11110000; // 3423 : 240 - 0xf0
      12'hD60: dout  = 8'b11110000; // 3424 : 240 - 0xf0 -- Background 0xac
      12'hD61: dout  = 8'b11110000; // 3425 : 240 - 0xf0
      12'hD62: dout  = 8'b11110000; // 3426 : 240 - 0xf0
      12'hD63: dout  = 8'b11110000; // 3427 : 240 - 0xf0
      12'hD64: dout  = 8'b11111111; // 3428 : 255 - 0xff
      12'hD65: dout  = 8'b11111111; // 3429 : 255 - 0xff
      12'hD66: dout  = 8'b11111111; // 3430 : 255 - 0xff
      12'hD67: dout  = 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout  = 8'b11111111; // 3432 : 255 - 0xff -- Background 0xad
      12'hD69: dout  = 8'b11111111; // 3433 : 255 - 0xff
      12'hD6A: dout  = 8'b11111111; // 3434 : 255 - 0xff
      12'hD6B: dout  = 8'b11111111; // 3435 : 255 - 0xff
      12'hD6C: dout  = 8'b00001111; // 3436 :  15 - 0xf
      12'hD6D: dout  = 8'b00001111; // 3437 :  15 - 0xf
      12'hD6E: dout  = 8'b00001111; // 3438 :  15 - 0xf
      12'hD6F: dout  = 8'b00001111; // 3439 :  15 - 0xf
      12'hD70: dout  = 8'b00001111; // 3440 :  15 - 0xf -- Background 0xae
      12'hD71: dout  = 8'b00001111; // 3441 :  15 - 0xf
      12'hD72: dout  = 8'b00001111; // 3442 :  15 - 0xf
      12'hD73: dout  = 8'b00001111; // 3443 :  15 - 0xf
      12'hD74: dout  = 8'b11110111; // 3444 : 247 - 0xf7
      12'hD75: dout  = 8'b11111011; // 3445 : 251 - 0xfb
      12'hD76: dout  = 8'b11111101; // 3446 : 253 - 0xfd
      12'hD77: dout  = 8'b11111110; // 3447 : 254 - 0xfe
      12'hD78: dout  = 8'b00000000; // 3448 :   0 - 0x0 -- Background 0xaf
      12'hD79: dout  = 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout  = 8'b00000000; // 3450 :   0 - 0x0
      12'hD7B: dout  = 8'b00000000; // 3451 :   0 - 0x0
      12'hD7C: dout  = 8'b00000000; // 3452 :   0 - 0x0
      12'hD7D: dout  = 8'b00000000; // 3453 :   0 - 0x0
      12'hD7E: dout  = 8'b00011000; // 3454 :  24 - 0x18
      12'hD7F: dout  = 8'b00011000; // 3455 :  24 - 0x18
      12'hD80: dout  = 8'b00011111; // 3456 :  31 - 0x1f -- Background 0xb0
      12'hD81: dout  = 8'b00111111; // 3457 :  63 - 0x3f
      12'hD82: dout  = 8'b01111111; // 3458 : 127 - 0x7f
      12'hD83: dout  = 8'b01111111; // 3459 : 127 - 0x7f
      12'hD84: dout  = 8'b01111111; // 3460 : 127 - 0x7f
      12'hD85: dout  = 8'b11111111; // 3461 : 255 - 0xff
      12'hD86: dout  = 8'b11111111; // 3462 : 255 - 0xff
      12'hD87: dout  = 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout  = 8'b11111111; // 3464 : 255 - 0xff -- Background 0xb1
      12'hD89: dout  = 8'b11111111; // 3465 : 255 - 0xff
      12'hD8A: dout  = 8'b11111111; // 3466 : 255 - 0xff
      12'hD8B: dout  = 8'b01111111; // 3467 : 127 - 0x7f
      12'hD8C: dout  = 8'b01111111; // 3468 : 127 - 0x7f
      12'hD8D: dout  = 8'b01111111; // 3469 : 127 - 0x7f
      12'hD8E: dout  = 8'b00111111; // 3470 :  63 - 0x3f
      12'hD8F: dout  = 8'b00011110; // 3471 :  30 - 0x1e
      12'hD90: dout  = 8'b11111000; // 3472 : 248 - 0xf8 -- Background 0xb2
      12'hD91: dout  = 8'b11111100; // 3473 : 252 - 0xfc
      12'hD92: dout  = 8'b11111110; // 3474 : 254 - 0xfe
      12'hD93: dout  = 8'b11111110; // 3475 : 254 - 0xfe
      12'hD94: dout  = 8'b11111110; // 3476 : 254 - 0xfe
      12'hD95: dout  = 8'b11111111; // 3477 : 255 - 0xff
      12'hD96: dout  = 8'b11111111; // 3478 : 255 - 0xff
      12'hD97: dout  = 8'b11111111; // 3479 : 255 - 0xff
      12'hD98: dout  = 8'b11111111; // 3480 : 255 - 0xff -- Background 0xb3
      12'hD99: dout  = 8'b11111111; // 3481 : 255 - 0xff
      12'hD9A: dout  = 8'b11111111; // 3482 : 255 - 0xff
      12'hD9B: dout  = 8'b11111110; // 3483 : 254 - 0xfe
      12'hD9C: dout  = 8'b11111110; // 3484 : 254 - 0xfe
      12'hD9D: dout  = 8'b11111110; // 3485 : 254 - 0xfe
      12'hD9E: dout  = 8'b11111100; // 3486 : 252 - 0xfc
      12'hD9F: dout  = 8'b01111000; // 3487 : 120 - 0x78
      12'hDA0: dout  = 8'b01111111; // 3488 : 127 - 0x7f -- Background 0xb4
      12'hDA1: dout  = 8'b10000000; // 3489 : 128 - 0x80
      12'hDA2: dout  = 8'b10000000; // 3490 : 128 - 0x80
      12'hDA3: dout  = 8'b10000000; // 3491 : 128 - 0x80
      12'hDA4: dout  = 8'b10000000; // 3492 : 128 - 0x80
      12'hDA5: dout  = 8'b10000000; // 3493 : 128 - 0x80
      12'hDA6: dout  = 8'b10000000; // 3494 : 128 - 0x80
      12'hDA7: dout  = 8'b10000000; // 3495 : 128 - 0x80
      12'hDA8: dout  = 8'b11011110; // 3496 : 222 - 0xde -- Background 0xb5
      12'hDA9: dout  = 8'b01100001; // 3497 :  97 - 0x61
      12'hDAA: dout  = 8'b01100001; // 3498 :  97 - 0x61
      12'hDAB: dout  = 8'b01100001; // 3499 :  97 - 0x61
      12'hDAC: dout  = 8'b01110001; // 3500 : 113 - 0x71
      12'hDAD: dout  = 8'b01011110; // 3501 :  94 - 0x5e
      12'hDAE: dout  = 8'b01111111; // 3502 : 127 - 0x7f
      12'hDAF: dout  = 8'b01100001; // 3503 :  97 - 0x61
      12'hDB0: dout  = 8'b10000000; // 3504 : 128 - 0x80 -- Background 0xb6
      12'hDB1: dout  = 8'b10000000; // 3505 : 128 - 0x80
      12'hDB2: dout  = 8'b11000000; // 3506 : 192 - 0xc0
      12'hDB3: dout  = 8'b11110000; // 3507 : 240 - 0xf0
      12'hDB4: dout  = 8'b10111111; // 3508 : 191 - 0xbf
      12'hDB5: dout  = 8'b10001111; // 3509 : 143 - 0x8f
      12'hDB6: dout  = 8'b10000001; // 3510 : 129 - 0x81
      12'hDB7: dout  = 8'b01111110; // 3511 : 126 - 0x7e
      12'hDB8: dout  = 8'b01100001; // 3512 :  97 - 0x61 -- Background 0xb7
      12'hDB9: dout  = 8'b01100001; // 3513 :  97 - 0x61
      12'hDBA: dout  = 8'b11000001; // 3514 : 193 - 0xc1
      12'hDBB: dout  = 8'b11000001; // 3515 : 193 - 0xc1
      12'hDBC: dout  = 8'b10000001; // 3516 : 129 - 0x81
      12'hDBD: dout  = 8'b10000001; // 3517 : 129 - 0x81
      12'hDBE: dout  = 8'b10000011; // 3518 : 131 - 0x83
      12'hDBF: dout  = 8'b11111110; // 3519 : 254 - 0xfe
      12'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout  = 8'b00000011; // 3522 :   3 - 0x3
      12'hDC3: dout  = 8'b00001111; // 3523 :  15 - 0xf
      12'hDC4: dout  = 8'b00011111; // 3524 :  31 - 0x1f
      12'hDC5: dout  = 8'b00111111; // 3525 :  63 - 0x3f
      12'hDC6: dout  = 8'b01111111; // 3526 : 127 - 0x7f
      12'hDC7: dout  = 8'b01111111; // 3527 : 127 - 0x7f
      12'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0 -- Background 0xb9
      12'hDC9: dout  = 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout  = 8'b11000000; // 3530 : 192 - 0xc0
      12'hDCB: dout  = 8'b11110000; // 3531 : 240 - 0xf0
      12'hDCC: dout  = 8'b11111000; // 3532 : 248 - 0xf8
      12'hDCD: dout  = 8'b11111100; // 3533 : 252 - 0xfc
      12'hDCE: dout  = 8'b11111110; // 3534 : 254 - 0xfe
      12'hDCF: dout  = 8'b11111110; // 3535 : 254 - 0xfe
      12'hDD0: dout  = 8'b11111111; // 3536 : 255 - 0xff -- Background 0xba
      12'hDD1: dout  = 8'b11111111; // 3537 : 255 - 0xff
      12'hDD2: dout  = 8'b11111111; // 3538 : 255 - 0xff
      12'hDD3: dout  = 8'b11111111; // 3539 : 255 - 0xff
      12'hDD4: dout  = 8'b11111111; // 3540 : 255 - 0xff
      12'hDD5: dout  = 8'b11111111; // 3541 : 255 - 0xff
      12'hDD6: dout  = 8'b11111111; // 3542 : 255 - 0xff
      12'hDD7: dout  = 8'b11111111; // 3543 : 255 - 0xff
      12'hDD8: dout  = 8'b11111111; // 3544 : 255 - 0xff -- Background 0xbb
      12'hDD9: dout  = 8'b11111111; // 3545 : 255 - 0xff
      12'hDDA: dout  = 8'b11111111; // 3546 : 255 - 0xff
      12'hDDB: dout  = 8'b11111111; // 3547 : 255 - 0xff
      12'hDDC: dout  = 8'b11111111; // 3548 : 255 - 0xff
      12'hDDD: dout  = 8'b11111111; // 3549 : 255 - 0xff
      12'hDDE: dout  = 8'b11111111; // 3550 : 255 - 0xff
      12'hDDF: dout  = 8'b11111111; // 3551 : 255 - 0xff
      12'hDE0: dout  = 8'b01111111; // 3552 : 127 - 0x7f -- Background 0xbc
      12'hDE1: dout  = 8'b01111111; // 3553 : 127 - 0x7f
      12'hDE2: dout  = 8'b01111111; // 3554 : 127 - 0x7f
      12'hDE3: dout  = 8'b00111111; // 3555 :  63 - 0x3f
      12'hDE4: dout  = 8'b00111111; // 3556 :  63 - 0x3f
      12'hDE5: dout  = 8'b00011111; // 3557 :  31 - 0x1f
      12'hDE6: dout  = 8'b00001111; // 3558 :  15 - 0xf
      12'hDE7: dout  = 8'b00000111; // 3559 :   7 - 0x7
      12'hDE8: dout  = 8'b11111110; // 3560 : 254 - 0xfe -- Background 0xbd
      12'hDE9: dout  = 8'b11111110; // 3561 : 254 - 0xfe
      12'hDEA: dout  = 8'b11111110; // 3562 : 254 - 0xfe
      12'hDEB: dout  = 8'b11111100; // 3563 : 252 - 0xfc
      12'hDEC: dout  = 8'b11111100; // 3564 : 252 - 0xfc
      12'hDED: dout  = 8'b11111000; // 3565 : 248 - 0xf8
      12'hDEE: dout  = 8'b11110000; // 3566 : 240 - 0xf0
      12'hDEF: dout  = 8'b11110000; // 3567 : 240 - 0xf0
      12'hDF0: dout  = 8'b00001111; // 3568 :  15 - 0xf -- Background 0xbe
      12'hDF1: dout  = 8'b00001111; // 3569 :  15 - 0xf
      12'hDF2: dout  = 8'b00001111; // 3570 :  15 - 0xf
      12'hDF3: dout  = 8'b00001111; // 3571 :  15 - 0xf
      12'hDF4: dout  = 8'b00001111; // 3572 :  15 - 0xf
      12'hDF5: dout  = 8'b00001111; // 3573 :  15 - 0xf
      12'hDF6: dout  = 8'b00000111; // 3574 :   7 - 0x7
      12'hDF7: dout  = 8'b00001111; // 3575 :  15 - 0xf
      12'hDF8: dout  = 8'b11110000; // 3576 : 240 - 0xf0 -- Background 0xbf
      12'hDF9: dout  = 8'b11110000; // 3577 : 240 - 0xf0
      12'hDFA: dout  = 8'b11110000; // 3578 : 240 - 0xf0
      12'hDFB: dout  = 8'b11110000; // 3579 : 240 - 0xf0
      12'hDFC: dout  = 8'b11110000; // 3580 : 240 - 0xf0
      12'hDFD: dout  = 8'b11110000; // 3581 : 240 - 0xf0
      12'hDFE: dout  = 8'b11100000; // 3582 : 224 - 0xe0
      12'hDFF: dout  = 8'b11110000; // 3583 : 240 - 0xf0
      12'hE00: dout  = 8'b10000001; // 3584 : 129 - 0x81 -- Background 0xc0
      12'hE01: dout  = 8'b11000001; // 3585 : 193 - 0xc1
      12'hE02: dout  = 8'b10100011; // 3586 : 163 - 0xa3
      12'hE03: dout  = 8'b10100011; // 3587 : 163 - 0xa3
      12'hE04: dout  = 8'b10011101; // 3588 : 157 - 0x9d
      12'hE05: dout  = 8'b10000001; // 3589 : 129 - 0x81
      12'hE06: dout  = 8'b10000001; // 3590 : 129 - 0x81
      12'hE07: dout  = 8'b10000001; // 3591 : 129 - 0x81
      12'hE08: dout  = 8'b11100011; // 3592 : 227 - 0xe3 -- Background 0xc1
      12'hE09: dout  = 8'b11110111; // 3593 : 247 - 0xf7
      12'hE0A: dout  = 8'b11000001; // 3594 : 193 - 0xc1
      12'hE0B: dout  = 8'b11000001; // 3595 : 193 - 0xc1
      12'hE0C: dout  = 8'b11000001; // 3596 : 193 - 0xc1
      12'hE0D: dout  = 8'b11000001; // 3597 : 193 - 0xc1
      12'hE0E: dout  = 8'b11110111; // 3598 : 247 - 0xf7
      12'hE0F: dout  = 8'b11100011; // 3599 : 227 - 0xe3
      12'hE10: dout  = 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout  = 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout  = 8'b00000111; // 3602 :   7 - 0x7
      12'hE13: dout  = 8'b00001111; // 3603 :  15 - 0xf
      12'hE14: dout  = 8'b00001100; // 3604 :  12 - 0xc
      12'hE15: dout  = 8'b00011011; // 3605 :  27 - 0x1b
      12'hE16: dout  = 8'b00011011; // 3606 :  27 - 0x1b
      12'hE17: dout  = 8'b00011011; // 3607 :  27 - 0x1b
      12'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0 -- Background 0xc3
      12'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout  = 8'b11100000; // 3610 : 224 - 0xe0
      12'hE1B: dout  = 8'b11110000; // 3611 : 240 - 0xf0
      12'hE1C: dout  = 8'b11110000; // 3612 : 240 - 0xf0
      12'hE1D: dout  = 8'b11111000; // 3613 : 248 - 0xf8
      12'hE1E: dout  = 8'b11111000; // 3614 : 248 - 0xf8
      12'hE1F: dout  = 8'b11111000; // 3615 : 248 - 0xf8
      12'hE20: dout  = 8'b00011011; // 3616 :  27 - 0x1b -- Background 0xc4
      12'hE21: dout  = 8'b00011011; // 3617 :  27 - 0x1b
      12'hE22: dout  = 8'b00011011; // 3618 :  27 - 0x1b
      12'hE23: dout  = 8'b00011011; // 3619 :  27 - 0x1b
      12'hE24: dout  = 8'b00011011; // 3620 :  27 - 0x1b
      12'hE25: dout  = 8'b00001111; // 3621 :  15 - 0xf
      12'hE26: dout  = 8'b00001111; // 3622 :  15 - 0xf
      12'hE27: dout  = 8'b00000111; // 3623 :   7 - 0x7
      12'hE28: dout  = 8'b11111000; // 3624 : 248 - 0xf8 -- Background 0xc5
      12'hE29: dout  = 8'b11111000; // 3625 : 248 - 0xf8
      12'hE2A: dout  = 8'b11111000; // 3626 : 248 - 0xf8
      12'hE2B: dout  = 8'b11111000; // 3627 : 248 - 0xf8
      12'hE2C: dout  = 8'b11111000; // 3628 : 248 - 0xf8
      12'hE2D: dout  = 8'b11110000; // 3629 : 240 - 0xf0
      12'hE2E: dout  = 8'b11110000; // 3630 : 240 - 0xf0
      12'hE2F: dout  = 8'b11100000; // 3631 : 224 - 0xe0
      12'hE30: dout  = 8'b11100000; // 3632 : 224 - 0xe0 -- Background 0xc6
      12'hE31: dout  = 8'b11111111; // 3633 : 255 - 0xff
      12'hE32: dout  = 8'b11111111; // 3634 : 255 - 0xff
      12'hE33: dout  = 8'b11111111; // 3635 : 255 - 0xff
      12'hE34: dout  = 8'b11111111; // 3636 : 255 - 0xff
      12'hE35: dout  = 8'b11111111; // 3637 : 255 - 0xff
      12'hE36: dout  = 8'b11111111; // 3638 : 255 - 0xff
      12'hE37: dout  = 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout  = 8'b00000111; // 3640 :   7 - 0x7 -- Background 0xc7
      12'hE39: dout  = 8'b11111111; // 3641 : 255 - 0xff
      12'hE3A: dout  = 8'b11111111; // 3642 : 255 - 0xff
      12'hE3B: dout  = 8'b11111111; // 3643 : 255 - 0xff
      12'hE3C: dout  = 8'b11111111; // 3644 : 255 - 0xff
      12'hE3D: dout  = 8'b11111111; // 3645 : 255 - 0xff
      12'hE3E: dout  = 8'b11111111; // 3646 : 255 - 0xff
      12'hE3F: dout  = 8'b11111111; // 3647 : 255 - 0xff
      12'hE40: dout  = 8'b11111111; // 3648 : 255 - 0xff -- Background 0xc8
      12'hE41: dout  = 8'b11111111; // 3649 : 255 - 0xff
      12'hE42: dout  = 8'b11111111; // 3650 : 255 - 0xff
      12'hE43: dout  = 8'b11111111; // 3651 : 255 - 0xff
      12'hE44: dout  = 8'b11111111; // 3652 : 255 - 0xff
      12'hE45: dout  = 8'b11111110; // 3653 : 254 - 0xfe
      12'hE46: dout  = 8'b11111111; // 3654 : 255 - 0xff
      12'hE47: dout  = 8'b11101111; // 3655 : 239 - 0xef
      12'hE48: dout  = 8'b11111111; // 3656 : 255 - 0xff -- Background 0xc9
      12'hE49: dout  = 8'b11011111; // 3657 : 223 - 0xdf
      12'hE4A: dout  = 8'b11101111; // 3658 : 239 - 0xef
      12'hE4B: dout  = 8'b10101111; // 3659 : 175 - 0xaf
      12'hE4C: dout  = 8'b10101111; // 3660 : 175 - 0xaf
      12'hE4D: dout  = 8'b01101111; // 3661 : 111 - 0x6f
      12'hE4E: dout  = 8'b11101111; // 3662 : 239 - 0xef
      12'hE4F: dout  = 8'b11100111; // 3663 : 231 - 0xe7
      12'hE50: dout  = 8'b00011111; // 3664 :  31 - 0x1f -- Background 0xca
      12'hE51: dout  = 8'b00011111; // 3665 :  31 - 0x1f
      12'hE52: dout  = 8'b00111111; // 3666 :  63 - 0x3f
      12'hE53: dout  = 8'b00111111; // 3667 :  63 - 0x3f
      12'hE54: dout  = 8'b01110000; // 3668 : 112 - 0x70
      12'hE55: dout  = 8'b01100011; // 3669 :  99 - 0x63
      12'hE56: dout  = 8'b11100111; // 3670 : 231 - 0xe7
      12'hE57: dout  = 8'b11100101; // 3671 : 229 - 0xe5
      12'hE58: dout  = 8'b11110000; // 3672 : 240 - 0xf0 -- Background 0xcb
      12'hE59: dout  = 8'b11110000; // 3673 : 240 - 0xf0
      12'hE5A: dout  = 8'b11111000; // 3674 : 248 - 0xf8
      12'hE5B: dout  = 8'b11111000; // 3675 : 248 - 0xf8
      12'hE5C: dout  = 8'b00001100; // 3676 :  12 - 0xc
      12'hE5D: dout  = 8'b11000100; // 3677 : 196 - 0xc4
      12'hE5E: dout  = 8'b11100100; // 3678 : 228 - 0xe4
      12'hE5F: dout  = 8'b10100110; // 3679 : 166 - 0xa6
      12'hE60: dout  = 8'b11101001; // 3680 : 233 - 0xe9 -- Background 0xcc
      12'hE61: dout  = 8'b11101001; // 3681 : 233 - 0xe9
      12'hE62: dout  = 8'b11101001; // 3682 : 233 - 0xe9
      12'hE63: dout  = 8'b11101111; // 3683 : 239 - 0xef
      12'hE64: dout  = 8'b11100010; // 3684 : 226 - 0xe2
      12'hE65: dout  = 8'b11100011; // 3685 : 227 - 0xe3
      12'hE66: dout  = 8'b11110000; // 3686 : 240 - 0xf0
      12'hE67: dout  = 8'b11111111; // 3687 : 255 - 0xff
      12'hE68: dout  = 8'b10010110; // 3688 : 150 - 0x96 -- Background 0xcd
      12'hE69: dout  = 8'b10010110; // 3689 : 150 - 0x96
      12'hE6A: dout  = 8'b10010110; // 3690 : 150 - 0x96
      12'hE6B: dout  = 8'b11110110; // 3691 : 246 - 0xf6
      12'hE6C: dout  = 8'b01000110; // 3692 :  70 - 0x46
      12'hE6D: dout  = 8'b11000110; // 3693 : 198 - 0xc6
      12'hE6E: dout  = 8'b00001110; // 3694 :  14 - 0xe
      12'hE6F: dout  = 8'b11111110; // 3695 : 254 - 0xfe
      12'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout  = 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout  = 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout  = 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout  = 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout  = 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout  = 8'b01111110; // 3702 : 126 - 0x7e
      12'hE77: dout  = 8'b00111100; // 3703 :  60 - 0x3c
      12'hE78: dout  = 8'b00111100; // 3704 :  60 - 0x3c -- Background 0xcf
      12'hE79: dout  = 8'b01000010; // 3705 :  66 - 0x42
      12'hE7A: dout  = 8'b10011001; // 3706 : 153 - 0x99
      12'hE7B: dout  = 8'b10100001; // 3707 : 161 - 0xa1
      12'hE7C: dout  = 8'b10100001; // 3708 : 161 - 0xa1
      12'hE7D: dout  = 8'b10011001; // 3709 : 153 - 0x99
      12'hE7E: dout  = 8'b01000010; // 3710 :  66 - 0x42
      12'hE7F: dout  = 8'b00111100; // 3711 :  60 - 0x3c
      12'hE80: dout  = 8'b00001111; // 3712 :  15 - 0xf -- Background 0xd0
      12'hE81: dout  = 8'b00011111; // 3713 :  31 - 0x1f
      12'hE82: dout  = 8'b00011111; // 3714 :  31 - 0x1f
      12'hE83: dout  = 8'b00111111; // 3715 :  63 - 0x3f
      12'hE84: dout  = 8'b00111111; // 3716 :  63 - 0x3f
      12'hE85: dout  = 8'b01111111; // 3717 : 127 - 0x7f
      12'hE86: dout  = 8'b01111111; // 3718 : 127 - 0x7f
      12'hE87: dout  = 8'b01111111; // 3719 : 127 - 0x7f
      12'hE88: dout  = 8'b11110000; // 3720 : 240 - 0xf0 -- Background 0xd1
      12'hE89: dout  = 8'b11111000; // 3721 : 248 - 0xf8
      12'hE8A: dout  = 8'b11111000; // 3722 : 248 - 0xf8
      12'hE8B: dout  = 8'b11111100; // 3723 : 252 - 0xfc
      12'hE8C: dout  = 8'b11111100; // 3724 : 252 - 0xfc
      12'hE8D: dout  = 8'b11111110; // 3725 : 254 - 0xfe
      12'hE8E: dout  = 8'b11111110; // 3726 : 254 - 0xfe
      12'hE8F: dout  = 8'b11111110; // 3727 : 254 - 0xfe
      12'hE90: dout  = 8'b01111111; // 3728 : 127 - 0x7f -- Background 0xd2
      12'hE91: dout  = 8'b01111111; // 3729 : 127 - 0x7f
      12'hE92: dout  = 8'b00111111; // 3730 :  63 - 0x3f
      12'hE93: dout  = 8'b00111111; // 3731 :  63 - 0x3f
      12'hE94: dout  = 8'b00111111; // 3732 :  63 - 0x3f
      12'hE95: dout  = 8'b00111111; // 3733 :  63 - 0x3f
      12'hE96: dout  = 8'b00011111; // 3734 :  31 - 0x1f
      12'hE97: dout  = 8'b00011111; // 3735 :  31 - 0x1f
      12'hE98: dout  = 8'b11111110; // 3736 : 254 - 0xfe -- Background 0xd3
      12'hE99: dout  = 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout  = 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout  = 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout  = 8'b11111100; // 3740 : 252 - 0xfc
      12'hE9D: dout  = 8'b11111100; // 3741 : 252 - 0xfc
      12'hE9E: dout  = 8'b11111110; // 3742 : 254 - 0xfe
      12'hE9F: dout  = 8'b11111110; // 3743 : 254 - 0xfe
      12'hEA0: dout  = 8'b01111111; // 3744 : 127 - 0x7f -- Background 0xd4
      12'hEA1: dout  = 8'b01111111; // 3745 : 127 - 0x7f
      12'hEA2: dout  = 8'b01111111; // 3746 : 127 - 0x7f
      12'hEA3: dout  = 8'b00111111; // 3747 :  63 - 0x3f
      12'hEA4: dout  = 8'b00111111; // 3748 :  63 - 0x3f
      12'hEA5: dout  = 8'b00111111; // 3749 :  63 - 0x3f
      12'hEA6: dout  = 8'b00111111; // 3750 :  63 - 0x3f
      12'hEA7: dout  = 8'b00011111; // 3751 :  31 - 0x1f
      12'hEA8: dout  = 8'b11111110; // 3752 : 254 - 0xfe -- Background 0xd5
      12'hEA9: dout  = 8'b11111110; // 3753 : 254 - 0xfe
      12'hEAA: dout  = 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout  = 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout  = 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout  = 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout  = 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout  = 8'b11111110; // 3759 : 254 - 0xfe
      12'hEB0: dout  = 8'b00011111; // 3760 :  31 - 0x1f -- Background 0xd6
      12'hEB1: dout  = 8'b00001111; // 3761 :  15 - 0xf
      12'hEB2: dout  = 8'b00001111; // 3762 :  15 - 0xf
      12'hEB3: dout  = 8'b00000111; // 3763 :   7 - 0x7
      12'hEB4: dout  = 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout  = 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout  = 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout  = 8'b11111110; // 3768 : 254 - 0xfe -- Background 0xd7
      12'hEB9: dout  = 8'b11111100; // 3769 : 252 - 0xfc
      12'hEBA: dout  = 8'b11111100; // 3770 : 252 - 0xfc
      12'hEBB: dout  = 8'b11111000; // 3771 : 248 - 0xf8
      12'hEBC: dout  = 8'b00000000; // 3772 :   0 - 0x0
      12'hEBD: dout  = 8'b00000000; // 3773 :   0 - 0x0
      12'hEBE: dout  = 8'b00000000; // 3774 :   0 - 0x0
      12'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout  = 8'b01111110; // 3776 : 126 - 0x7e -- Background 0xd8
      12'hEC1: dout  = 8'b01111110; // 3777 : 126 - 0x7e
      12'hEC2: dout  = 8'b01111110; // 3778 : 126 - 0x7e
      12'hEC3: dout  = 8'b01111110; // 3779 : 126 - 0x7e
      12'hEC4: dout  = 8'b01111111; // 3780 : 127 - 0x7f
      12'hEC5: dout  = 8'b01111111; // 3781 : 127 - 0x7f
      12'hEC6: dout  = 8'b01111111; // 3782 : 127 - 0x7f
      12'hEC7: dout  = 8'b01111111; // 3783 : 127 - 0x7f
      12'hEC8: dout  = 8'b11111111; // 3784 : 255 - 0xff -- Background 0xd9
      12'hEC9: dout  = 8'b11111111; // 3785 : 255 - 0xff
      12'hECA: dout  = 8'b11111111; // 3786 : 255 - 0xff
      12'hECB: dout  = 8'b11111111; // 3787 : 255 - 0xff
      12'hECC: dout  = 8'b11111111; // 3788 : 255 - 0xff
      12'hECD: dout  = 8'b11111111; // 3789 : 255 - 0xff
      12'hECE: dout  = 8'b11111111; // 3790 : 255 - 0xff
      12'hECF: dout  = 8'b11111110; // 3791 : 254 - 0xfe
      12'hED0: dout  = 8'b11111110; // 3792 : 254 - 0xfe -- Background 0xda
      12'hED1: dout  = 8'b11111110; // 3793 : 254 - 0xfe
      12'hED2: dout  = 8'b11111110; // 3794 : 254 - 0xfe
      12'hED3: dout  = 8'b11111110; // 3795 : 254 - 0xfe
      12'hED4: dout  = 8'b11111111; // 3796 : 255 - 0xff
      12'hED5: dout  = 8'b11111111; // 3797 : 255 - 0xff
      12'hED6: dout  = 8'b11111111; // 3798 : 255 - 0xff
      12'hED7: dout  = 8'b11111111; // 3799 : 255 - 0xff
      12'hED8: dout  = 8'b01111111; // 3800 : 127 - 0x7f -- Background 0xdb
      12'hED9: dout  = 8'b01111111; // 3801 : 127 - 0x7f
      12'hEDA: dout  = 8'b01111111; // 3802 : 127 - 0x7f
      12'hEDB: dout  = 8'b01111111; // 3803 : 127 - 0x7f
      12'hEDC: dout  = 8'b01111111; // 3804 : 127 - 0x7f
      12'hEDD: dout  = 8'b01111111; // 3805 : 127 - 0x7f
      12'hEDE: dout  = 8'b01111111; // 3806 : 127 - 0x7f
      12'hEDF: dout  = 8'b01111111; // 3807 : 127 - 0x7f
      12'hEE0: dout  = 8'b11111111; // 3808 : 255 - 0xff -- Background 0xdc
      12'hEE1: dout  = 8'b11111111; // 3809 : 255 - 0xff
      12'hEE2: dout  = 8'b11111111; // 3810 : 255 - 0xff
      12'hEE3: dout  = 8'b11111111; // 3811 : 255 - 0xff
      12'hEE4: dout  = 8'b11111100; // 3812 : 252 - 0xfc
      12'hEE5: dout  = 8'b11111110; // 3813 : 254 - 0xfe
      12'hEE6: dout  = 8'b11111110; // 3814 : 254 - 0xfe
      12'hEE7: dout  = 8'b01111110; // 3815 : 126 - 0x7e
      12'hEE8: dout  = 8'b11111111; // 3816 : 255 - 0xff -- Background 0xdd
      12'hEE9: dout  = 8'b11111111; // 3817 : 255 - 0xff
      12'hEEA: dout  = 8'b11111111; // 3818 : 255 - 0xff
      12'hEEB: dout  = 8'b11111111; // 3819 : 255 - 0xff
      12'hEEC: dout  = 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout  = 8'b00000000; // 3821 :   0 - 0x0
      12'hEEE: dout  = 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout  = 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout  = 8'b01111111; // 3824 : 127 - 0x7f -- Background 0xde
      12'hEF1: dout  = 8'b01111111; // 3825 : 127 - 0x7f
      12'hEF2: dout  = 8'b01111111; // 3826 : 127 - 0x7f
      12'hEF3: dout  = 8'b01111111; // 3827 : 127 - 0x7f
      12'hEF4: dout  = 8'b01111111; // 3828 : 127 - 0x7f
      12'hEF5: dout  = 8'b01111111; // 3829 : 127 - 0x7f
      12'hEF6: dout  = 8'b01111111; // 3830 : 127 - 0x7f
      12'hEF7: dout  = 8'b01111111; // 3831 : 127 - 0x7f
      12'hEF8: dout  = 8'b11111111; // 3832 : 255 - 0xff -- Background 0xdf
      12'hEF9: dout  = 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout  = 8'b11111111; // 3834 : 255 - 0xff
      12'hEFB: dout  = 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout  = 8'b11111111; // 3836 : 255 - 0xff
      12'hEFD: dout  = 8'b11111111; // 3837 : 255 - 0xff
      12'hEFE: dout  = 8'b11111111; // 3838 : 255 - 0xff
      12'hEFF: dout  = 8'b11111110; // 3839 : 254 - 0xfe
      12'hF00: dout  = 8'b01111110; // 3840 : 126 - 0x7e -- Background 0xe0
      12'hF01: dout  = 8'b01111110; // 3841 : 126 - 0x7e
      12'hF02: dout  = 8'b01111111; // 3842 : 127 - 0x7f
      12'hF03: dout  = 8'b01111111; // 3843 : 127 - 0x7f
      12'hF04: dout  = 8'b01111111; // 3844 : 127 - 0x7f
      12'hF05: dout  = 8'b01111111; // 3845 : 127 - 0x7f
      12'hF06: dout  = 8'b01111111; // 3846 : 127 - 0x7f
      12'hF07: dout  = 8'b01111111; // 3847 : 127 - 0x7f
      12'hF08: dout  = 8'b00111111; // 3848 :  63 - 0x3f -- Background 0xe1
      12'hF09: dout  = 8'b00111111; // 3849 :  63 - 0x3f
      12'hF0A: dout  = 8'b00111111; // 3850 :  63 - 0x3f
      12'hF0B: dout  = 8'b00111111; // 3851 :  63 - 0x3f
      12'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b01111110; // 3856 : 126 - 0x7e -- Background 0xe2
      12'hF11: dout  = 8'b01111100; // 3857 : 124 - 0x7c
      12'hF12: dout  = 8'b01111100; // 3858 : 124 - 0x7c
      12'hF13: dout  = 8'b01111000; // 3859 : 120 - 0x78
      12'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b11111110; // 3864 : 254 - 0xfe -- Background 0xe3
      12'hF19: dout  = 8'b11111110; // 3865 : 254 - 0xfe
      12'hF1A: dout  = 8'b11111111; // 3866 : 255 - 0xff
      12'hF1B: dout  = 8'b11111111; // 3867 : 255 - 0xff
      12'hF1C: dout  = 8'b01111111; // 3868 : 127 - 0x7f
      12'hF1D: dout  = 8'b01111111; // 3869 : 127 - 0x7f
      12'hF1E: dout  = 8'b01111111; // 3870 : 127 - 0x7f
      12'hF1F: dout  = 8'b01111111; // 3871 : 127 - 0x7f
      12'hF20: dout  = 8'b01111111; // 3872 : 127 - 0x7f -- Background 0xe4
      12'hF21: dout  = 8'b01111111; // 3873 : 127 - 0x7f
      12'hF22: dout  = 8'b00111111; // 3874 :  63 - 0x3f
      12'hF23: dout  = 8'b00111111; // 3875 :  63 - 0x3f
      12'hF24: dout  = 8'b00111111; // 3876 :  63 - 0x3f
      12'hF25: dout  = 8'b00111111; // 3877 :  63 - 0x3f
      12'hF26: dout  = 8'b00011111; // 3878 :  31 - 0x1f
      12'hF27: dout  = 8'b00011111; // 3879 :  31 - 0x1f
      12'hF28: dout  = 8'b00111111; // 3880 :  63 - 0x3f -- Background 0xe5
      12'hF29: dout  = 8'b10111111; // 3881 : 191 - 0xbf
      12'hF2A: dout  = 8'b11111111; // 3882 : 255 - 0xff
      12'hF2B: dout  = 8'b11111111; // 3883 : 255 - 0xff
      12'hF2C: dout  = 8'b11111100; // 3884 : 252 - 0xfc
      12'hF2D: dout  = 8'b11111100; // 3885 : 252 - 0xfc
      12'hF2E: dout  = 8'b11111110; // 3886 : 254 - 0xfe
      12'hF2F: dout  = 8'b11111110; // 3887 : 254 - 0xfe
      12'hF30: dout  = 8'b01111111; // 3888 : 127 - 0x7f -- Background 0xe6
      12'hF31: dout  = 8'b01111111; // 3889 : 127 - 0x7f
      12'hF32: dout  = 8'b01111110; // 3890 : 126 - 0x7e
      12'hF33: dout  = 8'b01111110; // 3891 : 126 - 0x7e
      12'hF34: dout  = 8'b01111111; // 3892 : 127 - 0x7f
      12'hF35: dout  = 8'b01111111; // 3893 : 127 - 0x7f
      12'hF36: dout  = 8'b01111111; // 3894 : 127 - 0x7f
      12'hF37: dout  = 8'b01111111; // 3895 : 127 - 0x7f
      12'hF38: dout  = 8'b01111110; // 3896 : 126 - 0x7e -- Background 0xe7
      12'hF39: dout  = 8'b01111110; // 3897 : 126 - 0x7e
      12'hF3A: dout  = 8'b01111110; // 3898 : 126 - 0x7e
      12'hF3B: dout  = 8'b01111110; // 3899 : 126 - 0x7e
      12'hF3C: dout  = 8'b01111111; // 3900 : 127 - 0x7f
      12'hF3D: dout  = 8'b01111111; // 3901 : 127 - 0x7f
      12'hF3E: dout  = 8'b01111111; // 3902 : 127 - 0x7f
      12'hF3F: dout  = 8'b01111111; // 3903 : 127 - 0x7f
      12'hF40: dout  = 8'b10000001; // 3904 : 129 - 0x81 -- Background 0xe8
      12'hF41: dout  = 8'b11000011; // 3905 : 195 - 0xc3
      12'hF42: dout  = 8'b11000011; // 3906 : 195 - 0xc3
      12'hF43: dout  = 8'b11100111; // 3907 : 231 - 0xe7
      12'hF44: dout  = 8'b11100111; // 3908 : 231 - 0xe7
      12'hF45: dout  = 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout  = 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout  = 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout  = 8'b00001111; // 3912 :  15 - 0xf -- Background 0xe9
      12'hF49: dout  = 8'b01000011; // 3913 :  67 - 0x43
      12'hF4A: dout  = 8'b01011011; // 3914 :  91 - 0x5b
      12'hF4B: dout  = 8'b01010011; // 3915 :  83 - 0x53
      12'hF4C: dout  = 8'b00110001; // 3916 :  49 - 0x31
      12'hF4D: dout  = 8'b00011001; // 3917 :  25 - 0x19
      12'hF4E: dout  = 8'b00001111; // 3918 :  15 - 0xf
      12'hF4F: dout  = 8'b00000111; // 3919 :   7 - 0x7
      12'hF50: dout  = 8'b11000001; // 3920 : 193 - 0xc1 -- Background 0xea
      12'hF51: dout  = 8'b11000011; // 3921 : 195 - 0xc3
      12'hF52: dout  = 8'b11000110; // 3922 : 198 - 0xc6
      12'hF53: dout  = 8'b10000100; // 3923 : 132 - 0x84
      12'hF54: dout  = 8'b11111100; // 3924 : 252 - 0xfc
      12'hF55: dout  = 8'b11111100; // 3925 : 252 - 0xfc
      12'hF56: dout  = 8'b00001110; // 3926 :  14 - 0xe
      12'hF57: dout  = 8'b00000010; // 3927 :   2 - 0x2
      12'hF58: dout  = 8'b00010000; // 3928 :  16 - 0x10 -- Background 0xeb
      12'hF59: dout  = 8'b00100000; // 3929 :  32 - 0x20
      12'hF5A: dout  = 8'b00100010; // 3930 :  34 - 0x22
      12'hF5B: dout  = 8'b10111010; // 3931 : 186 - 0xba
      12'hF5C: dout  = 8'b11100110; // 3932 : 230 - 0xe6
      12'hF5D: dout  = 8'b11100001; // 3933 : 225 - 0xe1
      12'hF5E: dout  = 8'b11000000; // 3934 : 192 - 0xc0
      12'hF5F: dout  = 8'b11000000; // 3935 : 192 - 0xc0
      12'hF60: dout  = 8'b00100000; // 3936 :  32 - 0x20 -- Background 0xec
      12'hF61: dout  = 8'b10100110; // 3937 : 166 - 0xa6
      12'hF62: dout  = 8'b01010100; // 3938 :  84 - 0x54
      12'hF63: dout  = 8'b00100110; // 3939 :  38 - 0x26
      12'hF64: dout  = 8'b00100000; // 3940 :  32 - 0x20
      12'hF65: dout  = 8'b11000110; // 3941 : 198 - 0xc6
      12'hF66: dout  = 8'b01010100; // 3942 :  84 - 0x54
      12'hF67: dout  = 8'b00100110; // 3943 :  38 - 0x26
      12'hF68: dout  = 8'b00100000; // 3944 :  32 - 0x20 -- Background 0xed
      12'hF69: dout  = 8'b10000101; // 3945 : 133 - 0x85
      12'hF6A: dout  = 8'b00000001; // 3946 :   1 - 0x1
      12'hF6B: dout  = 8'b01000100; // 3947 :  68 - 0x44
      12'hF6C: dout  = 8'b00100000; // 3948 :  32 - 0x20
      12'hF6D: dout  = 8'b10000110; // 3949 : 134 - 0x86
      12'hF6E: dout  = 8'b01010100; // 3950 :  84 - 0x54
      12'hF6F: dout  = 8'b01001000; // 3951 :  72 - 0x48
      12'hF70: dout  = 8'b00100000; // 3952 :  32 - 0x20 -- Background 0xee
      12'hF71: dout  = 8'b10111010; // 3953 : 186 - 0xba
      12'hF72: dout  = 8'b11001001; // 3954 : 201 - 0xc9
      12'hF73: dout  = 8'b01001010; // 3955 :  74 - 0x4a
      12'hF74: dout  = 8'b00100000; // 3956 :  32 - 0x20
      12'hF75: dout  = 8'b10100110; // 3957 : 166 - 0xa6
      12'hF76: dout  = 8'b00001010; // 3958 :  10 - 0xa
      12'hF77: dout  = 8'b11010000; // 3959 : 208 - 0xd0
      12'hF78: dout  = 8'b11010001; // 3960 : 209 - 0xd1 -- Background 0xef
      12'hF79: dout  = 8'b00100000; // 3961 :  32 - 0x20
      12'hF7A: dout  = 8'b11000110; // 3962 : 198 - 0xc6
      12'hF7B: dout  = 8'b00001010; // 3963 :  10 - 0xa
      12'hF7C: dout  = 8'b11010010; // 3964 : 210 - 0xd2
      12'hF7D: dout  = 8'b11010011; // 3965 : 211 - 0xd3
      12'hF7E: dout  = 8'b11011011; // 3966 : 219 - 0xdb
      12'hF7F: dout  = 8'b11011011; // 3967 : 219 - 0xdb
      12'hF80: dout  = 8'b00001010; // 3968 :  10 - 0xa -- Background 0xf0
      12'hF81: dout  = 8'b11010100; // 3969 : 212 - 0xd4
      12'hF82: dout  = 8'b11010101; // 3970 : 213 - 0xd5
      12'hF83: dout  = 8'b11010100; // 3971 : 212 - 0xd4
      12'hF84: dout  = 8'b11011001; // 3972 : 217 - 0xd9
      12'hF85: dout  = 8'b11011011; // 3973 : 219 - 0xdb
      12'hF86: dout  = 8'b11100010; // 3974 : 226 - 0xe2
      12'hF87: dout  = 8'b11010100; // 3975 : 212 - 0xd4
      12'hF88: dout  = 8'b11010110; // 3976 : 214 - 0xd6 -- Background 0xf1
      12'hF89: dout  = 8'b11010111; // 3977 : 215 - 0xd7
      12'hF8A: dout  = 8'b11100001; // 3978 : 225 - 0xe1
      12'hF8B: dout  = 8'b00100110; // 3979 :  38 - 0x26
      12'hF8C: dout  = 8'b11010110; // 3980 : 214 - 0xd6
      12'hF8D: dout  = 8'b11011101; // 3981 : 221 - 0xdd
      12'hF8E: dout  = 8'b11100001; // 3982 : 225 - 0xe1
      12'hF8F: dout  = 8'b11100001; // 3983 : 225 - 0xe1
      12'hF90: dout  = 8'b11011110; // 3984 : 222 - 0xde -- Background 0xf2
      12'hF91: dout  = 8'b11010001; // 3985 : 209 - 0xd1
      12'hF92: dout  = 8'b11011000; // 3986 : 216 - 0xd8
      12'hF93: dout  = 8'b11010000; // 3987 : 208 - 0xd0
      12'hF94: dout  = 8'b11010001; // 3988 : 209 - 0xd1
      12'hF95: dout  = 8'b00100110; // 3989 :  38 - 0x26
      12'hF96: dout  = 8'b11011110; // 3990 : 222 - 0xde
      12'hF97: dout  = 8'b11010001; // 3991 : 209 - 0xd1
      12'hF98: dout  = 8'b01000110; // 3992 :  70 - 0x46 -- Background 0xf3
      12'hF99: dout  = 8'b00010100; // 3993 :  20 - 0x14
      12'hF9A: dout  = 8'b11011011; // 3994 : 219 - 0xdb
      12'hF9B: dout  = 8'b01000010; // 3995 :  66 - 0x42
      12'hF9C: dout  = 8'b01000010; // 3996 :  66 - 0x42
      12'hF9D: dout  = 8'b11011011; // 3997 : 219 - 0xdb
      12'hF9E: dout  = 8'b01000010; // 3998 :  66 - 0x42
      12'hF9F: dout  = 8'b11011011; // 3999 : 219 - 0xdb
      12'hFA0: dout  = 8'b01000010; // 4000 :  66 - 0x42 -- Background 0xf4
      12'hFA1: dout  = 8'b11011011; // 4001 : 219 - 0xdb
      12'hFA2: dout  = 8'b01000010; // 4002 :  66 - 0x42
      12'hFA3: dout  = 8'b11011011; // 4003 : 219 - 0xdb
      12'hFA4: dout  = 8'b01000010; // 4004 :  66 - 0x42
      12'hFA5: dout  = 8'b00100110; // 4005 :  38 - 0x26
      12'hFA6: dout  = 8'b00100001; // 4006 :  33 - 0x21
      12'hFA7: dout  = 8'b01100110; // 4007 : 102 - 0x66
      12'hFA8: dout  = 8'b11011011; // 4008 : 219 - 0xdb -- Background 0xf5
      12'hFA9: dout  = 8'b00100110; // 4009 :  38 - 0x26
      12'hFAA: dout  = 8'b11011011; // 4010 : 219 - 0xdb
      12'hFAB: dout  = 8'b11011111; // 4011 : 223 - 0xdf
      12'hFAC: dout  = 8'b11011011; // 4012 : 219 - 0xdb
      12'hFAD: dout  = 8'b11011111; // 4013 : 223 - 0xdf
      12'hFAE: dout  = 8'b11011011; // 4014 : 219 - 0xdb
      12'hFAF: dout  = 8'b11011011; // 4015 : 219 - 0xdb
      12'hFB0: dout  = 8'b11011011; // 4016 : 219 - 0xdb -- Background 0xf6
      12'hFB1: dout  = 8'b11011110; // 4017 : 222 - 0xde
      12'hFB2: dout  = 8'b01000011; // 4018 :  67 - 0x43
      12'hFB3: dout  = 8'b11011011; // 4019 : 219 - 0xdb
      12'hFB4: dout  = 8'b11100000; // 4020 : 224 - 0xe0
      12'hFB5: dout  = 8'b11011011; // 4021 : 219 - 0xdb
      12'hFB6: dout  = 8'b11011011; // 4022 : 219 - 0xdb
      12'hFB7: dout  = 8'b11011011; // 4023 : 219 - 0xdb
      12'hFB8: dout  = 8'b11100011; // 4024 : 227 - 0xe3 -- Background 0xf7
      12'hFB9: dout  = 8'b00100110; // 4025 :  38 - 0x26
      12'hFBA: dout  = 8'b00100001; // 4026 :  33 - 0x21
      12'hFBB: dout  = 8'b10100110; // 4027 : 166 - 0xa6
      12'hFBC: dout  = 8'b00010100; // 4028 :  20 - 0x14
      12'hFBD: dout  = 8'b11011011; // 4029 : 219 - 0xdb
      12'hFBE: dout  = 8'b11011011; // 4030 : 219 - 0xdb
      12'hFBF: dout  = 8'b11011011; // 4031 : 219 - 0xdb
      12'hFC0: dout  = 8'b11011011; // 4032 : 219 - 0xdb -- Background 0xf8
      12'hFC1: dout  = 8'b11011001; // 4033 : 217 - 0xd9
      12'hFC2: dout  = 8'b11011011; // 4034 : 219 - 0xdb
      12'hFC3: dout  = 8'b11011011; // 4035 : 219 - 0xdb
      12'hFC4: dout  = 8'b11010100; // 4036 : 212 - 0xd4
      12'hFC5: dout  = 8'b11011001; // 4037 : 217 - 0xd9
      12'hFC6: dout  = 8'b11010100; // 4038 : 212 - 0xd4
      12'hFC7: dout  = 8'b11011001; // 4039 : 217 - 0xd9
      12'hFC8: dout  = 8'b10010101; // 4040 : 149 - 0x95 -- Background 0xf9
      12'hFC9: dout  = 8'b10010101; // 4041 : 149 - 0x95
      12'hFCA: dout  = 8'b10010101; // 4042 : 149 - 0x95
      12'hFCB: dout  = 8'b10010101; // 4043 : 149 - 0x95
      12'hFCC: dout  = 8'b10010101; // 4044 : 149 - 0x95
      12'hFCD: dout  = 8'b10010111; // 4045 : 151 - 0x97
      12'hFCE: dout  = 8'b10011000; // 4046 : 152 - 0x98
      12'hFCF: dout  = 8'b01111000; // 4047 : 120 - 0x78
      12'hFD0: dout  = 8'b10010101; // 4048 : 149 - 0x95 -- Background 0xfa
      12'hFD1: dout  = 8'b01111010; // 4049 : 122 - 0x7a
      12'hFD2: dout  = 8'b00100001; // 4050 :  33 - 0x21
      12'hFD3: dout  = 8'b11101101; // 4051 : 237 - 0xed
      12'hFD4: dout  = 8'b00001110; // 4052 :  14 - 0xe
      12'hFD5: dout  = 8'b11001111; // 4053 : 207 - 0xcf
      12'hFD6: dout  = 8'b00000001; // 4054 :   1 - 0x1
      12'hFD7: dout  = 8'b00001001; // 4055 :   9 - 0x9
      12'hFD8: dout  = 8'b00010111; // 4056 :  23 - 0x17 -- Background 0xfb
      12'hFD9: dout  = 8'b00001101; // 4057 :  13 - 0xd
      12'hFDA: dout  = 8'b00011000; // 4058 :  24 - 0x18
      12'hFDB: dout  = 8'b00100010; // 4059 :  34 - 0x22
      12'hFDC: dout  = 8'b01001011; // 4060 :  75 - 0x4b
      12'hFDD: dout  = 8'b00001101; // 4061 :  13 - 0xd
      12'hFDE: dout  = 8'b00000001; // 4062 :   1 - 0x1
      12'hFDF: dout  = 8'b00100100; // 4063 :  36 - 0x24
      12'hFE0: dout  = 8'b00001010; // 4064 :  10 - 0xa -- Background 0xfc
      12'hFE1: dout  = 8'b00010110; // 4065 :  22 - 0x16
      12'hFE2: dout  = 8'b00001110; // 4066 :  14 - 0xe
      12'hFE3: dout  = 8'b00100010; // 4067 :  34 - 0x22
      12'hFE4: dout  = 8'b10001011; // 4068 : 139 - 0x8b
      12'hFE5: dout  = 8'b00001101; // 4069 :  13 - 0xd
      12'hFE6: dout  = 8'b00000010; // 4070 :   2 - 0x2
      12'hFE7: dout  = 8'b00100100; // 4071 :  36 - 0x24
      12'hFE8: dout  = 8'b00001010; // 4072 :  10 - 0xa -- Background 0xfd
      12'hFE9: dout  = 8'b00010110; // 4073 :  22 - 0x16
      12'hFEA: dout  = 8'b00001110; // 4074 :  14 - 0xe
      12'hFEB: dout  = 8'b00100010; // 4075 :  34 - 0x22
      12'hFEC: dout  = 8'b11101100; // 4076 : 236 - 0xec
      12'hFED: dout  = 8'b00000100; // 4077 :   4 - 0x4
      12'hFEE: dout  = 8'b00011101; // 4078 :  29 - 0x1d
      12'hFEF: dout  = 8'b00011000; // 4079 :  24 - 0x18
      12'hFF0: dout  = 8'b01010110; // 4080 :  86 - 0x56 -- Background 0xfe
      12'hFF1: dout  = 8'b01010101; // 4081 :  85 - 0x55
      12'hFF2: dout  = 8'b00100011; // 4082 :  35 - 0x23
      12'hFF3: dout  = 8'b11100010; // 4083 : 226 - 0xe2
      12'hFF4: dout  = 8'b00000100; // 4084 :   4 - 0x4
      12'hFF5: dout  = 8'b10011001; // 4085 : 153 - 0x99
      12'hFF6: dout  = 8'b10101010; // 4086 : 170 - 0xaa
      12'hFF7: dout  = 8'b10101010; // 4087 : 170 - 0xaa
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout  = 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout  = 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout  = 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout  = 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout  = 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout  = 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout  = 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
