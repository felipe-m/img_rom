//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA
  (
     //input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      13'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      13'h2: dout  = 8'b00000100; //    2 :   4 - 0x4
      13'h3: dout  = 8'b00000011; //    3 :   3 - 0x3
      13'h4: dout  = 8'b00000011; //    4 :   3 - 0x3
      13'h5: dout  = 8'b00000011; //    5 :   3 - 0x3
      13'h6: dout  = 8'b00000100; //    6 :   4 - 0x4
      13'h7: dout  = 8'b00111010; //    7 :  58 - 0x3a
      13'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout  = 8'b00000011; //   10 :   3 - 0x3
      13'hB: dout  = 8'b00000001; //   11 :   1 - 0x1
      13'hC: dout  = 8'b00000001; //   12 :   1 - 0x1
      13'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      13'hE: dout  = 8'b00000011; //   14 :   3 - 0x3
      13'hF: dout  = 8'b00000001; //   15 :   1 - 0x1
      13'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      13'h11: dout  = 8'b00111000; //   17 :  56 - 0x38
      13'h12: dout  = 8'b11000110; //   18 : 198 - 0xc6
      13'h13: dout  = 8'b11001011; //   19 : 203 - 0xcb
      13'h14: dout  = 8'b11011100; //   20 : 220 - 0xdc
      13'h15: dout  = 8'b00111010; //   21 :  58 - 0x3a
      13'h16: dout  = 8'b10011010; //   22 : 154 - 0x9a
      13'h17: dout  = 8'b10000001; //   23 : 129 - 0x81
      13'h18: dout  = 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      13'h1A: dout  = 8'b00111000; //   26 :  56 - 0x38
      13'h1B: dout  = 8'b10110100; //   27 : 180 - 0xb4
      13'h1C: dout  = 8'b10101000; //   28 : 168 - 0xa8
      13'h1D: dout  = 8'b11010100; //   29 : 212 - 0xd4
      13'h1E: dout  = 8'b01110100; //   30 : 116 - 0x74
      13'h1F: dout  = 8'b01111110; //   31 : 126 - 0x7e
      13'h20: dout  = 8'b01000101; //   32 :  69 - 0x45 -- Sprite 0x2
      13'h21: dout  = 8'b10000111; //   33 : 135 - 0x87
      13'h22: dout  = 8'b10000011; //   34 : 131 - 0x83
      13'h23: dout  = 8'b10000001; //   35 : 129 - 0x81
      13'h24: dout  = 8'b10000001; //   36 : 129 - 0x81
      13'h25: dout  = 8'b10000001; //   37 : 129 - 0x81
      13'h26: dout  = 8'b01000001; //   38 :  65 - 0x41
      13'h27: dout  = 8'b00100001; //   39 :  33 - 0x21
      13'h28: dout  = 8'b00111000; //   40 :  56 - 0x38
      13'h29: dout  = 8'b01111000; //   41 : 120 - 0x78
      13'h2A: dout  = 8'b01111100; //   42 : 124 - 0x7c
      13'h2B: dout  = 8'b01111110; //   43 : 126 - 0x7e
      13'h2C: dout  = 8'b01111110; //   44 : 126 - 0x7e
      13'h2D: dout  = 8'b01111110; //   45 : 126 - 0x7e
      13'h2E: dout  = 8'b00111110; //   46 :  62 - 0x3e
      13'h2F: dout  = 8'b00011110; //   47 :  30 - 0x1e
      13'h30: dout  = 8'b01111111; //   48 : 127 - 0x7f -- Sprite 0x3
      13'h31: dout  = 8'b01111110; //   49 : 126 - 0x7e
      13'h32: dout  = 8'b11111100; //   50 : 252 - 0xfc
      13'h33: dout  = 8'b00111000; //   51 :  56 - 0x38
      13'h34: dout  = 8'b00011000; //   52 :  24 - 0x18
      13'h35: dout  = 8'b10001100; //   53 : 140 - 0x8c
      13'h36: dout  = 8'b11000100; //   54 : 196 - 0xc4
      13'h37: dout  = 8'b11111100; //   55 : 252 - 0xfc
      13'h38: dout  = 8'b11110110; //   56 : 246 - 0xf6
      13'h39: dout  = 8'b11110000; //   57 : 240 - 0xf0
      13'h3A: dout  = 8'b00111000; //   58 :  56 - 0x38
      13'h3B: dout  = 8'b11010000; //   59 : 208 - 0xd0
      13'h3C: dout  = 8'b11100000; //   60 : 224 - 0xe0
      13'h3D: dout  = 8'b01110000; //   61 : 112 - 0x70
      13'h3E: dout  = 8'b10111000; //   62 : 184 - 0xb8
      13'h3F: dout  = 8'b01000000; //   63 :  64 - 0x40
      13'h40: dout  = 8'b00100011; //   64 :  35 - 0x23 -- Sprite 0x4
      13'h41: dout  = 8'b00100011; //   65 :  35 - 0x23
      13'h42: dout  = 8'b00100001; //   66 :  33 - 0x21
      13'h43: dout  = 8'b00100000; //   67 :  32 - 0x20
      13'h44: dout  = 8'b00010011; //   68 :  19 - 0x13
      13'h45: dout  = 8'b00001100; //   69 :  12 - 0xc
      13'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      13'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      13'h48: dout  = 8'b00011100; //   72 :  28 - 0x1c
      13'h49: dout  = 8'b00011100; //   73 :  28 - 0x1c
      13'h4A: dout  = 8'b00011110; //   74 :  30 - 0x1e
      13'h4B: dout  = 8'b00011111; //   75 :  31 - 0x1f
      13'h4C: dout  = 8'b00001100; //   76 :  12 - 0xc
      13'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      13'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      13'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      13'h50: dout  = 8'b11111100; //   80 : 252 - 0xfc -- Sprite 0x5
      13'h51: dout  = 8'b11111100; //   81 : 252 - 0xfc
      13'h52: dout  = 8'b11111100; //   82 : 252 - 0xfc
      13'h53: dout  = 8'b11111100; //   83 : 252 - 0xfc
      13'h54: dout  = 8'b10010000; //   84 : 144 - 0x90
      13'h55: dout  = 8'b10010000; //   85 : 144 - 0x90
      13'h56: dout  = 8'b10001000; //   86 : 136 - 0x88
      13'h57: dout  = 8'b11111000; //   87 : 248 - 0xf8
      13'h58: dout  = 8'b10101000; //   88 : 168 - 0xa8
      13'h59: dout  = 8'b01010000; //   89 :  80 - 0x50
      13'h5A: dout  = 8'b10101000; //   90 : 168 - 0xa8
      13'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      13'h5C: dout  = 8'b01100000; //   92 :  96 - 0x60
      13'h5D: dout  = 8'b01100000; //   93 :  96 - 0x60
      13'h5E: dout  = 8'b01110000; //   94 : 112 - 0x70
      13'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      13'h60: dout  = 8'b00100011; //   96 :  35 - 0x23 -- Sprite 0x6
      13'h61: dout  = 8'b00100011; //   97 :  35 - 0x23
      13'h62: dout  = 8'b00100001; //   98 :  33 - 0x21
      13'h63: dout  = 8'b00100000; //   99 :  32 - 0x20
      13'h64: dout  = 8'b00010011; //  100 :  19 - 0x13
      13'h65: dout  = 8'b00001101; //  101 :  13 - 0xd
      13'h66: dout  = 8'b00000010; //  102 :   2 - 0x2
      13'h67: dout  = 8'b00000001; //  103 :   1 - 0x1
      13'h68: dout  = 8'b00011100; //  104 :  28 - 0x1c
      13'h69: dout  = 8'b00011100; //  105 :  28 - 0x1c
      13'h6A: dout  = 8'b00011110; //  106 :  30 - 0x1e
      13'h6B: dout  = 8'b00011111; //  107 :  31 - 0x1f
      13'h6C: dout  = 8'b00001100; //  108 :  12 - 0xc
      13'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      13'h6E: dout  = 8'b00000001; //  110 :   1 - 0x1
      13'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      13'h70: dout  = 8'b11111100; //  112 : 252 - 0xfc -- Sprite 0x7
      13'h71: dout  = 8'b11111100; //  113 : 252 - 0xfc
      13'h72: dout  = 8'b11111100; //  114 : 252 - 0xfc
      13'h73: dout  = 8'b11111100; //  115 : 252 - 0xfc
      13'h74: dout  = 8'b10100100; //  116 : 164 - 0xa4
      13'h75: dout  = 8'b00100100; //  117 :  36 - 0x24
      13'h76: dout  = 8'b01010010; //  118 :  82 - 0x52
      13'h77: dout  = 8'b11101110; //  119 : 238 - 0xee
      13'h78: dout  = 8'b10101000; //  120 : 168 - 0xa8
      13'h79: dout  = 8'b01010000; //  121 :  80 - 0x50
      13'h7A: dout  = 8'b10101000; //  122 : 168 - 0xa8
      13'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      13'h7C: dout  = 8'b01011000; //  124 :  88 - 0x58
      13'h7D: dout  = 8'b11011000; //  125 : 216 - 0xd8
      13'h7E: dout  = 8'b10001100; //  126 : 140 - 0x8c
      13'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout  = 8'b00100011; //  128 :  35 - 0x23 -- Sprite 0x8
      13'h81: dout  = 8'b00100011; //  129 :  35 - 0x23
      13'h82: dout  = 8'b00100001; //  130 :  33 - 0x21
      13'h83: dout  = 8'b00100000; //  131 :  32 - 0x20
      13'h84: dout  = 8'b00010011; //  132 :  19 - 0x13
      13'h85: dout  = 8'b00001101; //  133 :  13 - 0xd
      13'h86: dout  = 8'b00000001; //  134 :   1 - 0x1
      13'h87: dout  = 8'b00000001; //  135 :   1 - 0x1
      13'h88: dout  = 8'b00011100; //  136 :  28 - 0x1c
      13'h89: dout  = 8'b00011100; //  137 :  28 - 0x1c
      13'h8A: dout  = 8'b00011110; //  138 :  30 - 0x1e
      13'h8B: dout  = 8'b00011111; //  139 :  31 - 0x1f
      13'h8C: dout  = 8'b00001100; //  140 :  12 - 0xc
      13'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      13'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      13'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      13'h90: dout  = 8'b11111110; //  144 : 254 - 0xfe -- Sprite 0x9
      13'h91: dout  = 8'b11111110; //  145 : 254 - 0xfe
      13'h92: dout  = 8'b11111110; //  146 : 254 - 0xfe
      13'h93: dout  = 8'b11111111; //  147 : 255 - 0xff
      13'h94: dout  = 8'b10010001; //  148 : 145 - 0x91
      13'h95: dout  = 8'b00101111; //  149 :  47 - 0x2f
      13'h96: dout  = 8'b01000000; //  150 :  64 - 0x40
      13'h97: dout  = 8'b11100000; //  151 : 224 - 0xe0
      13'h98: dout  = 8'b10101000; //  152 : 168 - 0xa8
      13'h99: dout  = 8'b01010100; //  153 :  84 - 0x54
      13'h9A: dout  = 8'b10101000; //  154 : 168 - 0xa8
      13'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      13'h9C: dout  = 8'b01101110; //  156 : 110 - 0x6e
      13'h9D: dout  = 8'b11000000; //  157 : 192 - 0xc0
      13'h9E: dout  = 8'b10000000; //  158 : 128 - 0x80
      13'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout  = 8'b00100011; //  160 :  35 - 0x23 -- Sprite 0xa
      13'hA1: dout  = 8'b00100011; //  161 :  35 - 0x23
      13'hA2: dout  = 8'b00100001; //  162 :  33 - 0x21
      13'hA3: dout  = 8'b00100000; //  163 :  32 - 0x20
      13'hA4: dout  = 8'b00010011; //  164 :  19 - 0x13
      13'hA5: dout  = 8'b00001110; //  165 :  14 - 0xe
      13'hA6: dout  = 8'b00000001; //  166 :   1 - 0x1
      13'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      13'hA8: dout  = 8'b00011100; //  168 :  28 - 0x1c
      13'hA9: dout  = 8'b00011100; //  169 :  28 - 0x1c
      13'hAA: dout  = 8'b00011110; //  170 :  30 - 0x1e
      13'hAB: dout  = 8'b00011111; //  171 :  31 - 0x1f
      13'hAC: dout  = 8'b00001100; //  172 :  12 - 0xc
      13'hAD: dout  = 8'b00000001; //  173 :   1 - 0x1
      13'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      13'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      13'hB0: dout  = 8'b11111110; //  176 : 254 - 0xfe -- Sprite 0xb
      13'hB1: dout  = 8'b11111110; //  177 : 254 - 0xfe
      13'hB2: dout  = 8'b11111110; //  178 : 254 - 0xfe
      13'hB3: dout  = 8'b11111100; //  179 : 252 - 0xfc
      13'hB4: dout  = 8'b00100100; //  180 :  36 - 0x24
      13'hB5: dout  = 8'b00100010; //  181 :  34 - 0x22
      13'hB6: dout  = 8'b11010010; //  182 : 210 - 0xd2
      13'hB7: dout  = 8'b00001111; //  183 :  15 - 0xf
      13'hB8: dout  = 8'b10101000; //  184 : 168 - 0xa8
      13'hB9: dout  = 8'b01010100; //  185 :  84 - 0x54
      13'hBA: dout  = 8'b10101000; //  186 : 168 - 0xa8
      13'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      13'hBC: dout  = 8'b11011000; //  188 : 216 - 0xd8
      13'hBD: dout  = 8'b11011100; //  189 : 220 - 0xdc
      13'hBE: dout  = 8'b00001100; //  190 :  12 - 0xc
      13'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout  = 8'b01111111; //  192 : 127 - 0x7f -- Sprite 0xc
      13'hC1: dout  = 8'b01111110; //  193 : 126 - 0x7e
      13'hC2: dout  = 8'b11111100; //  194 : 252 - 0xfc
      13'hC3: dout  = 8'b00000010; //  195 :   2 - 0x2
      13'hC4: dout  = 8'b00000100; //  196 :   4 - 0x4
      13'hC5: dout  = 8'b11111100; //  197 : 252 - 0xfc
      13'hC6: dout  = 8'b11111100; //  198 : 252 - 0xfc
      13'hC7: dout  = 8'b11111110; //  199 : 254 - 0xfe
      13'hC8: dout  = 8'b11110110; //  200 : 246 - 0xf6
      13'hC9: dout  = 8'b11110000; //  201 : 240 - 0xf0
      13'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      13'hCB: dout  = 8'b11111100; //  203 : 252 - 0xfc
      13'hCC: dout  = 8'b11111000; //  204 : 248 - 0xf8
      13'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      13'hCE: dout  = 8'b10101000; //  206 : 168 - 0xa8
      13'hCF: dout  = 8'b01010100; //  207 :  84 - 0x54
      13'hD0: dout  = 8'b01000101; //  208 :  69 - 0x45 -- Sprite 0xd
      13'hD1: dout  = 8'b10000111; //  209 : 135 - 0x87
      13'hD2: dout  = 8'b10000011; //  210 : 131 - 0x83
      13'hD3: dout  = 8'b10000010; //  211 : 130 - 0x82
      13'hD4: dout  = 8'b10000010; //  212 : 130 - 0x82
      13'hD5: dout  = 8'b10000100; //  213 : 132 - 0x84
      13'hD6: dout  = 8'b01000100; //  214 :  68 - 0x44
      13'hD7: dout  = 8'b00100100; //  215 :  36 - 0x24
      13'hD8: dout  = 8'b00111000; //  216 :  56 - 0x38
      13'hD9: dout  = 8'b01111000; //  217 : 120 - 0x78
      13'hDA: dout  = 8'b01111100; //  218 : 124 - 0x7c
      13'hDB: dout  = 8'b01111101; //  219 : 125 - 0x7d
      13'hDC: dout  = 8'b01111101; //  220 : 125 - 0x7d
      13'hDD: dout  = 8'b01111011; //  221 : 123 - 0x7b
      13'hDE: dout  = 8'b00111011; //  222 :  59 - 0x3b
      13'hDF: dout  = 8'b00011011; //  223 :  27 - 0x1b
      13'hE0: dout  = 8'b01111111; //  224 : 127 - 0x7f -- Sprite 0xe
      13'hE1: dout  = 8'b01111110; //  225 : 126 - 0x7e
      13'hE2: dout  = 8'b11111100; //  226 : 252 - 0xfc
      13'hE3: dout  = 8'b11111000; //  227 : 248 - 0xf8
      13'hE4: dout  = 8'b01111000; //  228 : 120 - 0x78
      13'hE5: dout  = 8'b01111100; //  229 : 124 - 0x7c
      13'hE6: dout  = 8'b11111100; //  230 : 252 - 0xfc
      13'hE7: dout  = 8'b11111110; //  231 : 254 - 0xfe
      13'hE8: dout  = 8'b11110110; //  232 : 246 - 0xf6
      13'hE9: dout  = 8'b11110000; //  233 : 240 - 0xf0
      13'hEA: dout  = 8'b01111000; //  234 : 120 - 0x78
      13'hEB: dout  = 8'b01110000; //  235 : 112 - 0x70
      13'hEC: dout  = 8'b10100000; //  236 : 160 - 0xa0
      13'hED: dout  = 8'b10010000; //  237 : 144 - 0x90
      13'hEE: dout  = 8'b00101000; //  238 :  40 - 0x28
      13'hEF: dout  = 8'b01010100; //  239 :  84 - 0x54
      13'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      13'hF1: dout  = 8'b00001111; //  241 :  15 - 0xf
      13'hF2: dout  = 8'b00000100; //  242 :   4 - 0x4
      13'hF3: dout  = 8'b00000011; //  243 :   3 - 0x3
      13'hF4: dout  = 8'b00000011; //  244 :   3 - 0x3
      13'hF5: dout  = 8'b00000011; //  245 :   3 - 0x3
      13'hF6: dout  = 8'b00000100; //  246 :   4 - 0x4
      13'hF7: dout  = 8'b00000010; //  247 :   2 - 0x2
      13'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0
      13'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      13'hFA: dout  = 8'b00000011; //  250 :   3 - 0x3
      13'hFB: dout  = 8'b00000001; //  251 :   1 - 0x1
      13'hFC: dout  = 8'b00000001; //  252 :   1 - 0x1
      13'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      13'hFE: dout  = 8'b00000011; //  254 :   3 - 0x3
      13'hFF: dout  = 8'b00000001; //  255 :   1 - 0x1
      13'h100: dout  = 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x10
      13'h101: dout  = 8'b00001100; //  257 :  12 - 0xc
      13'h102: dout  = 8'b00010000; //  258 :  16 - 0x10
      13'h103: dout  = 8'b00010000; //  259 :  16 - 0x10
      13'h104: dout  = 8'b00010000; //  260 :  16 - 0x10
      13'h105: dout  = 8'b00100000; //  261 :  32 - 0x20
      13'h106: dout  = 8'b00100000; //  262 :  32 - 0x20
      13'h107: dout  = 8'b00100001; //  263 :  33 - 0x21
      13'h108: dout  = 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout  = 8'b00000011; //  265 :   3 - 0x3
      13'h10A: dout  = 8'b00001111; //  266 :  15 - 0xf
      13'h10B: dout  = 8'b00001111; //  267 :  15 - 0xf
      13'h10C: dout  = 8'b00001111; //  268 :  15 - 0xf
      13'h10D: dout  = 8'b00011111; //  269 :  31 - 0x1f
      13'h10E: dout  = 8'b00011111; //  270 :  31 - 0x1f
      13'h10F: dout  = 8'b00011110; //  271 :  30 - 0x1e
      13'h110: dout  = 8'b11111111; //  272 : 255 - 0xff -- Sprite 0x11
      13'h111: dout  = 8'b01111110; //  273 : 126 - 0x7e
      13'h112: dout  = 8'b01111100; //  274 : 124 - 0x7c
      13'h113: dout  = 8'b01111000; //  275 : 120 - 0x78
      13'h114: dout  = 8'b01011000; //  276 :  88 - 0x58
      13'h115: dout  = 8'b10001100; //  277 : 140 - 0x8c
      13'h116: dout  = 8'b11000100; //  278 : 196 - 0xc4
      13'h117: dout  = 8'b11111100; //  279 : 252 - 0xfc
      13'h118: dout  = 8'b00110110; //  280 :  54 - 0x36
      13'h119: dout  = 8'b10110000; //  281 : 176 - 0xb0
      13'h11A: dout  = 8'b10111000; //  282 : 184 - 0xb8
      13'h11B: dout  = 8'b10010000; //  283 : 144 - 0x90
      13'h11C: dout  = 8'b10100000; //  284 : 160 - 0xa0
      13'h11D: dout  = 8'b01110000; //  285 : 112 - 0x70
      13'h11E: dout  = 8'b00111000; //  286 :  56 - 0x38
      13'h11F: dout  = 8'b01000000; //  287 :  64 - 0x40
      13'h120: dout  = 8'b00100011; //  288 :  35 - 0x23 -- Sprite 0x12
      13'h121: dout  = 8'b00100011; //  289 :  35 - 0x23
      13'h122: dout  = 8'b00100001; //  290 :  33 - 0x21
      13'h123: dout  = 8'b00100000; //  291 :  32 - 0x20
      13'h124: dout  = 8'b00010011; //  292 :  19 - 0x13
      13'h125: dout  = 8'b00001100; //  293 :  12 - 0xc
      13'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      13'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      13'h128: dout  = 8'b00011100; //  296 :  28 - 0x1c
      13'h129: dout  = 8'b00011100; //  297 :  28 - 0x1c
      13'h12A: dout  = 8'b00011110; //  298 :  30 - 0x1e
      13'h12B: dout  = 8'b00011111; //  299 :  31 - 0x1f
      13'h12C: dout  = 8'b00001100; //  300 :  12 - 0xc
      13'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      13'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      13'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      13'h130: dout  = 8'b00000001; //  304 :   1 - 0x1 -- Sprite 0x13
      13'h131: dout  = 8'b00000001; //  305 :   1 - 0x1
      13'h132: dout  = 8'b00000011; //  306 :   3 - 0x3
      13'h133: dout  = 8'b00000100; //  307 :   4 - 0x4
      13'h134: dout  = 8'b00001000; //  308 :   8 - 0x8
      13'h135: dout  = 8'b00010000; //  309 :  16 - 0x10
      13'h136: dout  = 8'b00010000; //  310 :  16 - 0x10
      13'h137: dout  = 8'b00100000; //  311 :  32 - 0x20
      13'h138: dout  = 8'b00000000; //  312 :   0 - 0x0
      13'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      13'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      13'h13B: dout  = 8'b00000011; //  315 :   3 - 0x3
      13'h13C: dout  = 8'b00000111; //  316 :   7 - 0x7
      13'h13D: dout  = 8'b00001111; //  317 :  15 - 0xf
      13'h13E: dout  = 8'b00001111; //  318 :  15 - 0xf
      13'h13F: dout  = 8'b00011111; //  319 :  31 - 0x1f
      13'h140: dout  = 8'b01111111; //  320 : 127 - 0x7f -- Sprite 0x14
      13'h141: dout  = 8'b11111110; //  321 : 254 - 0xfe
      13'h142: dout  = 8'b00000110; //  322 :   6 - 0x6
      13'h143: dout  = 8'b00000001; //  323 :   1 - 0x1
      13'h144: dout  = 8'b00000001; //  324 :   1 - 0x1
      13'h145: dout  = 8'b00000001; //  325 :   1 - 0x1
      13'h146: dout  = 8'b00000111; //  326 :   7 - 0x7
      13'h147: dout  = 8'b11111110; //  327 : 254 - 0xfe
      13'h148: dout  = 8'b11110110; //  328 : 246 - 0xf6
      13'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      13'h14A: dout  = 8'b11111000; //  330 : 248 - 0xf8
      13'h14B: dout  = 8'b11111110; //  331 : 254 - 0xfe
      13'h14C: dout  = 8'b11111110; //  332 : 254 - 0xfe
      13'h14D: dout  = 8'b11111110; //  333 : 254 - 0xfe
      13'h14E: dout  = 8'b11111000; //  334 : 248 - 0xf8
      13'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout  = 8'b00000101; //  336 :   5 - 0x5 -- Sprite 0x15
      13'h151: dout  = 8'b00000101; //  337 :   5 - 0x5
      13'h152: dout  = 8'b00000111; //  338 :   7 - 0x7
      13'h153: dout  = 8'b00000100; //  339 :   4 - 0x4
      13'h154: dout  = 8'b00000100; //  340 :   4 - 0x4
      13'h155: dout  = 8'b00001111; //  341 :  15 - 0xf
      13'h156: dout  = 8'b00110000; //  342 :  48 - 0x30
      13'h157: dout  = 8'b01000000; //  343 :  64 - 0x40
      13'h158: dout  = 8'b00000011; //  344 :   3 - 0x3
      13'h159: dout  = 8'b00000011; //  345 :   3 - 0x3
      13'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      13'h15B: dout  = 8'b00000011; //  347 :   3 - 0x3
      13'h15C: dout  = 8'b00000011; //  348 :   3 - 0x3
      13'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      13'h15E: dout  = 8'b00001111; //  350 :  15 - 0xf
      13'h15F: dout  = 8'b00111111; //  351 :  63 - 0x3f
      13'h160: dout  = 8'b11111100; //  352 : 252 - 0xfc -- Sprite 0x16
      13'h161: dout  = 8'b11111000; //  353 : 248 - 0xf8
      13'h162: dout  = 8'b11110000; //  354 : 240 - 0xf0
      13'h163: dout  = 8'b11100000; //  355 : 224 - 0xe0
      13'h164: dout  = 8'b01100000; //  356 :  96 - 0x60
      13'h165: dout  = 8'b11110000; //  357 : 240 - 0xf0
      13'h166: dout  = 8'b00011100; //  358 :  28 - 0x1c
      13'h167: dout  = 8'b00000010; //  359 :   2 - 0x2
      13'h168: dout  = 8'b11011000; //  360 : 216 - 0xd8
      13'h169: dout  = 8'b11000000; //  361 : 192 - 0xc0
      13'h16A: dout  = 8'b11100000; //  362 : 224 - 0xe0
      13'h16B: dout  = 8'b01000000; //  363 :  64 - 0x40
      13'h16C: dout  = 8'b10000000; //  364 : 128 - 0x80
      13'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      13'h16E: dout  = 8'b11100000; //  366 : 224 - 0xe0
      13'h16F: dout  = 8'b11111100; //  367 : 252 - 0xfc
      13'h170: dout  = 8'b10000000; //  368 : 128 - 0x80 -- Sprite 0x17
      13'h171: dout  = 8'b10000000; //  369 : 128 - 0x80
      13'h172: dout  = 8'b10000000; //  370 : 128 - 0x80
      13'h173: dout  = 8'b10000011; //  371 : 131 - 0x83
      13'h174: dout  = 8'b01001111; //  372 :  79 - 0x4f
      13'h175: dout  = 8'b00110010; //  373 :  50 - 0x32
      13'h176: dout  = 8'b00000010; //  374 :   2 - 0x2
      13'h177: dout  = 8'b00000011; //  375 :   3 - 0x3
      13'h178: dout  = 8'b01111111; //  376 : 127 - 0x7f
      13'h179: dout  = 8'b01111111; //  377 : 127 - 0x7f
      13'h17A: dout  = 8'b01111111; //  378 : 127 - 0x7f
      13'h17B: dout  = 8'b01111100; //  379 : 124 - 0x7c
      13'h17C: dout  = 8'b00110000; //  380 :  48 - 0x30
      13'h17D: dout  = 8'b00000001; //  381 :   1 - 0x1
      13'h17E: dout  = 8'b00000001; //  382 :   1 - 0x1
      13'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout  = 8'b00000010; //  384 :   2 - 0x2 -- Sprite 0x18
      13'h181: dout  = 8'b00000001; //  385 :   1 - 0x1
      13'h182: dout  = 8'b00000010; //  386 :   2 - 0x2
      13'h183: dout  = 8'b11111100; //  387 : 252 - 0xfc
      13'h184: dout  = 8'b11000000; //  388 : 192 - 0xc0
      13'h185: dout  = 8'b01000000; //  389 :  64 - 0x40
      13'h186: dout  = 8'b00100000; //  390 :  32 - 0x20
      13'h187: dout  = 8'b11100000; //  391 : 224 - 0xe0
      13'h188: dout  = 8'b11111100; //  392 : 252 - 0xfc
      13'h189: dout  = 8'b11111110; //  393 : 254 - 0xfe
      13'h18A: dout  = 8'b11111100; //  394 : 252 - 0xfc
      13'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      13'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      13'h18D: dout  = 8'b10000000; //  397 : 128 - 0x80
      13'h18E: dout  = 8'b11000000; //  398 : 192 - 0xc0
      13'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      13'h190: dout  = 8'b00001011; //  400 :  11 - 0xb -- Sprite 0x19
      13'h191: dout  = 8'b00001011; //  401 :  11 - 0xb
      13'h192: dout  = 8'b00001111; //  402 :  15 - 0xf
      13'h193: dout  = 8'b00001001; //  403 :   9 - 0x9
      13'h194: dout  = 8'b00001000; //  404 :   8 - 0x8
      13'h195: dout  = 8'b00001001; //  405 :   9 - 0x9
      13'h196: dout  = 8'b00001111; //  406 :  15 - 0xf
      13'h197: dout  = 8'b00110000; //  407 :  48 - 0x30
      13'h198: dout  = 8'b00000111; //  408 :   7 - 0x7
      13'h199: dout  = 8'b00000111; //  409 :   7 - 0x7
      13'h19A: dout  = 8'b00000001; //  410 :   1 - 0x1
      13'h19B: dout  = 8'b00000110; //  411 :   6 - 0x6
      13'h19C: dout  = 8'b00000111; //  412 :   7 - 0x7
      13'h19D: dout  = 8'b00000110; //  413 :   6 - 0x6
      13'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout  = 8'b00001111; //  415 :  15 - 0xf
      13'h1A0: dout  = 8'b11111000; //  416 : 248 - 0xf8 -- Sprite 0x1a
      13'h1A1: dout  = 8'b11110000; //  417 : 240 - 0xf0
      13'h1A2: dout  = 8'b11100000; //  418 : 224 - 0xe0
      13'h1A3: dout  = 8'b11000000; //  419 : 192 - 0xc0
      13'h1A4: dout  = 8'b11000000; //  420 : 192 - 0xc0
      13'h1A5: dout  = 8'b11000000; //  421 : 192 - 0xc0
      13'h1A6: dout  = 8'b11111000; //  422 : 248 - 0xf8
      13'h1A7: dout  = 8'b00011111; //  423 :  31 - 0x1f
      13'h1A8: dout  = 8'b10110000; //  424 : 176 - 0xb0
      13'h1A9: dout  = 8'b10000000; //  425 : 128 - 0x80
      13'h1AA: dout  = 8'b11000000; //  426 : 192 - 0xc0
      13'h1AB: dout  = 8'b10000000; //  427 : 128 - 0x80
      13'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      13'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      13'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      13'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      13'h1B0: dout  = 8'b01000000; //  432 :  64 - 0x40 -- Sprite 0x1b
      13'h1B1: dout  = 8'b01000000; //  433 :  64 - 0x40
      13'h1B2: dout  = 8'b10000000; //  434 : 128 - 0x80
      13'h1B3: dout  = 8'b10000000; //  435 : 128 - 0x80
      13'h1B4: dout  = 8'b01000000; //  436 :  64 - 0x40
      13'h1B5: dout  = 8'b00111111; //  437 :  63 - 0x3f
      13'h1B6: dout  = 8'b00000100; //  438 :   4 - 0x4
      13'h1B7: dout  = 8'b00000111; //  439 :   7 - 0x7
      13'h1B8: dout  = 8'b00111111; //  440 :  63 - 0x3f
      13'h1B9: dout  = 8'b00111111; //  441 :  63 - 0x3f
      13'h1BA: dout  = 8'b01111111; //  442 : 127 - 0x7f
      13'h1BB: dout  = 8'b01111111; //  443 : 127 - 0x7f
      13'h1BC: dout  = 8'b00111111; //  444 :  63 - 0x3f
      13'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      13'h1BE: dout  = 8'b00000011; //  446 :   3 - 0x3
      13'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      13'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x1c
      13'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      13'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      13'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      13'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      13'h1C5: dout  = 8'b11111111; //  453 : 255 - 0xff
      13'h1C6: dout  = 8'b01000000; //  454 :  64 - 0x40
      13'h1C7: dout  = 8'b11000000; //  455 : 192 - 0xc0
      13'h1C8: dout  = 8'b11111111; //  456 : 255 - 0xff
      13'h1C9: dout  = 8'b11111111; //  457 : 255 - 0xff
      13'h1CA: dout  = 8'b11111111; //  458 : 255 - 0xff
      13'h1CB: dout  = 8'b11111111; //  459 : 255 - 0xff
      13'h1CC: dout  = 8'b11111111; //  460 : 255 - 0xff
      13'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      13'h1CE: dout  = 8'b10000000; //  462 : 128 - 0x80
      13'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      13'h1D0: dout  = 8'b11000000; //  464 : 192 - 0xc0 -- Sprite 0x1d
      13'h1D1: dout  = 8'b00100000; //  465 :  32 - 0x20
      13'h1D2: dout  = 8'b00100000; //  466 :  32 - 0x20
      13'h1D3: dout  = 8'b00100000; //  467 :  32 - 0x20
      13'h1D4: dout  = 8'b01000000; //  468 :  64 - 0x40
      13'h1D5: dout  = 8'b10000000; //  469 : 128 - 0x80
      13'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      13'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      13'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0
      13'h1D9: dout  = 8'b11000000; //  473 : 192 - 0xc0
      13'h1DA: dout  = 8'b11000000; //  474 : 192 - 0xc0
      13'h1DB: dout  = 8'b11000000; //  475 : 192 - 0xc0
      13'h1DC: dout  = 8'b10000000; //  476 : 128 - 0x80
      13'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      13'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout  = 8'b01111111; //  480 : 127 - 0x7f -- Sprite 0x1e
      13'h1E1: dout  = 8'b01100010; //  481 :  98 - 0x62
      13'h1E2: dout  = 8'b11000100; //  482 : 196 - 0xc4
      13'h1E3: dout  = 8'b00011000; //  483 :  24 - 0x18
      13'h1E4: dout  = 8'b00111100; //  484 :  60 - 0x3c
      13'h1E5: dout  = 8'b11111110; //  485 : 254 - 0xfe
      13'h1E6: dout  = 8'b11111110; //  486 : 254 - 0xfe
      13'h1E7: dout  = 8'b11111110; //  487 : 254 - 0xfe
      13'h1E8: dout  = 8'b11100000; //  488 : 224 - 0xe0
      13'h1E9: dout  = 8'b10011100; //  489 : 156 - 0x9c
      13'h1EA: dout  = 8'b00111000; //  490 :  56 - 0x38
      13'h1EB: dout  = 8'b11100000; //  491 : 224 - 0xe0
      13'h1EC: dout  = 8'b11001000; //  492 : 200 - 0xc8
      13'h1ED: dout  = 8'b00010100; //  493 :  20 - 0x14
      13'h1EE: dout  = 8'b10101000; //  494 : 168 - 0xa8
      13'h1EF: dout  = 8'b01010100; //  495 :  84 - 0x54
      13'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x1f
      13'h1F1: dout  = 8'b00111000; //  497 :  56 - 0x38
      13'h1F2: dout  = 8'b11000110; //  498 : 198 - 0xc6
      13'h1F3: dout  = 8'b11001011; //  499 : 203 - 0xcb
      13'h1F4: dout  = 8'b11011100; //  500 : 220 - 0xdc
      13'h1F5: dout  = 8'b00111010; //  501 :  58 - 0x3a
      13'h1F6: dout  = 8'b10011010; //  502 : 154 - 0x9a
      13'h1F7: dout  = 8'b11100001; //  503 : 225 - 0xe1
      13'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0
      13'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      13'h1FA: dout  = 8'b00111000; //  506 :  56 - 0x38
      13'h1FB: dout  = 8'b10110100; //  507 : 180 - 0xb4
      13'h1FC: dout  = 8'b10101000; //  508 : 168 - 0xa8
      13'h1FD: dout  = 8'b11010100; //  509 : 212 - 0xd4
      13'h1FE: dout  = 8'b01110100; //  510 : 116 - 0x74
      13'h1FF: dout  = 8'b00011110; //  511 :  30 - 0x1e
      13'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      13'h201: dout  = 8'b00011100; //  513 :  28 - 0x1c
      13'h202: dout  = 8'b00010011; //  514 :  19 - 0x13
      13'h203: dout  = 8'b00001000; //  515 :   8 - 0x8
      13'h204: dout  = 8'b00010000; //  516 :  16 - 0x10
      13'h205: dout  = 8'b00001000; //  517 :   8 - 0x8
      13'h206: dout  = 8'b00010000; //  518 :  16 - 0x10
      13'h207: dout  = 8'b00010000; //  519 :  16 - 0x10
      13'h208: dout  = 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      13'h20A: dout  = 8'b00001100; //  522 :  12 - 0xc
      13'h20B: dout  = 8'b00000111; //  523 :   7 - 0x7
      13'h20C: dout  = 8'b00001111; //  524 :  15 - 0xf
      13'h20D: dout  = 8'b00000111; //  525 :   7 - 0x7
      13'h20E: dout  = 8'b00001111; //  526 :  15 - 0xf
      13'h20F: dout  = 8'b00001111; //  527 :  15 - 0xf
      13'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      13'h211: dout  = 8'b00111000; //  529 :  56 - 0x38
      13'h212: dout  = 8'b11001000; //  530 : 200 - 0xc8
      13'h213: dout  = 8'b00010000; //  531 :  16 - 0x10
      13'h214: dout  = 8'b00001000; //  532 :   8 - 0x8
      13'h215: dout  = 8'b00010000; //  533 :  16 - 0x10
      13'h216: dout  = 8'b00001000; //  534 :   8 - 0x8
      13'h217: dout  = 8'b00001000; //  535 :   8 - 0x8
      13'h218: dout  = 8'b00000000; //  536 :   0 - 0x0
      13'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      13'h21A: dout  = 8'b00110000; //  538 :  48 - 0x30
      13'h21B: dout  = 8'b11100000; //  539 : 224 - 0xe0
      13'h21C: dout  = 8'b11110000; //  540 : 240 - 0xf0
      13'h21D: dout  = 8'b11100000; //  541 : 224 - 0xe0
      13'h21E: dout  = 8'b11110000; //  542 : 240 - 0xf0
      13'h21F: dout  = 8'b11110000; //  543 : 240 - 0xf0
      13'h220: dout  = 8'b00001000; //  544 :   8 - 0x8 -- Sprite 0x22
      13'h221: dout  = 8'b00011100; //  545 :  28 - 0x1c
      13'h222: dout  = 8'b00100111; //  546 :  39 - 0x27
      13'h223: dout  = 8'b00101111; //  547 :  47 - 0x2f
      13'h224: dout  = 8'b00011111; //  548 :  31 - 0x1f
      13'h225: dout  = 8'b00001111; //  549 :  15 - 0xf
      13'h226: dout  = 8'b00001111; //  550 :  15 - 0xf
      13'h227: dout  = 8'b00001111; //  551 :  15 - 0xf
      13'h228: dout  = 8'b00000111; //  552 :   7 - 0x7
      13'h229: dout  = 8'b00000011; //  553 :   3 - 0x3
      13'h22A: dout  = 8'b00011000; //  554 :  24 - 0x18
      13'h22B: dout  = 8'b00010101; //  555 :  21 - 0x15
      13'h22C: dout  = 8'b00000010; //  556 :   2 - 0x2
      13'h22D: dout  = 8'b00000101; //  557 :   5 - 0x5
      13'h22E: dout  = 8'b00000010; //  558 :   2 - 0x2
      13'h22F: dout  = 8'b00000100; //  559 :   4 - 0x4
      13'h230: dout  = 8'b00010000; //  560 :  16 - 0x10 -- Sprite 0x23
      13'h231: dout  = 8'b00111100; //  561 :  60 - 0x3c
      13'h232: dout  = 8'b11000010; //  562 : 194 - 0xc2
      13'h233: dout  = 8'b10000010; //  563 : 130 - 0x82
      13'h234: dout  = 8'b10000010; //  564 : 130 - 0x82
      13'h235: dout  = 8'b10000010; //  565 : 130 - 0x82
      13'h236: dout  = 8'b00010010; //  566 :  18 - 0x12
      13'h237: dout  = 8'b00011100; //  567 :  28 - 0x1c
      13'h238: dout  = 8'b11100000; //  568 : 224 - 0xe0
      13'h239: dout  = 8'b11000000; //  569 : 192 - 0xc0
      13'h23A: dout  = 8'b00111100; //  570 :  60 - 0x3c
      13'h23B: dout  = 8'b01111100; //  571 : 124 - 0x7c
      13'h23C: dout  = 8'b01111100; //  572 : 124 - 0x7c
      13'h23D: dout  = 8'b01111100; //  573 : 124 - 0x7c
      13'h23E: dout  = 8'b11101100; //  574 : 236 - 0xec
      13'h23F: dout  = 8'b11100000; //  575 : 224 - 0xe0
      13'h240: dout  = 8'b00001111; //  576 :  15 - 0xf -- Sprite 0x24
      13'h241: dout  = 8'b00001110; //  577 :  14 - 0xe
      13'h242: dout  = 8'b00010100; //  578 :  20 - 0x14
      13'h243: dout  = 8'b00010100; //  579 :  20 - 0x14
      13'h244: dout  = 8'b00010010; //  580 :  18 - 0x12
      13'h245: dout  = 8'b00100101; //  581 :  37 - 0x25
      13'h246: dout  = 8'b01000100; //  582 :  68 - 0x44
      13'h247: dout  = 8'b00111000; //  583 :  56 - 0x38
      13'h248: dout  = 8'b00000010; //  584 :   2 - 0x2
      13'h249: dout  = 8'b00000101; //  585 :   5 - 0x5
      13'h24A: dout  = 8'b00001011; //  586 :  11 - 0xb
      13'h24B: dout  = 8'b00001011; //  587 :  11 - 0xb
      13'h24C: dout  = 8'b00001101; //  588 :  13 - 0xd
      13'h24D: dout  = 8'b00011000; //  589 :  24 - 0x18
      13'h24E: dout  = 8'b00111000; //  590 :  56 - 0x38
      13'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout  = 8'b00010000; //  592 :  16 - 0x10 -- Sprite 0x25
      13'h251: dout  = 8'b00010000; //  593 :  16 - 0x10
      13'h252: dout  = 8'b00010000; //  594 :  16 - 0x10
      13'h253: dout  = 8'b00101100; //  595 :  44 - 0x2c
      13'h254: dout  = 8'b01000100; //  596 :  68 - 0x44
      13'h255: dout  = 8'b11000100; //  597 : 196 - 0xc4
      13'h256: dout  = 8'b00111000; //  598 :  56 - 0x38
      13'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      13'h258: dout  = 8'b11100000; //  600 : 224 - 0xe0
      13'h259: dout  = 8'b11100000; //  601 : 224 - 0xe0
      13'h25A: dout  = 8'b11100000; //  602 : 224 - 0xe0
      13'h25B: dout  = 8'b11010000; //  603 : 208 - 0xd0
      13'h25C: dout  = 8'b10111000; //  604 : 184 - 0xb8
      13'h25D: dout  = 8'b00111000; //  605 :  56 - 0x38
      13'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      13'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      13'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      13'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      13'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      13'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      13'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      13'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      13'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      13'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      13'h268: dout  = 8'b00000000; //  616 :   0 - 0x0
      13'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      13'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      13'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      13'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      13'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      13'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      13'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x27
      13'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      13'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      13'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      13'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      13'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      13'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      13'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      13'h278: dout  = 8'b00000000; //  632 :   0 - 0x0
      13'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      13'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      13'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      13'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      13'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      13'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      13'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      13'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      13'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      13'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      13'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      13'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      13'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      13'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      13'h288: dout  = 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      13'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      13'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      13'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      13'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      13'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      13'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      13'h290: dout  = 8'b00100000; //  656 :  32 - 0x20 -- Sprite 0x29
      13'h291: dout  = 8'b00100000; //  657 :  32 - 0x20
      13'h292: dout  = 8'b00100000; //  658 :  32 - 0x20
      13'h293: dout  = 8'b00100000; //  659 :  32 - 0x20
      13'h294: dout  = 8'b00010011; //  660 :  19 - 0x13
      13'h295: dout  = 8'b00001101; //  661 :  13 - 0xd
      13'h296: dout  = 8'b00000010; //  662 :   2 - 0x2
      13'h297: dout  = 8'b00000001; //  663 :   1 - 0x1
      13'h298: dout  = 8'b00011111; //  664 :  31 - 0x1f
      13'h299: dout  = 8'b00011111; //  665 :  31 - 0x1f
      13'h29A: dout  = 8'b00011111; //  666 :  31 - 0x1f
      13'h29B: dout  = 8'b00011111; //  667 :  31 - 0x1f
      13'h29C: dout  = 8'b00001100; //  668 :  12 - 0xc
      13'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      13'h29E: dout  = 8'b00000001; //  670 :   1 - 0x1
      13'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      13'h2A0: dout  = 8'b00100000; //  672 :  32 - 0x20 -- Sprite 0x2a
      13'h2A1: dout  = 8'b00100000; //  673 :  32 - 0x20
      13'h2A2: dout  = 8'b00100000; //  674 :  32 - 0x20
      13'h2A3: dout  = 8'b00100000; //  675 :  32 - 0x20
      13'h2A4: dout  = 8'b00010011; //  676 :  19 - 0x13
      13'h2A5: dout  = 8'b00001101; //  677 :  13 - 0xd
      13'h2A6: dout  = 8'b00000001; //  678 :   1 - 0x1
      13'h2A7: dout  = 8'b00000001; //  679 :   1 - 0x1
      13'h2A8: dout  = 8'b00011111; //  680 :  31 - 0x1f
      13'h2A9: dout  = 8'b00011111; //  681 :  31 - 0x1f
      13'h2AA: dout  = 8'b00011111; //  682 :  31 - 0x1f
      13'h2AB: dout  = 8'b00011111; //  683 :  31 - 0x1f
      13'h2AC: dout  = 8'b00001100; //  684 :  12 - 0xc
      13'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      13'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      13'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      13'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x2b
      13'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      13'h2B2: dout  = 8'b00000000; //  690 :   0 - 0x0
      13'h2B3: dout  = 8'b00000000; //  691 :   0 - 0x0
      13'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      13'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      13'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      13'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      13'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0
      13'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      13'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      13'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      13'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      13'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      13'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      13'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      13'h2C1: dout  = 8'b00000000; //  705 :   0 - 0x0
      13'h2C2: dout  = 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout  = 8'b00000000; //  707 :   0 - 0x0
      13'h2C4: dout  = 8'b00000000; //  708 :   0 - 0x0
      13'h2C5: dout  = 8'b00000000; //  709 :   0 - 0x0
      13'h2C6: dout  = 8'b00000000; //  710 :   0 - 0x0
      13'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0
      13'h2C9: dout  = 8'b00000000; //  713 :   0 - 0x0
      13'h2CA: dout  = 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      13'h2CC: dout  = 8'b00000000; //  716 :   0 - 0x0
      13'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      13'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      13'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      13'h2D0: dout  = 8'b00111100; //  720 :  60 - 0x3c -- Sprite 0x2d
      13'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      13'h2D2: dout  = 8'b10000001; //  722 : 129 - 0x81
      13'h2D3: dout  = 8'b10011001; //  723 : 153 - 0x99
      13'h2D4: dout  = 8'b10011001; //  724 : 153 - 0x99
      13'h2D5: dout  = 8'b10000001; //  725 : 129 - 0x81
      13'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      13'h2D7: dout  = 8'b00111100; //  727 :  60 - 0x3c
      13'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0
      13'h2D9: dout  = 8'b01111110; //  729 : 126 - 0x7e
      13'h2DA: dout  = 8'b01000010; //  730 :  66 - 0x42
      13'h2DB: dout  = 8'b01000010; //  731 :  66 - 0x42
      13'h2DC: dout  = 8'b01000010; //  732 :  66 - 0x42
      13'h2DD: dout  = 8'b01000010; //  733 :  66 - 0x42
      13'h2DE: dout  = 8'b01111110; //  734 : 126 - 0x7e
      13'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      13'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      13'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      13'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      13'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      13'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      13'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      13'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0
      13'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      13'h2EA: dout  = 8'b00000000; //  746 :   0 - 0x0
      13'h2EB: dout  = 8'b00000000; //  747 :   0 - 0x0
      13'h2EC: dout  = 8'b00000000; //  748 :   0 - 0x0
      13'h2ED: dout  = 8'b00000000; //  749 :   0 - 0x0
      13'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      13'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      13'h2F0: dout  = 8'b10011111; //  752 : 159 - 0x9f -- Sprite 0x2f
      13'h2F1: dout  = 8'b10011110; //  753 : 158 - 0x9e
      13'h2F2: dout  = 8'b10011100; //  754 : 156 - 0x9c
      13'h2F3: dout  = 8'b00011000; //  755 :  24 - 0x18
      13'h2F4: dout  = 8'b00111000; //  756 :  56 - 0x38
      13'h2F5: dout  = 8'b11111100; //  757 : 252 - 0xfc
      13'h2F6: dout  = 8'b11111100; //  758 : 252 - 0xfc
      13'h2F7: dout  = 8'b11111100; //  759 : 252 - 0xfc
      13'h2F8: dout  = 8'b01100110; //  760 : 102 - 0x66
      13'h2F9: dout  = 8'b01100000; //  761 :  96 - 0x60
      13'h2FA: dout  = 8'b01101000; //  762 : 104 - 0x68
      13'h2FB: dout  = 8'b11100000; //  763 : 224 - 0xe0
      13'h2FC: dout  = 8'b11000000; //  764 : 192 - 0xc0
      13'h2FD: dout  = 8'b00010000; //  765 :  16 - 0x10
      13'h2FE: dout  = 8'b00101000; //  766 :  40 - 0x28
      13'h2FF: dout  = 8'b01010000; //  767 :  80 - 0x50
      13'h300: dout  = 8'b01111111; //  768 : 127 - 0x7f -- Sprite 0x30
      13'h301: dout  = 8'b01111110; //  769 : 126 - 0x7e
      13'h302: dout  = 8'b11111100; //  770 : 252 - 0xfc
      13'h303: dout  = 8'b00111000; //  771 :  56 - 0x38
      13'h304: dout  = 8'b00111000; //  772 :  56 - 0x38
      13'h305: dout  = 8'b00000100; //  773 :   4 - 0x4
      13'h306: dout  = 8'b10000100; //  774 : 132 - 0x84
      13'h307: dout  = 8'b11111100; //  775 : 252 - 0xfc
      13'h308: dout  = 8'b11110110; //  776 : 246 - 0xf6
      13'h309: dout  = 8'b11110000; //  777 : 240 - 0xf0
      13'h30A: dout  = 8'b00111000; //  778 :  56 - 0x38
      13'h30B: dout  = 8'b11010000; //  779 : 208 - 0xd0
      13'h30C: dout  = 8'b11000000; //  780 : 192 - 0xc0
      13'h30D: dout  = 8'b11111000; //  781 : 248 - 0xf8
      13'h30E: dout  = 8'b01111000; //  782 : 120 - 0x78
      13'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout  = 8'b01111111; //  784 : 127 - 0x7f -- Sprite 0x31
      13'h311: dout  = 8'b01111110; //  785 : 126 - 0x7e
      13'h312: dout  = 8'b11111100; //  786 : 252 - 0xfc
      13'h313: dout  = 8'b00111000; //  787 :  56 - 0x38
      13'h314: dout  = 8'b00111000; //  788 :  56 - 0x38
      13'h315: dout  = 8'b00011100; //  789 :  28 - 0x1c
      13'h316: dout  = 8'b10000100; //  790 : 132 - 0x84
      13'h317: dout  = 8'b11000100; //  791 : 196 - 0xc4
      13'h318: dout  = 8'b11110110; //  792 : 246 - 0xf6
      13'h319: dout  = 8'b11110000; //  793 : 240 - 0xf0
      13'h31A: dout  = 8'b00111000; //  794 :  56 - 0x38
      13'h31B: dout  = 8'b11010000; //  795 : 208 - 0xd0
      13'h31C: dout  = 8'b11000000; //  796 : 192 - 0xc0
      13'h31D: dout  = 8'b11100000; //  797 : 224 - 0xe0
      13'h31E: dout  = 8'b01111000; //  798 : 120 - 0x78
      13'h31F: dout  = 8'b00111000; //  799 :  56 - 0x38
      13'h320: dout  = 8'b01111111; //  800 : 127 - 0x7f -- Sprite 0x32
      13'h321: dout  = 8'b01111110; //  801 : 126 - 0x7e
      13'h322: dout  = 8'b11111100; //  802 : 252 - 0xfc
      13'h323: dout  = 8'b00111000; //  803 :  56 - 0x38
      13'h324: dout  = 8'b00100100; //  804 :  36 - 0x24
      13'h325: dout  = 8'b00000100; //  805 :   4 - 0x4
      13'h326: dout  = 8'b10011100; //  806 : 156 - 0x9c
      13'h327: dout  = 8'b11111100; //  807 : 252 - 0xfc
      13'h328: dout  = 8'b11110110; //  808 : 246 - 0xf6
      13'h329: dout  = 8'b11110000; //  809 : 240 - 0xf0
      13'h32A: dout  = 8'b00111000; //  810 :  56 - 0x38
      13'h32B: dout  = 8'b11000000; //  811 : 192 - 0xc0
      13'h32C: dout  = 8'b11011000; //  812 : 216 - 0xd8
      13'h32D: dout  = 8'b11111000; //  813 : 248 - 0xf8
      13'h32E: dout  = 8'b01100000; //  814 :  96 - 0x60
      13'h32F: dout  = 8'b00010000; //  815 :  16 - 0x10
      13'h330: dout  = 8'b00100011; //  816 :  35 - 0x23 -- Sprite 0x33
      13'h331: dout  = 8'b00100011; //  817 :  35 - 0x23
      13'h332: dout  = 8'b00100001; //  818 :  33 - 0x21
      13'h333: dout  = 8'b00100000; //  819 :  32 - 0x20
      13'h334: dout  = 8'b00010011; //  820 :  19 - 0x13
      13'h335: dout  = 8'b00001101; //  821 :  13 - 0xd
      13'h336: dout  = 8'b00000001; //  822 :   1 - 0x1
      13'h337: dout  = 8'b00000001; //  823 :   1 - 0x1
      13'h338: dout  = 8'b00011100; //  824 :  28 - 0x1c
      13'h339: dout  = 8'b00011100; //  825 :  28 - 0x1c
      13'h33A: dout  = 8'b00011110; //  826 :  30 - 0x1e
      13'h33B: dout  = 8'b00011111; //  827 :  31 - 0x1f
      13'h33C: dout  = 8'b00001100; //  828 :  12 - 0xc
      13'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      13'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      13'h340: dout  = 8'b11111100; //  832 : 252 - 0xfc -- Sprite 0x34
      13'h341: dout  = 8'b11111100; //  833 : 252 - 0xfc
      13'h342: dout  = 8'b11111100; //  834 : 252 - 0xfc
      13'h343: dout  = 8'b11111100; //  835 : 252 - 0xfc
      13'h344: dout  = 8'b10100100; //  836 : 164 - 0xa4
      13'h345: dout  = 8'b00100100; //  837 :  36 - 0x24
      13'h346: dout  = 8'b00010010; //  838 :  18 - 0x12
      13'h347: dout  = 8'b11101110; //  839 : 238 - 0xee
      13'h348: dout  = 8'b10000000; //  840 : 128 - 0x80
      13'h349: dout  = 8'b01010000; //  841 :  80 - 0x50
      13'h34A: dout  = 8'b10101000; //  842 : 168 - 0xa8
      13'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      13'h34C: dout  = 8'b01011000; //  844 :  88 - 0x58
      13'h34D: dout  = 8'b11011000; //  845 : 216 - 0xd8
      13'h34E: dout  = 8'b11101100; //  846 : 236 - 0xec
      13'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      13'h350: dout  = 8'b00100011; //  848 :  35 - 0x23 -- Sprite 0x35
      13'h351: dout  = 8'b00100011; //  849 :  35 - 0x23
      13'h352: dout  = 8'b00100001; //  850 :  33 - 0x21
      13'h353: dout  = 8'b00100000; //  851 :  32 - 0x20
      13'h354: dout  = 8'b00010011; //  852 :  19 - 0x13
      13'h355: dout  = 8'b00001110; //  853 :  14 - 0xe
      13'h356: dout  = 8'b00000010; //  854 :   2 - 0x2
      13'h357: dout  = 8'b00000001; //  855 :   1 - 0x1
      13'h358: dout  = 8'b00011100; //  856 :  28 - 0x1c
      13'h359: dout  = 8'b00011100; //  857 :  28 - 0x1c
      13'h35A: dout  = 8'b00011110; //  858 :  30 - 0x1e
      13'h35B: dout  = 8'b00011111; //  859 :  31 - 0x1f
      13'h35C: dout  = 8'b00001100; //  860 :  12 - 0xc
      13'h35D: dout  = 8'b00000001; //  861 :   1 - 0x1
      13'h35E: dout  = 8'b00000001; //  862 :   1 - 0x1
      13'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout  = 8'b11111100; //  864 : 252 - 0xfc -- Sprite 0x36
      13'h361: dout  = 8'b11111100; //  865 : 252 - 0xfc
      13'h362: dout  = 8'b11111100; //  866 : 252 - 0xfc
      13'h363: dout  = 8'b11111100; //  867 : 252 - 0xfc
      13'h364: dout  = 8'b10100110; //  868 : 166 - 0xa6
      13'h365: dout  = 8'b00110001; //  869 :  49 - 0x31
      13'h366: dout  = 8'b01001001; //  870 :  73 - 0x49
      13'h367: dout  = 8'b11000110; //  871 : 198 - 0xc6
      13'h368: dout  = 8'b10101000; //  872 : 168 - 0xa8
      13'h369: dout  = 8'b01010000; //  873 :  80 - 0x50
      13'h36A: dout  = 8'b10101000; //  874 : 168 - 0xa8
      13'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      13'h36C: dout  = 8'b01011000; //  876 :  88 - 0x58
      13'h36D: dout  = 8'b11001110; //  877 : 206 - 0xce
      13'h36E: dout  = 8'b10000110; //  878 : 134 - 0x86
      13'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      13'h370: dout  = 8'b11111100; //  880 : 252 - 0xfc -- Sprite 0x37
      13'h371: dout  = 8'b11111100; //  881 : 252 - 0xfc
      13'h372: dout  = 8'b11111100; //  882 : 252 - 0xfc
      13'h373: dout  = 8'b11111100; //  883 : 252 - 0xfc
      13'h374: dout  = 8'b10100100; //  884 : 164 - 0xa4
      13'h375: dout  = 8'b00100100; //  885 :  36 - 0x24
      13'h376: dout  = 8'b00010010; //  886 :  18 - 0x12
      13'h377: dout  = 8'b11101110; //  887 : 238 - 0xee
      13'h378: dout  = 8'b10101000; //  888 : 168 - 0xa8
      13'h379: dout  = 8'b01010000; //  889 :  80 - 0x50
      13'h37A: dout  = 8'b10101000; //  890 : 168 - 0xa8
      13'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      13'h37C: dout  = 8'b01011000; //  892 :  88 - 0x58
      13'h37D: dout  = 8'b11011000; //  893 : 216 - 0xd8
      13'h37E: dout  = 8'b11101100; //  894 : 236 - 0xec
      13'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      13'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      13'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      13'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      13'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      13'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      13'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      13'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      13'h388: dout  = 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      13'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      13'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      13'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      13'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      13'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      13'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x39
      13'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      13'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      13'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      13'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      13'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      13'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout  = 8'b00000000; //  920 :   0 - 0x0
      13'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      13'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      13'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      13'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      13'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      13'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      13'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      13'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      13'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      13'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      13'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      13'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      13'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      13'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      13'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      13'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      13'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      13'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      13'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0
      13'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      13'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      13'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      13'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      13'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      13'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      13'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      13'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      13'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      13'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      13'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      13'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      13'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      13'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      13'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      13'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      13'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      13'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      13'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      13'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      13'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      13'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0
      13'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      13'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      13'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      13'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      13'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      13'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      13'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      13'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      13'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      13'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      13'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      13'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      13'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      13'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      13'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      13'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      13'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      13'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      13'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      13'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      13'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      13'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      13'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      13'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      13'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      13'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      13'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      13'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      13'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0
      13'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      13'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      13'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      13'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      13'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      13'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      13'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      13'h401: dout  = 8'b00111110; // 1025 :  62 - 0x3e
      13'h402: dout  = 8'b01111111; // 1026 : 127 - 0x7f
      13'h403: dout  = 8'b01111111; // 1027 : 127 - 0x7f
      13'h404: dout  = 8'b01111111; // 1028 : 127 - 0x7f
      13'h405: dout  = 8'b01111111; // 1029 : 127 - 0x7f
      13'h406: dout  = 8'b01111111; // 1030 : 127 - 0x7f
      13'h407: dout  = 8'b00111110; // 1031 :  62 - 0x3e
      13'h408: dout  = 8'b00111100; // 1032 :  60 - 0x3c
      13'h409: dout  = 8'b01111100; // 1033 : 124 - 0x7c
      13'h40A: dout  = 8'b11100110; // 1034 : 230 - 0xe6
      13'h40B: dout  = 8'b11101110; // 1035 : 238 - 0xee
      13'h40C: dout  = 8'b11110110; // 1036 : 246 - 0xf6
      13'h40D: dout  = 8'b11100110; // 1037 : 230 - 0xe6
      13'h40E: dout  = 8'b00111100; // 1038 :  60 - 0x3c
      13'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      13'h411: dout  = 8'b00111100; // 1041 :  60 - 0x3c
      13'h412: dout  = 8'b00011100; // 1042 :  28 - 0x1c
      13'h413: dout  = 8'b00011100; // 1043 :  28 - 0x1c
      13'h414: dout  = 8'b00011100; // 1044 :  28 - 0x1c
      13'h415: dout  = 8'b00011100; // 1045 :  28 - 0x1c
      13'h416: dout  = 8'b00011100; // 1046 :  28 - 0x1c
      13'h417: dout  = 8'b00011100; // 1047 :  28 - 0x1c
      13'h418: dout  = 8'b00111000; // 1048 :  56 - 0x38
      13'h419: dout  = 8'b01111000; // 1049 : 120 - 0x78
      13'h41A: dout  = 8'b00111000; // 1050 :  56 - 0x38
      13'h41B: dout  = 8'b00111000; // 1051 :  56 - 0x38
      13'h41C: dout  = 8'b00111000; // 1052 :  56 - 0x38
      13'h41D: dout  = 8'b00111000; // 1053 :  56 - 0x38
      13'h41E: dout  = 8'b00111000; // 1054 :  56 - 0x38
      13'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      13'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x42
      13'h421: dout  = 8'b01111100; // 1057 : 124 - 0x7c
      13'h422: dout  = 8'b01111111; // 1058 : 127 - 0x7f
      13'h423: dout  = 8'b01100111; // 1059 : 103 - 0x67
      13'h424: dout  = 8'b00111111; // 1060 :  63 - 0x3f
      13'h425: dout  = 8'b01111110; // 1061 : 126 - 0x7e
      13'h426: dout  = 8'b01111111; // 1062 : 127 - 0x7f
      13'h427: dout  = 8'b01111111; // 1063 : 127 - 0x7f
      13'h428: dout  = 8'b01111100; // 1064 : 124 - 0x7c
      13'h429: dout  = 8'b11111110; // 1065 : 254 - 0xfe
      13'h42A: dout  = 8'b11100110; // 1066 : 230 - 0xe6
      13'h42B: dout  = 8'b00011110; // 1067 :  30 - 0x1e
      13'h42C: dout  = 8'b01111100; // 1068 : 124 - 0x7c
      13'h42D: dout  = 8'b11100000; // 1069 : 224 - 0xe0
      13'h42E: dout  = 8'b11111110; // 1070 : 254 - 0xfe
      13'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      13'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      13'h431: dout  = 8'b01111110; // 1073 : 126 - 0x7e
      13'h432: dout  = 8'b01111111; // 1074 : 127 - 0x7f
      13'h433: dout  = 8'b01111111; // 1075 : 127 - 0x7f
      13'h434: dout  = 8'b00011111; // 1076 :  31 - 0x1f
      13'h435: dout  = 8'b01110111; // 1077 : 119 - 0x77
      13'h436: dout  = 8'b01111111; // 1078 : 127 - 0x7f
      13'h437: dout  = 8'b01111110; // 1079 : 126 - 0x7e
      13'h438: dout  = 8'b01111100; // 1080 : 124 - 0x7c
      13'h439: dout  = 8'b11111100; // 1081 : 252 - 0xfc
      13'h43A: dout  = 8'b11100110; // 1082 : 230 - 0xe6
      13'h43B: dout  = 8'b00011100; // 1083 :  28 - 0x1c
      13'h43C: dout  = 8'b01100110; // 1084 : 102 - 0x66
      13'h43D: dout  = 8'b11101110; // 1085 : 238 - 0xee
      13'h43E: dout  = 8'b11111100; // 1086 : 252 - 0xfc
      13'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      13'h441: dout  = 8'b00001110; // 1089 :  14 - 0xe
      13'h442: dout  = 8'b00011110; // 1090 :  30 - 0x1e
      13'h443: dout  = 8'b00111110; // 1091 :  62 - 0x3e
      13'h444: dout  = 8'b01111110; // 1092 : 126 - 0x7e
      13'h445: dout  = 8'b01111111; // 1093 : 127 - 0x7f
      13'h446: dout  = 8'b01111110; // 1094 : 126 - 0x7e
      13'h447: dout  = 8'b00001100; // 1095 :  12 - 0xc
      13'h448: dout  = 8'b00001100; // 1096 :  12 - 0xc
      13'h449: dout  = 8'b00011100; // 1097 :  28 - 0x1c
      13'h44A: dout  = 8'b00111100; // 1098 :  60 - 0x3c
      13'h44B: dout  = 8'b01111100; // 1099 : 124 - 0x7c
      13'h44C: dout  = 8'b11101100; // 1100 : 236 - 0xec
      13'h44D: dout  = 8'b11111110; // 1101 : 254 - 0xfe
      13'h44E: dout  = 8'b00001100; // 1102 :  12 - 0xc
      13'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      13'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x45
      13'h451: dout  = 8'b01111111; // 1105 : 127 - 0x7f
      13'h452: dout  = 8'b01111111; // 1106 : 127 - 0x7f
      13'h453: dout  = 8'b01111111; // 1107 : 127 - 0x7f
      13'h454: dout  = 8'b01111111; // 1108 : 127 - 0x7f
      13'h455: dout  = 8'b01110111; // 1109 : 119 - 0x77
      13'h456: dout  = 8'b01111111; // 1110 : 127 - 0x7f
      13'h457: dout  = 8'b01111110; // 1111 : 126 - 0x7e
      13'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe
      13'h459: dout  = 8'b11111110; // 1113 : 254 - 0xfe
      13'h45A: dout  = 8'b11100000; // 1114 : 224 - 0xe0
      13'h45B: dout  = 8'b11111110; // 1115 : 254 - 0xfe
      13'h45C: dout  = 8'b00000110; // 1116 :   6 - 0x6
      13'h45D: dout  = 8'b11101110; // 1117 : 238 - 0xee
      13'h45E: dout  = 8'b11111100; // 1118 : 252 - 0xfc
      13'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      13'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x46
      13'h461: dout  = 8'b00111110; // 1121 :  62 - 0x3e
      13'h462: dout  = 8'b01111110; // 1122 : 126 - 0x7e
      13'h463: dout  = 8'b01111111; // 1123 : 127 - 0x7f
      13'h464: dout  = 8'b01111111; // 1124 : 127 - 0x7f
      13'h465: dout  = 8'b01110111; // 1125 : 119 - 0x77
      13'h466: dout  = 8'b01111111; // 1126 : 127 - 0x7f
      13'h467: dout  = 8'b00111110; // 1127 :  62 - 0x3e
      13'h468: dout  = 8'b00111100; // 1128 :  60 - 0x3c
      13'h469: dout  = 8'b01111100; // 1129 : 124 - 0x7c
      13'h46A: dout  = 8'b11100000; // 1130 : 224 - 0xe0
      13'h46B: dout  = 8'b11111110; // 1131 : 254 - 0xfe
      13'h46C: dout  = 8'b11100110; // 1132 : 230 - 0xe6
      13'h46D: dout  = 8'b11101110; // 1133 : 238 - 0xee
      13'h46E: dout  = 8'b00111100; // 1134 :  60 - 0x3c
      13'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x47
      13'h471: dout  = 8'b01111110; // 1137 : 126 - 0x7e
      13'h472: dout  = 8'b01111110; // 1138 : 126 - 0x7e
      13'h473: dout  = 8'b00011110; // 1139 :  30 - 0x1e
      13'h474: dout  = 8'b00011100; // 1140 :  28 - 0x1c
      13'h475: dout  = 8'b00111100; // 1141 :  60 - 0x3c
      13'h476: dout  = 8'b00111000; // 1142 :  56 - 0x38
      13'h477: dout  = 8'b00111000; // 1143 :  56 - 0x38
      13'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe
      13'h479: dout  = 8'b11111100; // 1145 : 252 - 0xfc
      13'h47A: dout  = 8'b00001100; // 1146 :  12 - 0xc
      13'h47B: dout  = 8'b00111000; // 1147 :  56 - 0x38
      13'h47C: dout  = 8'b00111000; // 1148 :  56 - 0x38
      13'h47D: dout  = 8'b01110000; // 1149 : 112 - 0x70
      13'h47E: dout  = 8'b01110000; // 1150 : 112 - 0x70
      13'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      13'h481: dout  = 8'b00111110; // 1153 :  62 - 0x3e
      13'h482: dout  = 8'b01111111; // 1154 : 127 - 0x7f
      13'h483: dout  = 8'b01111111; // 1155 : 127 - 0x7f
      13'h484: dout  = 8'b01111111; // 1156 : 127 - 0x7f
      13'h485: dout  = 8'b01111111; // 1157 : 127 - 0x7f
      13'h486: dout  = 8'b01111111; // 1158 : 127 - 0x7f
      13'h487: dout  = 8'b00111110; // 1159 :  62 - 0x3e
      13'h488: dout  = 8'b00111110; // 1160 :  62 - 0x3e
      13'h489: dout  = 8'b01111100; // 1161 : 124 - 0x7c
      13'h48A: dout  = 8'b11100110; // 1162 : 230 - 0xe6
      13'h48B: dout  = 8'b10111100; // 1163 : 188 - 0xbc
      13'h48C: dout  = 8'b11100110; // 1164 : 230 - 0xe6
      13'h48D: dout  = 8'b11101110; // 1165 : 238 - 0xee
      13'h48E: dout  = 8'b00111100; // 1166 :  60 - 0x3c
      13'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      13'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x49
      13'h491: dout  = 8'b00111110; // 1169 :  62 - 0x3e
      13'h492: dout  = 8'b01111111; // 1170 : 127 - 0x7f
      13'h493: dout  = 8'b01110111; // 1171 : 119 - 0x77
      13'h494: dout  = 8'b01111111; // 1172 : 127 - 0x7f
      13'h495: dout  = 8'b01111111; // 1173 : 127 - 0x7f
      13'h496: dout  = 8'b00111111; // 1174 :  63 - 0x3f
      13'h497: dout  = 8'b00111110; // 1175 :  62 - 0x3e
      13'h498: dout  = 8'b00111100; // 1176 :  60 - 0x3c
      13'h499: dout  = 8'b01111100; // 1177 : 124 - 0x7c
      13'h49A: dout  = 8'b11100110; // 1178 : 230 - 0xe6
      13'h49B: dout  = 8'b11101110; // 1179 : 238 - 0xee
      13'h49C: dout  = 8'b11111110; // 1180 : 254 - 0xfe
      13'h49D: dout  = 8'b10000110; // 1181 : 134 - 0x86
      13'h49E: dout  = 8'b01111100; // 1182 : 124 - 0x7c
      13'h49F: dout  = 8'b01000000; // 1183 :  64 - 0x40
      13'h4A0: dout  = 8'b11111111; // 1184 : 255 - 0xff -- Sprite 0x4a
      13'h4A1: dout  = 8'b10011001; // 1185 : 153 - 0x99
      13'h4A2: dout  = 8'b10011001; // 1186 : 153 - 0x99
      13'h4A3: dout  = 8'b10011001; // 1187 : 153 - 0x99
      13'h4A4: dout  = 8'b10011001; // 1188 : 153 - 0x99
      13'h4A5: dout  = 8'b10011001; // 1189 : 153 - 0x99
      13'h4A6: dout  = 8'b10011001; // 1190 : 153 - 0x99
      13'h4A7: dout  = 8'b11111111; // 1191 : 255 - 0xff
      13'h4A8: dout  = 8'b11101110; // 1192 : 238 - 0xee
      13'h4A9: dout  = 8'b11101110; // 1193 : 238 - 0xee
      13'h4AA: dout  = 8'b11101110; // 1194 : 238 - 0xee
      13'h4AB: dout  = 8'b11101110; // 1195 : 238 - 0xee
      13'h4AC: dout  = 8'b11101110; // 1196 : 238 - 0xee
      13'h4AD: dout  = 8'b11101110; // 1197 : 238 - 0xee
      13'h4AE: dout  = 8'b11101110; // 1198 : 238 - 0xee
      13'h4AF: dout  = 8'b10001000; // 1199 : 136 - 0x88
      13'h4B0: dout  = 8'b11110000; // 1200 : 240 - 0xf0 -- Sprite 0x4b
      13'h4B1: dout  = 8'b10010000; // 1201 : 144 - 0x90
      13'h4B2: dout  = 8'b10010000; // 1202 : 144 - 0x90
      13'h4B3: dout  = 8'b10010000; // 1203 : 144 - 0x90
      13'h4B4: dout  = 8'b10010000; // 1204 : 144 - 0x90
      13'h4B5: dout  = 8'b10010000; // 1205 : 144 - 0x90
      13'h4B6: dout  = 8'b10010000; // 1206 : 144 - 0x90
      13'h4B7: dout  = 8'b11110000; // 1207 : 240 - 0xf0
      13'h4B8: dout  = 8'b11100000; // 1208 : 224 - 0xe0
      13'h4B9: dout  = 8'b11100000; // 1209 : 224 - 0xe0
      13'h4BA: dout  = 8'b11100000; // 1210 : 224 - 0xe0
      13'h4BB: dout  = 8'b11100000; // 1211 : 224 - 0xe0
      13'h4BC: dout  = 8'b11100000; // 1212 : 224 - 0xe0
      13'h4BD: dout  = 8'b11100000; // 1213 : 224 - 0xe0
      13'h4BE: dout  = 8'b11100000; // 1214 : 224 - 0xe0
      13'h4BF: dout  = 8'b10000000; // 1215 : 128 - 0x80
      13'h4C0: dout  = 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x4c
      13'h4C1: dout  = 8'b11111111; // 1217 : 255 - 0xff
      13'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      13'h4C3: dout  = 8'b11111111; // 1219 : 255 - 0xff
      13'h4C4: dout  = 8'b11111111; // 1220 : 255 - 0xff
      13'h4C5: dout  = 8'b11111111; // 1221 : 255 - 0xff
      13'h4C6: dout  = 8'b11111111; // 1222 : 255 - 0xff
      13'h4C7: dout  = 8'b11111111; // 1223 : 255 - 0xff
      13'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout  = 8'b01111111; // 1225 : 127 - 0x7f
      13'h4CA: dout  = 8'b01111111; // 1226 : 127 - 0x7f
      13'h4CB: dout  = 8'b01111111; // 1227 : 127 - 0x7f
      13'h4CC: dout  = 8'b01111111; // 1228 : 127 - 0x7f
      13'h4CD: dout  = 8'b01111111; // 1229 : 127 - 0x7f
      13'h4CE: dout  = 8'b01111111; // 1230 : 127 - 0x7f
      13'h4CF: dout  = 8'b01111111; // 1231 : 127 - 0x7f
      13'h4D0: dout  = 8'b11111111; // 1232 : 255 - 0xff -- Sprite 0x4d
      13'h4D1: dout  = 8'b11111111; // 1233 : 255 - 0xff
      13'h4D2: dout  = 8'b11111111; // 1234 : 255 - 0xff
      13'h4D3: dout  = 8'b11111111; // 1235 : 255 - 0xff
      13'h4D4: dout  = 8'b11111111; // 1236 : 255 - 0xff
      13'h4D5: dout  = 8'b11111111; // 1237 : 255 - 0xff
      13'h4D6: dout  = 8'b11111111; // 1238 : 255 - 0xff
      13'h4D7: dout  = 8'b11111111; // 1239 : 255 - 0xff
      13'h4D8: dout  = 8'b01111111; // 1240 : 127 - 0x7f
      13'h4D9: dout  = 8'b01111111; // 1241 : 127 - 0x7f
      13'h4DA: dout  = 8'b01111111; // 1242 : 127 - 0x7f
      13'h4DB: dout  = 8'b01111111; // 1243 : 127 - 0x7f
      13'h4DC: dout  = 8'b01111111; // 1244 : 127 - 0x7f
      13'h4DD: dout  = 8'b01111111; // 1245 : 127 - 0x7f
      13'h4DE: dout  = 8'b01111111; // 1246 : 127 - 0x7f
      13'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout  = 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x4e
      13'h4E1: dout  = 8'b11111111; // 1249 : 255 - 0xff
      13'h4E2: dout  = 8'b11111111; // 1250 : 255 - 0xff
      13'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      13'h4E4: dout  = 8'b11111111; // 1252 : 255 - 0xff
      13'h4E5: dout  = 8'b11111111; // 1253 : 255 - 0xff
      13'h4E6: dout  = 8'b11111111; // 1254 : 255 - 0xff
      13'h4E7: dout  = 8'b11111111; // 1255 : 255 - 0xff
      13'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout  = 8'b11111110; // 1257 : 254 - 0xfe
      13'h4EA: dout  = 8'b11111110; // 1258 : 254 - 0xfe
      13'h4EB: dout  = 8'b11111110; // 1259 : 254 - 0xfe
      13'h4EC: dout  = 8'b11111110; // 1260 : 254 - 0xfe
      13'h4ED: dout  = 8'b11111110; // 1261 : 254 - 0xfe
      13'h4EE: dout  = 8'b11111110; // 1262 : 254 - 0xfe
      13'h4EF: dout  = 8'b11111110; // 1263 : 254 - 0xfe
      13'h4F0: dout  = 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x4f
      13'h4F1: dout  = 8'b11111111; // 1265 : 255 - 0xff
      13'h4F2: dout  = 8'b11111111; // 1266 : 255 - 0xff
      13'h4F3: dout  = 8'b11111111; // 1267 : 255 - 0xff
      13'h4F4: dout  = 8'b11111111; // 1268 : 255 - 0xff
      13'h4F5: dout  = 8'b11111111; // 1269 : 255 - 0xff
      13'h4F6: dout  = 8'b11111111; // 1270 : 255 - 0xff
      13'h4F7: dout  = 8'b11111111; // 1271 : 255 - 0xff
      13'h4F8: dout  = 8'b11111110; // 1272 : 254 - 0xfe
      13'h4F9: dout  = 8'b11111110; // 1273 : 254 - 0xfe
      13'h4FA: dout  = 8'b11111110; // 1274 : 254 - 0xfe
      13'h4FB: dout  = 8'b11111110; // 1275 : 254 - 0xfe
      13'h4FC: dout  = 8'b11111110; // 1276 : 254 - 0xfe
      13'h4FD: dout  = 8'b11111110; // 1277 : 254 - 0xfe
      13'h4FE: dout  = 8'b11111110; // 1278 : 254 - 0xfe
      13'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      13'h500: dout  = 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0x50
      13'h501: dout  = 8'b00101000; // 1281 :  40 - 0x28
      13'h502: dout  = 8'b11101110; // 1282 : 238 - 0xee
      13'h503: dout  = 8'b10000010; // 1283 : 130 - 0x82
      13'h504: dout  = 8'b01000100; // 1284 :  68 - 0x44
      13'h505: dout  = 8'b01000100; // 1285 :  68 - 0x44
      13'h506: dout  = 8'b10010010; // 1286 : 146 - 0x92
      13'h507: dout  = 8'b11101110; // 1287 : 238 - 0xee
      13'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      13'h50A: dout  = 8'b00000000; // 1290 :   0 - 0x0
      13'h50B: dout  = 8'b00000000; // 1291 :   0 - 0x0
      13'h50C: dout  = 8'b00000000; // 1292 :   0 - 0x0
      13'h50D: dout  = 8'b00000000; // 1293 :   0 - 0x0
      13'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      13'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      13'h510: dout  = 8'b00010000; // 1296 :  16 - 0x10 -- Sprite 0x51
      13'h511: dout  = 8'b00101000; // 1297 :  40 - 0x28
      13'h512: dout  = 8'b11101110; // 1298 : 238 - 0xee
      13'h513: dout  = 8'b10000010; // 1299 : 130 - 0x82
      13'h514: dout  = 8'b01000100; // 1300 :  68 - 0x44
      13'h515: dout  = 8'b01000100; // 1301 :  68 - 0x44
      13'h516: dout  = 8'b10010010; // 1302 : 146 - 0x92
      13'h517: dout  = 8'b11101110; // 1303 : 238 - 0xee
      13'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout  = 8'b00010000; // 1305 :  16 - 0x10
      13'h51A: dout  = 8'b00010000; // 1306 :  16 - 0x10
      13'h51B: dout  = 8'b01111100; // 1307 : 124 - 0x7c
      13'h51C: dout  = 8'b00111000; // 1308 :  56 - 0x38
      13'h51D: dout  = 8'b00111000; // 1309 :  56 - 0x38
      13'h51E: dout  = 8'b01101100; // 1310 : 108 - 0x6c
      13'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      13'h520: dout  = 8'b00010000; // 1312 :  16 - 0x10 -- Sprite 0x52
      13'h521: dout  = 8'b00111000; // 1313 :  56 - 0x38
      13'h522: dout  = 8'b11111110; // 1314 : 254 - 0xfe
      13'h523: dout  = 8'b11111110; // 1315 : 254 - 0xfe
      13'h524: dout  = 8'b01111100; // 1316 : 124 - 0x7c
      13'h525: dout  = 8'b01111100; // 1317 : 124 - 0x7c
      13'h526: dout  = 8'b11111110; // 1318 : 254 - 0xfe
      13'h527: dout  = 8'b11101110; // 1319 : 238 - 0xee
      13'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout  = 8'b00010000; // 1321 :  16 - 0x10
      13'h52A: dout  = 8'b00010000; // 1322 :  16 - 0x10
      13'h52B: dout  = 8'b01111100; // 1323 : 124 - 0x7c
      13'h52C: dout  = 8'b00111000; // 1324 :  56 - 0x38
      13'h52D: dout  = 8'b00111000; // 1325 :  56 - 0x38
      13'h52E: dout  = 8'b01101100; // 1326 : 108 - 0x6c
      13'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      13'h530: dout  = 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      13'h531: dout  = 8'b11111111; // 1329 : 255 - 0xff
      13'h532: dout  = 8'b11111111; // 1330 : 255 - 0xff
      13'h533: dout  = 8'b11111111; // 1331 : 255 - 0xff
      13'h534: dout  = 8'b11111111; // 1332 : 255 - 0xff
      13'h535: dout  = 8'b11111111; // 1333 : 255 - 0xff
      13'h536: dout  = 8'b11111111; // 1334 : 255 - 0xff
      13'h537: dout  = 8'b11111111; // 1335 : 255 - 0xff
      13'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout  = 8'b00000000; // 1338 :   0 - 0x0
      13'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      13'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      13'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      13'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0x54
      13'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      13'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      13'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      13'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      13'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      13'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      13'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      13'h548: dout  = 8'b11111111; // 1352 : 255 - 0xff
      13'h549: dout  = 8'b11111111; // 1353 : 255 - 0xff
      13'h54A: dout  = 8'b11111111; // 1354 : 255 - 0xff
      13'h54B: dout  = 8'b11111111; // 1355 : 255 - 0xff
      13'h54C: dout  = 8'b11111111; // 1356 : 255 - 0xff
      13'h54D: dout  = 8'b11111111; // 1357 : 255 - 0xff
      13'h54E: dout  = 8'b11111111; // 1358 : 255 - 0xff
      13'h54F: dout  = 8'b11111111; // 1359 : 255 - 0xff
      13'h550: dout  = 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      13'h551: dout  = 8'b11111111; // 1361 : 255 - 0xff
      13'h552: dout  = 8'b11111111; // 1362 : 255 - 0xff
      13'h553: dout  = 8'b11111111; // 1363 : 255 - 0xff
      13'h554: dout  = 8'b11111111; // 1364 : 255 - 0xff
      13'h555: dout  = 8'b11111111; // 1365 : 255 - 0xff
      13'h556: dout  = 8'b11111111; // 1366 : 255 - 0xff
      13'h557: dout  = 8'b11111111; // 1367 : 255 - 0xff
      13'h558: dout  = 8'b11111111; // 1368 : 255 - 0xff
      13'h559: dout  = 8'b11111111; // 1369 : 255 - 0xff
      13'h55A: dout  = 8'b11111111; // 1370 : 255 - 0xff
      13'h55B: dout  = 8'b11111111; // 1371 : 255 - 0xff
      13'h55C: dout  = 8'b11111111; // 1372 : 255 - 0xff
      13'h55D: dout  = 8'b11111111; // 1373 : 255 - 0xff
      13'h55E: dout  = 8'b11111111; // 1374 : 255 - 0xff
      13'h55F: dout  = 8'b11111111; // 1375 : 255 - 0xff
      13'h560: dout  = 8'b00101010; // 1376 :  42 - 0x2a -- Sprite 0x56
      13'h561: dout  = 8'b01000101; // 1377 :  69 - 0x45
      13'h562: dout  = 8'b00001000; // 1378 :   8 - 0x8
      13'h563: dout  = 8'b00010101; // 1379 :  21 - 0x15
      13'h564: dout  = 8'b00100000; // 1380 :  32 - 0x20
      13'h565: dout  = 8'b01000101; // 1381 :  69 - 0x45
      13'h566: dout  = 8'b10101000; // 1382 : 168 - 0xa8
      13'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      13'h568: dout  = 8'b00000010; // 1384 :   2 - 0x2
      13'h569: dout  = 8'b00000101; // 1385 :   5 - 0x5
      13'h56A: dout  = 8'b10101010; // 1386 : 170 - 0xaa
      13'h56B: dout  = 8'b01010001; // 1387 :  81 - 0x51
      13'h56C: dout  = 8'b10101010; // 1388 : 170 - 0xaa
      13'h56D: dout  = 8'b01010001; // 1389 :  81 - 0x51
      13'h56E: dout  = 8'b10100010; // 1390 : 162 - 0xa2
      13'h56F: dout  = 8'b00000100; // 1391 :   4 - 0x4
      13'h570: dout  = 8'b00001000; // 1392 :   8 - 0x8 -- Sprite 0x57
      13'h571: dout  = 8'b01010101; // 1393 :  85 - 0x55
      13'h572: dout  = 8'b10100000; // 1394 : 160 - 0xa0
      13'h573: dout  = 8'b00010000; // 1395 :  16 - 0x10
      13'h574: dout  = 8'b10000000; // 1396 : 128 - 0x80
      13'h575: dout  = 8'b00010100; // 1397 :  20 - 0x14
      13'h576: dout  = 8'b00100010; // 1398 :  34 - 0x22
      13'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout  = 8'b00001000; // 1400 :   8 - 0x8
      13'h579: dout  = 8'b01010101; // 1401 :  85 - 0x55
      13'h57A: dout  = 8'b00101010; // 1402 :  42 - 0x2a
      13'h57B: dout  = 8'b01010101; // 1403 :  85 - 0x55
      13'h57C: dout  = 8'b00101010; // 1404 :  42 - 0x2a
      13'h57D: dout  = 8'b01000101; // 1405 :  69 - 0x45
      13'h57E: dout  = 8'b00001010; // 1406 :  10 - 0xa
      13'h57F: dout  = 8'b00010000; // 1407 :  16 - 0x10
      13'h580: dout  = 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      13'h581: dout  = 8'b11010101; // 1409 : 213 - 0xd5
      13'h582: dout  = 8'b10100000; // 1410 : 160 - 0xa0
      13'h583: dout  = 8'b11010000; // 1411 : 208 - 0xd0
      13'h584: dout  = 8'b10001111; // 1412 : 143 - 0x8f
      13'h585: dout  = 8'b11001000; // 1413 : 200 - 0xc8
      13'h586: dout  = 8'b10001000; // 1414 : 136 - 0x88
      13'h587: dout  = 8'b11001000; // 1415 : 200 - 0xc8
      13'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0
      13'h589: dout  = 8'b00111111; // 1417 :  63 - 0x3f
      13'h58A: dout  = 8'b01011111; // 1418 :  95 - 0x5f
      13'h58B: dout  = 8'b01101111; // 1419 : 111 - 0x6f
      13'h58C: dout  = 8'b01110000; // 1420 : 112 - 0x70
      13'h58D: dout  = 8'b01110111; // 1421 : 119 - 0x77
      13'h58E: dout  = 8'b01110111; // 1422 : 119 - 0x77
      13'h58F: dout  = 8'b01110111; // 1423 : 119 - 0x77
      13'h590: dout  = 8'b10001000; // 1424 : 136 - 0x88 -- Sprite 0x59
      13'h591: dout  = 8'b11001000; // 1425 : 200 - 0xc8
      13'h592: dout  = 8'b10001000; // 1426 : 136 - 0x88
      13'h593: dout  = 8'b11001111; // 1427 : 207 - 0xcf
      13'h594: dout  = 8'b10010000; // 1428 : 144 - 0x90
      13'h595: dout  = 8'b11100000; // 1429 : 224 - 0xe0
      13'h596: dout  = 8'b11101010; // 1430 : 234 - 0xea
      13'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      13'h598: dout  = 8'b01110111; // 1432 : 119 - 0x77
      13'h599: dout  = 8'b01110111; // 1433 : 119 - 0x77
      13'h59A: dout  = 8'b01110111; // 1434 : 119 - 0x77
      13'h59B: dout  = 8'b01110000; // 1435 : 112 - 0x70
      13'h59C: dout  = 8'b01101111; // 1436 : 111 - 0x6f
      13'h59D: dout  = 8'b01011111; // 1437 :  95 - 0x5f
      13'h59E: dout  = 8'b00010101; // 1438 :  21 - 0x15
      13'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      13'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      13'h5A1: dout  = 8'b01011011; // 1441 :  91 - 0x5b
      13'h5A2: dout  = 8'b00000111; // 1442 :   7 - 0x7
      13'h5A3: dout  = 8'b00001001; // 1443 :   9 - 0x9
      13'h5A4: dout  = 8'b11110011; // 1444 : 243 - 0xf3
      13'h5A5: dout  = 8'b00010001; // 1445 :  17 - 0x11
      13'h5A6: dout  = 8'b00010011; // 1446 :  19 - 0x13
      13'h5A7: dout  = 8'b00010001; // 1447 :  17 - 0x11
      13'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0
      13'h5A9: dout  = 8'b11111100; // 1449 : 252 - 0xfc
      13'h5AA: dout  = 8'b11111000; // 1450 : 248 - 0xf8
      13'h5AB: dout  = 8'b11110110; // 1451 : 246 - 0xf6
      13'h5AC: dout  = 8'b00001100; // 1452 :  12 - 0xc
      13'h5AD: dout  = 8'b11101110; // 1453 : 238 - 0xee
      13'h5AE: dout  = 8'b11101100; // 1454 : 236 - 0xec
      13'h5AF: dout  = 8'b11101110; // 1455 : 238 - 0xee
      13'h5B0: dout  = 8'b00010011; // 1456 :  19 - 0x13 -- Sprite 0x5b
      13'h5B1: dout  = 8'b00010001; // 1457 :  17 - 0x11
      13'h5B2: dout  = 8'b00010011; // 1458 :  19 - 0x13
      13'h5B3: dout  = 8'b11110001; // 1459 : 241 - 0xf1
      13'h5B4: dout  = 8'b00001011; // 1460 :  11 - 0xb
      13'h5B5: dout  = 8'b00000101; // 1461 :   5 - 0x5
      13'h5B6: dout  = 8'b10101011; // 1462 : 171 - 0xab
      13'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      13'h5B8: dout  = 8'b11101100; // 1464 : 236 - 0xec
      13'h5B9: dout  = 8'b11101110; // 1465 : 238 - 0xee
      13'h5BA: dout  = 8'b11101100; // 1466 : 236 - 0xec
      13'h5BB: dout  = 8'b00001110; // 1467 :  14 - 0xe
      13'h5BC: dout  = 8'b11110100; // 1468 : 244 - 0xf4
      13'h5BD: dout  = 8'b11111010; // 1469 : 250 - 0xfa
      13'h5BE: dout  = 8'b01010100; // 1470 :  84 - 0x54
      13'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      13'h5C0: dout  = 8'b00011100; // 1472 :  28 - 0x1c -- Sprite 0x5c
      13'h5C1: dout  = 8'b00100010; // 1473 :  34 - 0x22
      13'h5C2: dout  = 8'b01000001; // 1474 :  65 - 0x41
      13'h5C3: dout  = 8'b01000001; // 1475 :  65 - 0x41
      13'h5C4: dout  = 8'b01000001; // 1476 :  65 - 0x41
      13'h5C5: dout  = 8'b00100010; // 1477 :  34 - 0x22
      13'h5C6: dout  = 8'b00100010; // 1478 :  34 - 0x22
      13'h5C7: dout  = 8'b00011100; // 1479 :  28 - 0x1c
      13'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout  = 8'b00011100; // 1481 :  28 - 0x1c
      13'h5CA: dout  = 8'b00111110; // 1482 :  62 - 0x3e
      13'h5CB: dout  = 8'b00111110; // 1483 :  62 - 0x3e
      13'h5CC: dout  = 8'b00111110; // 1484 :  62 - 0x3e
      13'h5CD: dout  = 8'b00011100; // 1485 :  28 - 0x1c
      13'h5CE: dout  = 8'b00011100; // 1486 :  28 - 0x1c
      13'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      13'h5D0: dout  = 8'b00001000; // 1488 :   8 - 0x8 -- Sprite 0x5d
      13'h5D1: dout  = 8'b00010000; // 1489 :  16 - 0x10
      13'h5D2: dout  = 8'b00010000; // 1490 :  16 - 0x10
      13'h5D3: dout  = 8'b00001000; // 1491 :   8 - 0x8
      13'h5D4: dout  = 8'b00000100; // 1492 :   4 - 0x4
      13'h5D5: dout  = 8'b00000100; // 1493 :   4 - 0x4
      13'h5D6: dout  = 8'b00001000; // 1494 :   8 - 0x8
      13'h5D7: dout  = 8'b00010000; // 1495 :  16 - 0x10
      13'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      13'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      13'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      13'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      13'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      13'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      13'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      13'h5E0: dout  = 8'b00110110; // 1504 :  54 - 0x36 -- Sprite 0x5e
      13'h5E1: dout  = 8'b01101011; // 1505 : 107 - 0x6b
      13'h5E2: dout  = 8'b01001001; // 1506 :  73 - 0x49
      13'h5E3: dout  = 8'b01000001; // 1507 :  65 - 0x41
      13'h5E4: dout  = 8'b01000001; // 1508 :  65 - 0x41
      13'h5E5: dout  = 8'b00100010; // 1509 :  34 - 0x22
      13'h5E6: dout  = 8'b00010100; // 1510 :  20 - 0x14
      13'h5E7: dout  = 8'b00001000; // 1511 :   8 - 0x8
      13'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout  = 8'b00010100; // 1513 :  20 - 0x14
      13'h5EA: dout  = 8'b00110110; // 1514 :  54 - 0x36
      13'h5EB: dout  = 8'b00111110; // 1515 :  62 - 0x3e
      13'h5EC: dout  = 8'b00111110; // 1516 :  62 - 0x3e
      13'h5ED: dout  = 8'b00011100; // 1517 :  28 - 0x1c
      13'h5EE: dout  = 8'b00001000; // 1518 :   8 - 0x8
      13'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      13'h5F0: dout  = 8'b00111110; // 1520 :  62 - 0x3e -- Sprite 0x5f
      13'h5F1: dout  = 8'b01101011; // 1521 : 107 - 0x6b
      13'h5F2: dout  = 8'b00100010; // 1522 :  34 - 0x22
      13'h5F3: dout  = 8'b01100011; // 1523 :  99 - 0x63
      13'h5F4: dout  = 8'b00100010; // 1524 :  34 - 0x22
      13'h5F5: dout  = 8'b01100011; // 1525 :  99 - 0x63
      13'h5F6: dout  = 8'b00100010; // 1526 :  34 - 0x22
      13'h5F7: dout  = 8'b01111111; // 1527 : 127 - 0x7f
      13'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0
      13'h5F9: dout  = 8'b00010100; // 1529 :  20 - 0x14
      13'h5FA: dout  = 8'b00011100; // 1530 :  28 - 0x1c
      13'h5FB: dout  = 8'b00011100; // 1531 :  28 - 0x1c
      13'h5FC: dout  = 8'b00011100; // 1532 :  28 - 0x1c
      13'h5FD: dout  = 8'b00011100; // 1533 :  28 - 0x1c
      13'h5FE: dout  = 8'b00011100; // 1534 :  28 - 0x1c
      13'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      13'h600: dout  = 8'b11111111; // 1536 : 255 - 0xff -- Sprite 0x60
      13'h601: dout  = 8'b11111111; // 1537 : 255 - 0xff
      13'h602: dout  = 8'b11111111; // 1538 : 255 - 0xff
      13'h603: dout  = 8'b11111111; // 1539 : 255 - 0xff
      13'h604: dout  = 8'b11010101; // 1540 : 213 - 0xd5
      13'h605: dout  = 8'b10101010; // 1541 : 170 - 0xaa
      13'h606: dout  = 8'b11010101; // 1542 : 213 - 0xd5
      13'h607: dout  = 8'b11111111; // 1543 : 255 - 0xff
      13'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout  = 8'b01111111; // 1545 : 127 - 0x7f
      13'h60A: dout  = 8'b01111111; // 1546 : 127 - 0x7f
      13'h60B: dout  = 8'b01111111; // 1547 : 127 - 0x7f
      13'h60C: dout  = 8'b01111111; // 1548 : 127 - 0x7f
      13'h60D: dout  = 8'b01111111; // 1549 : 127 - 0x7f
      13'h60E: dout  = 8'b00101010; // 1550 :  42 - 0x2a
      13'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      13'h610: dout  = 8'b11111111; // 1552 : 255 - 0xff -- Sprite 0x61
      13'h611: dout  = 8'b11111111; // 1553 : 255 - 0xff
      13'h612: dout  = 8'b11111111; // 1554 : 255 - 0xff
      13'h613: dout  = 8'b11111111; // 1555 : 255 - 0xff
      13'h614: dout  = 8'b01010101; // 1556 :  85 - 0x55
      13'h615: dout  = 8'b10101010; // 1557 : 170 - 0xaa
      13'h616: dout  = 8'b01010101; // 1558 :  85 - 0x55
      13'h617: dout  = 8'b11111111; // 1559 : 255 - 0xff
      13'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0
      13'h619: dout  = 8'b11111111; // 1561 : 255 - 0xff
      13'h61A: dout  = 8'b11111111; // 1562 : 255 - 0xff
      13'h61B: dout  = 8'b11111111; // 1563 : 255 - 0xff
      13'h61C: dout  = 8'b11111111; // 1564 : 255 - 0xff
      13'h61D: dout  = 8'b11111111; // 1565 : 255 - 0xff
      13'h61E: dout  = 8'b10101010; // 1566 : 170 - 0xaa
      13'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      13'h620: dout  = 8'b11111111; // 1568 : 255 - 0xff -- Sprite 0x62
      13'h621: dout  = 8'b11111111; // 1569 : 255 - 0xff
      13'h622: dout  = 8'b11111111; // 1570 : 255 - 0xff
      13'h623: dout  = 8'b11111111; // 1571 : 255 - 0xff
      13'h624: dout  = 8'b01010101; // 1572 :  85 - 0x55
      13'h625: dout  = 8'b10101011; // 1573 : 171 - 0xab
      13'h626: dout  = 8'b01010101; // 1574 :  85 - 0x55
      13'h627: dout  = 8'b11111111; // 1575 : 255 - 0xff
      13'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0
      13'h629: dout  = 8'b11111110; // 1577 : 254 - 0xfe
      13'h62A: dout  = 8'b11111110; // 1578 : 254 - 0xfe
      13'h62B: dout  = 8'b11111110; // 1579 : 254 - 0xfe
      13'h62C: dout  = 8'b11111110; // 1580 : 254 - 0xfe
      13'h62D: dout  = 8'b11111110; // 1581 : 254 - 0xfe
      13'h62E: dout  = 8'b10101010; // 1582 : 170 - 0xaa
      13'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0x63
      13'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      13'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      13'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      13'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      13'h635: dout  = 8'b00000000; // 1589 :   0 - 0x0
      13'h636: dout  = 8'b00000000; // 1590 :   0 - 0x0
      13'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      13'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0
      13'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      13'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      13'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      13'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      13'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      13'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      13'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout  = 8'b00000001; // 1600 :   1 - 0x1 -- Sprite 0x64
      13'h641: dout  = 8'b00000001; // 1601 :   1 - 0x1
      13'h642: dout  = 8'b00000011; // 1602 :   3 - 0x3
      13'h643: dout  = 8'b00000011; // 1603 :   3 - 0x3
      13'h644: dout  = 8'b00000110; // 1604 :   6 - 0x6
      13'h645: dout  = 8'b00000110; // 1605 :   6 - 0x6
      13'h646: dout  = 8'b00001100; // 1606 :  12 - 0xc
      13'h647: dout  = 8'b00001100; // 1607 :  12 - 0xc
      13'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      13'h64A: dout  = 8'b00000001; // 1610 :   1 - 0x1
      13'h64B: dout  = 8'b00000001; // 1611 :   1 - 0x1
      13'h64C: dout  = 8'b00000011; // 1612 :   3 - 0x3
      13'h64D: dout  = 8'b00000011; // 1613 :   3 - 0x3
      13'h64E: dout  = 8'b00000111; // 1614 :   7 - 0x7
      13'h64F: dout  = 8'b00000111; // 1615 :   7 - 0x7
      13'h650: dout  = 8'b00011000; // 1616 :  24 - 0x18 -- Sprite 0x65
      13'h651: dout  = 8'b00011000; // 1617 :  24 - 0x18
      13'h652: dout  = 8'b00110000; // 1618 :  48 - 0x30
      13'h653: dout  = 8'b00110000; // 1619 :  48 - 0x30
      13'h654: dout  = 8'b01100000; // 1620 :  96 - 0x60
      13'h655: dout  = 8'b01100000; // 1621 :  96 - 0x60
      13'h656: dout  = 8'b11101010; // 1622 : 234 - 0xea
      13'h657: dout  = 8'b11111111; // 1623 : 255 - 0xff
      13'h658: dout  = 8'b00001111; // 1624 :  15 - 0xf
      13'h659: dout  = 8'b00001111; // 1625 :  15 - 0xf
      13'h65A: dout  = 8'b00011111; // 1626 :  31 - 0x1f
      13'h65B: dout  = 8'b00011111; // 1627 :  31 - 0x1f
      13'h65C: dout  = 8'b00111111; // 1628 :  63 - 0x3f
      13'h65D: dout  = 8'b00111111; // 1629 :  63 - 0x3f
      13'h65E: dout  = 8'b01010101; // 1630 :  85 - 0x55
      13'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout  = 8'b10000000; // 1632 : 128 - 0x80 -- Sprite 0x66
      13'h661: dout  = 8'b10000000; // 1633 : 128 - 0x80
      13'h662: dout  = 8'b11000000; // 1634 : 192 - 0xc0
      13'h663: dout  = 8'b01000000; // 1635 :  64 - 0x40
      13'h664: dout  = 8'b10100000; // 1636 : 160 - 0xa0
      13'h665: dout  = 8'b01100000; // 1637 :  96 - 0x60
      13'h666: dout  = 8'b00110000; // 1638 :  48 - 0x30
      13'h667: dout  = 8'b00010000; // 1639 :  16 - 0x10
      13'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      13'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      13'h66B: dout  = 8'b10000000; // 1643 : 128 - 0x80
      13'h66C: dout  = 8'b01000000; // 1644 :  64 - 0x40
      13'h66D: dout  = 8'b10000000; // 1645 : 128 - 0x80
      13'h66E: dout  = 8'b11000000; // 1646 : 192 - 0xc0
      13'h66F: dout  = 8'b11100000; // 1647 : 224 - 0xe0
      13'h670: dout  = 8'b00101000; // 1648 :  40 - 0x28 -- Sprite 0x67
      13'h671: dout  = 8'b00011000; // 1649 :  24 - 0x18
      13'h672: dout  = 8'b00001100; // 1650 :  12 - 0xc
      13'h673: dout  = 8'b00010100; // 1651 :  20 - 0x14
      13'h674: dout  = 8'b00001010; // 1652 :  10 - 0xa
      13'h675: dout  = 8'b00000110; // 1653 :   6 - 0x6
      13'h676: dout  = 8'b10101011; // 1654 : 171 - 0xab
      13'h677: dout  = 8'b11111111; // 1655 : 255 - 0xff
      13'h678: dout  = 8'b11010000; // 1656 : 208 - 0xd0
      13'h679: dout  = 8'b11100000; // 1657 : 224 - 0xe0
      13'h67A: dout  = 8'b11110000; // 1658 : 240 - 0xf0
      13'h67B: dout  = 8'b11101000; // 1659 : 232 - 0xe8
      13'h67C: dout  = 8'b11110100; // 1660 : 244 - 0xf4
      13'h67D: dout  = 8'b11111000; // 1661 : 248 - 0xf8
      13'h67E: dout  = 8'b01010100; // 1662 :  84 - 0x54
      13'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      13'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      13'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      13'h684: dout  = 8'b00000000; // 1668 :   0 - 0x0
      13'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      13'h686: dout  = 8'b00000000; // 1670 :   0 - 0x0
      13'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      13'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      13'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      13'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      13'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      13'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      13'h68E: dout  = 8'b00000000; // 1678 :   0 - 0x0
      13'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      13'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      13'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      13'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      13'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      13'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      13'h695: dout  = 8'b00000000; // 1685 :   0 - 0x0
      13'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      13'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      13'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout  = 8'b00000000; // 1689 :   0 - 0x0
      13'h69A: dout  = 8'b00000000; // 1690 :   0 - 0x0
      13'h69B: dout  = 8'b00000000; // 1691 :   0 - 0x0
      13'h69C: dout  = 8'b00000000; // 1692 :   0 - 0x0
      13'h69D: dout  = 8'b00000000; // 1693 :   0 - 0x0
      13'h69E: dout  = 8'b00000000; // 1694 :   0 - 0x0
      13'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      13'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      13'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      13'h6A4: dout  = 8'b00000000; // 1700 :   0 - 0x0
      13'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      13'h6A6: dout  = 8'b00000000; // 1702 :   0 - 0x0
      13'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      13'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0
      13'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      13'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      13'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      13'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      13'h6AD: dout  = 8'b00000000; // 1709 :   0 - 0x0
      13'h6AE: dout  = 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      13'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      13'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      13'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      13'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      13'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      13'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      13'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      13'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0
      13'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      13'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      13'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      13'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      13'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      13'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      13'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      13'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      13'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      13'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      13'h6C4: dout  = 8'b00000000; // 1732 :   0 - 0x0
      13'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      13'h6C6: dout  = 8'b00000000; // 1734 :   0 - 0x0
      13'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      13'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0
      13'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      13'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      13'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      13'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      13'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      13'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      13'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      13'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      13'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      13'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      13'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      13'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      13'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      13'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      13'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout  = 8'b00000000; // 1753 :   0 - 0x0
      13'h6DA: dout  = 8'b00000000; // 1754 :   0 - 0x0
      13'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      13'h6DC: dout  = 8'b00000000; // 1756 :   0 - 0x0
      13'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      13'h6DE: dout  = 8'b00000000; // 1758 :   0 - 0x0
      13'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      13'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      13'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      13'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      13'h6E6: dout  = 8'b00000000; // 1766 :   0 - 0x0
      13'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      13'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0
      13'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      13'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      13'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      13'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      13'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      13'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0x6f
      13'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      13'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      13'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      13'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      13'h6F5: dout  = 8'b00000000; // 1781 :   0 - 0x0
      13'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      13'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      13'h6F8: dout  = 8'b00000000; // 1784 :   0 - 0x0
      13'h6F9: dout  = 8'b00000000; // 1785 :   0 - 0x0
      13'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      13'h6FB: dout  = 8'b00000000; // 1787 :   0 - 0x0
      13'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      13'h6FD: dout  = 8'b00000000; // 1789 :   0 - 0x0
      13'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      13'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      13'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      13'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      13'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      13'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      13'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      13'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      13'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0
      13'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      13'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      13'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      13'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      13'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      13'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      13'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      13'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0x71
      13'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      13'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      13'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      13'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      13'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      13'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      13'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      13'h718: dout  = 8'b00000000; // 1816 :   0 - 0x0
      13'h719: dout  = 8'b00000000; // 1817 :   0 - 0x0
      13'h71A: dout  = 8'b00000000; // 1818 :   0 - 0x0
      13'h71B: dout  = 8'b00000000; // 1819 :   0 - 0x0
      13'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      13'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      13'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      13'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      13'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0x72
      13'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      13'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      13'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      13'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      13'h725: dout  = 8'b00000000; // 1829 :   0 - 0x0
      13'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      13'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      13'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0
      13'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      13'h72A: dout  = 8'b00000000; // 1834 :   0 - 0x0
      13'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      13'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      13'h72D: dout  = 8'b00000000; // 1837 :   0 - 0x0
      13'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      13'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      13'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0x73
      13'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      13'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      13'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      13'h734: dout  = 8'b00000000; // 1844 :   0 - 0x0
      13'h735: dout  = 8'b00000000; // 1845 :   0 - 0x0
      13'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      13'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      13'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0
      13'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      13'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      13'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      13'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      13'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      13'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      13'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      13'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      13'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      13'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      13'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      13'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      13'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      13'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      13'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      13'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0
      13'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      13'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      13'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      13'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      13'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      13'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      13'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      13'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      13'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      13'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      13'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      13'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      13'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      13'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      13'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      13'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0
      13'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      13'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      13'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      13'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      13'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      13'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      13'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      13'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0x76
      13'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      13'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      13'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      13'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      13'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      13'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      13'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      13'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0
      13'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      13'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      13'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      13'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      13'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      13'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      13'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      13'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0x77
      13'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      13'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      13'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      13'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      13'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      13'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      13'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      13'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0
      13'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      13'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      13'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      13'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      13'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      13'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      13'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      13'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      13'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      13'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      13'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      13'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      13'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      13'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      13'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      13'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0
      13'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      13'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      13'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      13'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      13'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      13'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      13'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      13'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      13'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      13'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      13'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      13'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      13'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      13'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      13'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      13'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0
      13'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      13'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      13'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      13'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      13'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      13'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      13'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      13'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      13'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      13'h7A2: dout  = 8'b00000000; // 1954 :   0 - 0x0
      13'h7A3: dout  = 8'b00000000; // 1955 :   0 - 0x0
      13'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      13'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      13'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      13'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      13'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0
      13'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      13'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      13'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      13'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      13'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      13'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      13'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      13'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      13'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      13'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      13'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      13'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      13'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      13'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      13'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      13'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0
      13'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      13'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      13'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      13'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      13'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      13'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      13'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      13'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      13'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      13'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      13'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      13'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      13'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      13'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      13'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      13'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      13'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      13'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      13'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      13'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      13'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      13'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      13'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      13'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      13'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      13'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      13'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      13'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      13'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      13'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      13'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0
      13'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      13'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      13'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      13'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      13'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      13'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      13'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      13'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      13'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      13'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      13'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      13'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      13'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      13'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      13'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0
      13'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      13'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      13'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      13'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      13'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      13'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      13'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      13'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      13'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      13'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      13'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      13'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      13'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      13'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      13'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      13'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0
      13'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      13'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      13'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      13'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      13'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      13'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      13'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
      13'h800: dout  = 8'b00000011; // 2048 :   3 - 0x3 -- Sprite 0x80
      13'h801: dout  = 8'b00001111; // 2049 :  15 - 0xf
      13'h802: dout  = 8'b00011100; // 2050 :  28 - 0x1c
      13'h803: dout  = 8'b00110000; // 2051 :  48 - 0x30
      13'h804: dout  = 8'b00100000; // 2052 :  32 - 0x20
      13'h805: dout  = 8'b01000000; // 2053 :  64 - 0x40
      13'h806: dout  = 8'b01000000; // 2054 :  64 - 0x40
      13'h807: dout  = 8'b01111111; // 2055 : 127 - 0x7f
      13'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0
      13'h809: dout  = 8'b00000011; // 2057 :   3 - 0x3
      13'h80A: dout  = 8'b00001111; // 2058 :  15 - 0xf
      13'h80B: dout  = 8'b00011111; // 2059 :  31 - 0x1f
      13'h80C: dout  = 8'b00011111; // 2060 :  31 - 0x1f
      13'h80D: dout  = 8'b00111111; // 2061 :  63 - 0x3f
      13'h80E: dout  = 8'b00111111; // 2062 :  63 - 0x3f
      13'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      13'h810: dout  = 8'b00000001; // 2064 :   1 - 0x1 -- Sprite 0x81
      13'h811: dout  = 8'b00000001; // 2065 :   1 - 0x1
      13'h812: dout  = 8'b00000001; // 2066 :   1 - 0x1
      13'h813: dout  = 8'b00000001; // 2067 :   1 - 0x1
      13'h814: dout  = 8'b00000001; // 2068 :   1 - 0x1
      13'h815: dout  = 8'b00000001; // 2069 :   1 - 0x1
      13'h816: dout  = 8'b00000011; // 2070 :   3 - 0x3
      13'h817: dout  = 8'b00000011; // 2071 :   3 - 0x3
      13'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0
      13'h819: dout  = 8'b00000000; // 2073 :   0 - 0x0
      13'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      13'h81B: dout  = 8'b00000000; // 2075 :   0 - 0x0
      13'h81C: dout  = 8'b00000000; // 2076 :   0 - 0x0
      13'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      13'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      13'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      13'h820: dout  = 8'b11000000; // 2080 : 192 - 0xc0 -- Sprite 0x82
      13'h821: dout  = 8'b11110000; // 2081 : 240 - 0xf0
      13'h822: dout  = 8'b00111000; // 2082 :  56 - 0x38
      13'h823: dout  = 8'b00001110; // 2083 :  14 - 0xe
      13'h824: dout  = 8'b00011110; // 2084 :  30 - 0x1e
      13'h825: dout  = 8'b00011110; // 2085 :  30 - 0x1e
      13'h826: dout  = 8'b00000010; // 2086 :   2 - 0x2
      13'h827: dout  = 8'b11111110; // 2087 : 254 - 0xfe
      13'h828: dout  = 8'b00000000; // 2088 :   0 - 0x0
      13'h829: dout  = 8'b11000000; // 2089 : 192 - 0xc0
      13'h82A: dout  = 8'b11110000; // 2090 : 240 - 0xf0
      13'h82B: dout  = 8'b11110000; // 2091 : 240 - 0xf0
      13'h82C: dout  = 8'b11101100; // 2092 : 236 - 0xec
      13'h82D: dout  = 8'b11100000; // 2093 : 224 - 0xe0
      13'h82E: dout  = 8'b11111100; // 2094 : 252 - 0xfc
      13'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      13'h830: dout  = 8'b10000000; // 2096 : 128 - 0x80 -- Sprite 0x83
      13'h831: dout  = 8'b10000000; // 2097 : 128 - 0x80
      13'h832: dout  = 8'b10000000; // 2098 : 128 - 0x80
      13'h833: dout  = 8'b10000000; // 2099 : 128 - 0x80
      13'h834: dout  = 8'b10000000; // 2100 : 128 - 0x80
      13'h835: dout  = 8'b11100000; // 2101 : 224 - 0xe0
      13'h836: dout  = 8'b00010000; // 2102 :  16 - 0x10
      13'h837: dout  = 8'b11110000; // 2103 : 240 - 0xf0
      13'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0
      13'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      13'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      13'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      13'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      13'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      13'h83E: dout  = 8'b11100000; // 2110 : 224 - 0xe0
      13'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      13'h840: dout  = 8'b00000011; // 2112 :   3 - 0x3 -- Sprite 0x84
      13'h841: dout  = 8'b00001111; // 2113 :  15 - 0xf
      13'h842: dout  = 8'b00011100; // 2114 :  28 - 0x1c
      13'h843: dout  = 8'b00110000; // 2115 :  48 - 0x30
      13'h844: dout  = 8'b00100000; // 2116 :  32 - 0x20
      13'h845: dout  = 8'b01000000; // 2117 :  64 - 0x40
      13'h846: dout  = 8'b01000000; // 2118 :  64 - 0x40
      13'h847: dout  = 8'b01111111; // 2119 : 127 - 0x7f
      13'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0
      13'h849: dout  = 8'b00000011; // 2121 :   3 - 0x3
      13'h84A: dout  = 8'b00001111; // 2122 :  15 - 0xf
      13'h84B: dout  = 8'b00011111; // 2123 :  31 - 0x1f
      13'h84C: dout  = 8'b00011111; // 2124 :  31 - 0x1f
      13'h84D: dout  = 8'b00111111; // 2125 :  63 - 0x3f
      13'h84E: dout  = 8'b00111111; // 2126 :  63 - 0x3f
      13'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      13'h850: dout  = 8'b00000011; // 2128 :   3 - 0x3 -- Sprite 0x85
      13'h851: dout  = 8'b00000110; // 2129 :   6 - 0x6
      13'h852: dout  = 8'b00000110; // 2130 :   6 - 0x6
      13'h853: dout  = 8'b00011100; // 2131 :  28 - 0x1c
      13'h854: dout  = 8'b00011000; // 2132 :  24 - 0x18
      13'h855: dout  = 8'b00110110; // 2133 :  54 - 0x36
      13'h856: dout  = 8'b00110001; // 2134 :  49 - 0x31
      13'h857: dout  = 8'b00001111; // 2135 :  15 - 0xf
      13'h858: dout  = 8'b00000000; // 2136 :   0 - 0x0
      13'h859: dout  = 8'b00000000; // 2137 :   0 - 0x0
      13'h85A: dout  = 8'b00000000; // 2138 :   0 - 0x0
      13'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      13'h85C: dout  = 8'b00000000; // 2140 :   0 - 0x0
      13'h85D: dout  = 8'b00001000; // 2141 :   8 - 0x8
      13'h85E: dout  = 8'b00001110; // 2142 :  14 - 0xe
      13'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      13'h860: dout  = 8'b11000000; // 2144 : 192 - 0xc0 -- Sprite 0x86
      13'h861: dout  = 8'b11110000; // 2145 : 240 - 0xf0
      13'h862: dout  = 8'b00111000; // 2146 :  56 - 0x38
      13'h863: dout  = 8'b00001110; // 2147 :  14 - 0xe
      13'h864: dout  = 8'b00011110; // 2148 :  30 - 0x1e
      13'h865: dout  = 8'b00011110; // 2149 :  30 - 0x1e
      13'h866: dout  = 8'b00000010; // 2150 :   2 - 0x2
      13'h867: dout  = 8'b11111110; // 2151 : 254 - 0xfe
      13'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0
      13'h869: dout  = 8'b11000000; // 2153 : 192 - 0xc0
      13'h86A: dout  = 8'b11110000; // 2154 : 240 - 0xf0
      13'h86B: dout  = 8'b11110000; // 2155 : 240 - 0xf0
      13'h86C: dout  = 8'b11101100; // 2156 : 236 - 0xec
      13'h86D: dout  = 8'b11100000; // 2157 : 224 - 0xe0
      13'h86E: dout  = 8'b11111100; // 2158 : 252 - 0xfc
      13'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      13'h870: dout  = 8'b11000000; // 2160 : 192 - 0xc0 -- Sprite 0x87
      13'h871: dout  = 8'b01100000; // 2161 :  96 - 0x60
      13'h872: dout  = 8'b01100000; // 2162 :  96 - 0x60
      13'h873: dout  = 8'b00110000; // 2163 :  48 - 0x30
      13'h874: dout  = 8'b00111110; // 2164 :  62 - 0x3e
      13'h875: dout  = 8'b00011001; // 2165 :  25 - 0x19
      13'h876: dout  = 8'b00110011; // 2166 :  51 - 0x33
      13'h877: dout  = 8'b00111100; // 2167 :  60 - 0x3c
      13'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0
      13'h879: dout  = 8'b00000000; // 2169 :   0 - 0x0
      13'h87A: dout  = 8'b00000000; // 2170 :   0 - 0x0
      13'h87B: dout  = 8'b00000000; // 2171 :   0 - 0x0
      13'h87C: dout  = 8'b00000000; // 2172 :   0 - 0x0
      13'h87D: dout  = 8'b00000110; // 2173 :   6 - 0x6
      13'h87E: dout  = 8'b00001100; // 2174 :  12 - 0xc
      13'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      13'h880: dout  = 8'b00000011; // 2176 :   3 - 0x3 -- Sprite 0x88
      13'h881: dout  = 8'b00000111; // 2177 :   7 - 0x7
      13'h882: dout  = 8'b00000111; // 2178 :   7 - 0x7
      13'h883: dout  = 8'b00001011; // 2179 :  11 - 0xb
      13'h884: dout  = 8'b00010000; // 2180 :  16 - 0x10
      13'h885: dout  = 8'b01100000; // 2181 :  96 - 0x60
      13'h886: dout  = 8'b11110000; // 2182 : 240 - 0xf0
      13'h887: dout  = 8'b11110000; // 2183 : 240 - 0xf0
      13'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout  = 8'b00000011; // 2185 :   3 - 0x3
      13'h88A: dout  = 8'b00000011; // 2186 :   3 - 0x3
      13'h88B: dout  = 8'b00000100; // 2187 :   4 - 0x4
      13'h88C: dout  = 8'b00001111; // 2188 :  15 - 0xf
      13'h88D: dout  = 8'b00011111; // 2189 :  31 - 0x1f
      13'h88E: dout  = 8'b01101111; // 2190 : 111 - 0x6f
      13'h88F: dout  = 8'b01101111; // 2191 : 111 - 0x6f
      13'h890: dout  = 8'b11110000; // 2192 : 240 - 0xf0 -- Sprite 0x89
      13'h891: dout  = 8'b11110000; // 2193 : 240 - 0xf0
      13'h892: dout  = 8'b01100000; // 2194 :  96 - 0x60
      13'h893: dout  = 8'b00010000; // 2195 :  16 - 0x10
      13'h894: dout  = 8'b00001011; // 2196 :  11 - 0xb
      13'h895: dout  = 8'b00000111; // 2197 :   7 - 0x7
      13'h896: dout  = 8'b00000111; // 2198 :   7 - 0x7
      13'h897: dout  = 8'b00000011; // 2199 :   3 - 0x3
      13'h898: dout  = 8'b01101111; // 2200 : 111 - 0x6f
      13'h899: dout  = 8'b01101111; // 2201 : 111 - 0x6f
      13'h89A: dout  = 8'b00011111; // 2202 :  31 - 0x1f
      13'h89B: dout  = 8'b00001111; // 2203 :  15 - 0xf
      13'h89C: dout  = 8'b00000100; // 2204 :   4 - 0x4
      13'h89D: dout  = 8'b00000011; // 2205 :   3 - 0x3
      13'h89E: dout  = 8'b00000011; // 2206 :   3 - 0x3
      13'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      13'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Sprite 0x8a
      13'h8A1: dout  = 8'b00011100; // 2209 :  28 - 0x1c
      13'h8A2: dout  = 8'b00111111; // 2210 :  63 - 0x3f
      13'h8A3: dout  = 8'b01111000; // 2211 : 120 - 0x78
      13'h8A4: dout  = 8'b01110000; // 2212 : 112 - 0x70
      13'h8A5: dout  = 8'b01100000; // 2213 :  96 - 0x60
      13'h8A6: dout  = 8'b00100000; // 2214 :  32 - 0x20
      13'h8A7: dout  = 8'b00100000; // 2215 :  32 - 0x20
      13'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      13'h8AA: dout  = 8'b00011000; // 2218 :  24 - 0x18
      13'h8AB: dout  = 8'b00110111; // 2219 :  55 - 0x37
      13'h8AC: dout  = 8'b00101111; // 2220 :  47 - 0x2f
      13'h8AD: dout  = 8'b00011111; // 2221 :  31 - 0x1f
      13'h8AE: dout  = 8'b00011111; // 2222 :  31 - 0x1f
      13'h8AF: dout  = 8'b00011111; // 2223 :  31 - 0x1f
      13'h8B0: dout  = 8'b00100000; // 2224 :  32 - 0x20 -- Sprite 0x8b
      13'h8B1: dout  = 8'b00100000; // 2225 :  32 - 0x20
      13'h8B2: dout  = 8'b01100000; // 2226 :  96 - 0x60
      13'h8B3: dout  = 8'b01110000; // 2227 : 112 - 0x70
      13'h8B4: dout  = 8'b01111000; // 2228 : 120 - 0x78
      13'h8B5: dout  = 8'b00111111; // 2229 :  63 - 0x3f
      13'h8B6: dout  = 8'b00011100; // 2230 :  28 - 0x1c
      13'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      13'h8B8: dout  = 8'b00011111; // 2232 :  31 - 0x1f
      13'h8B9: dout  = 8'b00011111; // 2233 :  31 - 0x1f
      13'h8BA: dout  = 8'b00011111; // 2234 :  31 - 0x1f
      13'h8BB: dout  = 8'b00101111; // 2235 :  47 - 0x2f
      13'h8BC: dout  = 8'b00110111; // 2236 :  55 - 0x37
      13'h8BD: dout  = 8'b00011000; // 2237 :  24 - 0x18
      13'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      13'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      13'h8C0: dout  = 8'b00000011; // 2240 :   3 - 0x3 -- Sprite 0x8c
      13'h8C1: dout  = 8'b00001100; // 2241 :  12 - 0xc
      13'h8C2: dout  = 8'b00011110; // 2242 :  30 - 0x1e
      13'h8C3: dout  = 8'b00100110; // 2243 :  38 - 0x26
      13'h8C4: dout  = 8'b01000110; // 2244 :  70 - 0x46
      13'h8C5: dout  = 8'b01100100; // 2245 : 100 - 0x64
      13'h8C6: dout  = 8'b01110000; // 2246 : 112 - 0x70
      13'h8C7: dout  = 8'b11110000; // 2247 : 240 - 0xf0
      13'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout  = 8'b00000011; // 2249 :   3 - 0x3
      13'h8CA: dout  = 8'b00000001; // 2250 :   1 - 0x1
      13'h8CB: dout  = 8'b00011001; // 2251 :  25 - 0x19
      13'h8CC: dout  = 8'b00111001; // 2252 :  57 - 0x39
      13'h8CD: dout  = 8'b00011011; // 2253 :  27 - 0x1b
      13'h8CE: dout  = 8'b00001111; // 2254 :  15 - 0xf
      13'h8CF: dout  = 8'b00001111; // 2255 :  15 - 0xf
      13'h8D0: dout  = 8'b10101010; // 2256 : 170 - 0xaa -- Sprite 0x8d
      13'h8D1: dout  = 8'b11111111; // 2257 : 255 - 0xff
      13'h8D2: dout  = 8'b01111111; // 2258 : 127 - 0x7f
      13'h8D3: dout  = 8'b00111001; // 2259 :  57 - 0x39
      13'h8D4: dout  = 8'b00011001; // 2260 :  25 - 0x19
      13'h8D5: dout  = 8'b00001011; // 2261 :  11 - 0xb
      13'h8D6: dout  = 8'b00001000; // 2262 :   8 - 0x8
      13'h8D7: dout  = 8'b00000111; // 2263 :   7 - 0x7
      13'h8D8: dout  = 8'b01111111; // 2264 : 127 - 0x7f
      13'h8D9: dout  = 8'b01111111; // 2265 : 127 - 0x7f
      13'h8DA: dout  = 8'b00111111; // 2266 :  63 - 0x3f
      13'h8DB: dout  = 8'b00010111; // 2267 :  23 - 0x17
      13'h8DC: dout  = 8'b00000110; // 2268 :   6 - 0x6
      13'h8DD: dout  = 8'b00000100; // 2269 :   4 - 0x4
      13'h8DE: dout  = 8'b00000111; // 2270 :   7 - 0x7
      13'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      13'h8E0: dout  = 8'b11000000; // 2272 : 192 - 0xc0 -- Sprite 0x8e
      13'h8E1: dout  = 8'b00110000; // 2273 :  48 - 0x30
      13'h8E2: dout  = 8'b00001000; // 2274 :   8 - 0x8
      13'h8E3: dout  = 8'b01000100; // 2275 :  68 - 0x44
      13'h8E4: dout  = 8'b01100010; // 2276 :  98 - 0x62
      13'h8E5: dout  = 8'b01100010; // 2277 :  98 - 0x62
      13'h8E6: dout  = 8'b00000001; // 2278 :   1 - 0x1
      13'h8E7: dout  = 8'b00111111; // 2279 :  63 - 0x3f
      13'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0
      13'h8E9: dout  = 8'b11000000; // 2281 : 192 - 0xc0
      13'h8EA: dout  = 8'b11110000; // 2282 : 240 - 0xf0
      13'h8EB: dout  = 8'b10111000; // 2283 : 184 - 0xb8
      13'h8EC: dout  = 8'b10011100; // 2284 : 156 - 0x9c
      13'h8ED: dout  = 8'b11111100; // 2285 : 252 - 0xfc
      13'h8EE: dout  = 8'b11111110; // 2286 : 254 - 0xfe
      13'h8EF: dout  = 8'b11000000; // 2287 : 192 - 0xc0
      13'h8F0: dout  = 8'b10001011; // 2288 : 139 - 0x8b -- Sprite 0x8f
      13'h8F1: dout  = 8'b11000001; // 2289 : 193 - 0xc1
      13'h8F2: dout  = 8'b11111110; // 2290 : 254 - 0xfe
      13'h8F3: dout  = 8'b11111100; // 2291 : 252 - 0xfc
      13'h8F4: dout  = 8'b11110000; // 2292 : 240 - 0xf0
      13'h8F5: dout  = 8'b11110000; // 2293 : 240 - 0xf0
      13'h8F6: dout  = 8'b11111000; // 2294 : 248 - 0xf8
      13'h8F7: dout  = 8'b11110000; // 2295 : 240 - 0xf0
      13'h8F8: dout  = 8'b11111110; // 2296 : 254 - 0xfe
      13'h8F9: dout  = 8'b11111110; // 2297 : 254 - 0xfe
      13'h8FA: dout  = 8'b11111000; // 2298 : 248 - 0xf8
      13'h8FB: dout  = 8'b11110000; // 2299 : 240 - 0xf0
      13'h8FC: dout  = 8'b11000000; // 2300 : 192 - 0xc0
      13'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      13'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      13'h8FF: dout  = 8'b10000000; // 2303 : 128 - 0x80
      13'h900: dout  = 8'b00000011; // 2304 :   3 - 0x3 -- Sprite 0x90
      13'h901: dout  = 8'b00001110; // 2305 :  14 - 0xe
      13'h902: dout  = 8'b00010110; // 2306 :  22 - 0x16
      13'h903: dout  = 8'b00100110; // 2307 :  38 - 0x26
      13'h904: dout  = 8'b01100011; // 2308 :  99 - 0x63
      13'h905: dout  = 8'b01110010; // 2309 : 114 - 0x72
      13'h906: dout  = 8'b01110000; // 2310 : 112 - 0x70
      13'h907: dout  = 8'b11010000; // 2311 : 208 - 0xd0
      13'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout  = 8'b00000001; // 2313 :   1 - 0x1
      13'h90A: dout  = 8'b00001001; // 2314 :   9 - 0x9
      13'h90B: dout  = 8'b00011001; // 2315 :  25 - 0x19
      13'h90C: dout  = 8'b00011100; // 2316 :  28 - 0x1c
      13'h90D: dout  = 8'b00001101; // 2317 :  13 - 0xd
      13'h90E: dout  = 8'b00001111; // 2318 :  15 - 0xf
      13'h90F: dout  = 8'b00101111; // 2319 :  47 - 0x2f
      13'h910: dout  = 8'b10101010; // 2320 : 170 - 0xaa -- Sprite 0x91
      13'h911: dout  = 8'b11111111; // 2321 : 255 - 0xff
      13'h912: dout  = 8'b01111111; // 2322 : 127 - 0x7f
      13'h913: dout  = 8'b00111100; // 2323 :  60 - 0x3c
      13'h914: dout  = 8'b00011100; // 2324 :  28 - 0x1c
      13'h915: dout  = 8'b00000100; // 2325 :   4 - 0x4
      13'h916: dout  = 8'b00000010; // 2326 :   2 - 0x2
      13'h917: dout  = 8'b00000001; // 2327 :   1 - 0x1
      13'h918: dout  = 8'b01111111; // 2328 : 127 - 0x7f
      13'h919: dout  = 8'b01111111; // 2329 : 127 - 0x7f
      13'h91A: dout  = 8'b00111111; // 2330 :  63 - 0x3f
      13'h91B: dout  = 8'b00011011; // 2331 :  27 - 0x1b
      13'h91C: dout  = 8'b00000011; // 2332 :   3 - 0x3
      13'h91D: dout  = 8'b00000011; // 2333 :   3 - 0x3
      13'h91E: dout  = 8'b00000001; // 2334 :   1 - 0x1
      13'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout  = 8'b11000000; // 2336 : 192 - 0xc0 -- Sprite 0x92
      13'h921: dout  = 8'b00110000; // 2337 :  48 - 0x30
      13'h922: dout  = 8'b00001000; // 2338 :   8 - 0x8
      13'h923: dout  = 8'b00100100; // 2339 :  36 - 0x24
      13'h924: dout  = 8'b00110010; // 2340 :  50 - 0x32
      13'h925: dout  = 8'b00110010; // 2341 :  50 - 0x32
      13'h926: dout  = 8'b00000001; // 2342 :   1 - 0x1
      13'h927: dout  = 8'b00011111; // 2343 :  31 - 0x1f
      13'h928: dout  = 8'b00000000; // 2344 :   0 - 0x0
      13'h929: dout  = 8'b11000000; // 2345 : 192 - 0xc0
      13'h92A: dout  = 8'b11110000; // 2346 : 240 - 0xf0
      13'h92B: dout  = 8'b11011000; // 2347 : 216 - 0xd8
      13'h92C: dout  = 8'b11001100; // 2348 : 204 - 0xcc
      13'h92D: dout  = 8'b11111100; // 2349 : 252 - 0xfc
      13'h92E: dout  = 8'b11111110; // 2350 : 254 - 0xfe
      13'h92F: dout  = 8'b11100000; // 2351 : 224 - 0xe0
      13'h930: dout  = 8'b10001011; // 2352 : 139 - 0x8b -- Sprite 0x93
      13'h931: dout  = 8'b11000001; // 2353 : 193 - 0xc1
      13'h932: dout  = 8'b11111110; // 2354 : 254 - 0xfe
      13'h933: dout  = 8'b11111100; // 2355 : 252 - 0xfc
      13'h934: dout  = 8'b11110000; // 2356 : 240 - 0xf0
      13'h935: dout  = 8'b11000000; // 2357 : 192 - 0xc0
      13'h936: dout  = 8'b00100000; // 2358 :  32 - 0x20
      13'h937: dout  = 8'b11100000; // 2359 : 224 - 0xe0
      13'h938: dout  = 8'b11111110; // 2360 : 254 - 0xfe
      13'h939: dout  = 8'b11111110; // 2361 : 254 - 0xfe
      13'h93A: dout  = 8'b11111000; // 2362 : 248 - 0xf8
      13'h93B: dout  = 8'b01110000; // 2363 : 112 - 0x70
      13'h93C: dout  = 8'b01000000; // 2364 :  64 - 0x40
      13'h93D: dout  = 8'b00000000; // 2365 :   0 - 0x0
      13'h93E: dout  = 8'b11000000; // 2366 : 192 - 0xc0
      13'h93F: dout  = 8'b00100000; // 2367 :  32 - 0x20
      13'h940: dout  = 8'b00000011; // 2368 :   3 - 0x3 -- Sprite 0x94
      13'h941: dout  = 8'b00001111; // 2369 :  15 - 0xf
      13'h942: dout  = 8'b00010011; // 2370 :  19 - 0x13
      13'h943: dout  = 8'b00110001; // 2371 :  49 - 0x31
      13'h944: dout  = 8'b01111001; // 2372 : 121 - 0x79
      13'h945: dout  = 8'b01011001; // 2373 :  89 - 0x59
      13'h946: dout  = 8'b01001000; // 2374 :  72 - 0x48
      13'h947: dout  = 8'b11001100; // 2375 : 204 - 0xcc
      13'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0
      13'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      13'h94A: dout  = 8'b00001100; // 2378 :  12 - 0xc
      13'h94B: dout  = 8'b00001110; // 2379 :  14 - 0xe
      13'h94C: dout  = 8'b00000110; // 2380 :   6 - 0x6
      13'h94D: dout  = 8'b00100110; // 2381 :  38 - 0x26
      13'h94E: dout  = 8'b00110111; // 2382 :  55 - 0x37
      13'h94F: dout  = 8'b00110011; // 2383 :  51 - 0x33
      13'h950: dout  = 8'b10010101; // 2384 : 149 - 0x95 -- Sprite 0x95
      13'h951: dout  = 8'b11111111; // 2385 : 255 - 0xff
      13'h952: dout  = 8'b01111111; // 2386 : 127 - 0x7f
      13'h953: dout  = 8'b00111110; // 2387 :  62 - 0x3e
      13'h954: dout  = 8'b00011111; // 2388 :  31 - 0x1f
      13'h955: dout  = 8'b00001111; // 2389 :  15 - 0xf
      13'h956: dout  = 8'b00001111; // 2390 :  15 - 0xf
      13'h957: dout  = 8'b00000111; // 2391 :   7 - 0x7
      13'h958: dout  = 8'b01111111; // 2392 : 127 - 0x7f
      13'h959: dout  = 8'b01111111; // 2393 : 127 - 0x7f
      13'h95A: dout  = 8'b00111111; // 2394 :  63 - 0x3f
      13'h95B: dout  = 8'b00011111; // 2395 :  31 - 0x1f
      13'h95C: dout  = 8'b00001110; // 2396 :  14 - 0xe
      13'h95D: dout  = 8'b00000000; // 2397 :   0 - 0x0
      13'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      13'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      13'h960: dout  = 8'b11000000; // 2400 : 192 - 0xc0 -- Sprite 0x96
      13'h961: dout  = 8'b00110000; // 2401 :  48 - 0x30
      13'h962: dout  = 8'b00001000; // 2402 :   8 - 0x8
      13'h963: dout  = 8'b10010100; // 2403 : 148 - 0x94
      13'h964: dout  = 8'b10011010; // 2404 : 154 - 0x9a
      13'h965: dout  = 8'b00011010; // 2405 :  26 - 0x1a
      13'h966: dout  = 8'b00000001; // 2406 :   1 - 0x1
      13'h967: dout  = 8'b00001111; // 2407 :  15 - 0xf
      13'h968: dout  = 8'b00000000; // 2408 :   0 - 0x0
      13'h969: dout  = 8'b11000000; // 2409 : 192 - 0xc0
      13'h96A: dout  = 8'b11110000; // 2410 : 240 - 0xf0
      13'h96B: dout  = 8'b01101000; // 2411 : 104 - 0x68
      13'h96C: dout  = 8'b01100100; // 2412 : 100 - 0x64
      13'h96D: dout  = 8'b11111100; // 2413 : 252 - 0xfc
      13'h96E: dout  = 8'b11111110; // 2414 : 254 - 0xfe
      13'h96F: dout  = 8'b11110000; // 2415 : 240 - 0xf0
      13'h970: dout  = 8'b01000101; // 2416 :  69 - 0x45 -- Sprite 0x97
      13'h971: dout  = 8'b11100001; // 2417 : 225 - 0xe1
      13'h972: dout  = 8'b11111110; // 2418 : 254 - 0xfe
      13'h973: dout  = 8'b01111100; // 2419 : 124 - 0x7c
      13'h974: dout  = 8'b00110000; // 2420 :  48 - 0x30
      13'h975: dout  = 8'b00110000; // 2421 :  48 - 0x30
      13'h976: dout  = 8'b10001000; // 2422 : 136 - 0x88
      13'h977: dout  = 8'b01111000; // 2423 : 120 - 0x78
      13'h978: dout  = 8'b11111111; // 2424 : 255 - 0xff
      13'h979: dout  = 8'b11111110; // 2425 : 254 - 0xfe
      13'h97A: dout  = 8'b11111100; // 2426 : 252 - 0xfc
      13'h97B: dout  = 8'b10110000; // 2427 : 176 - 0xb0
      13'h97C: dout  = 8'b11000000; // 2428 : 192 - 0xc0
      13'h97D: dout  = 8'b11000000; // 2429 : 192 - 0xc0
      13'h97E: dout  = 8'b01110000; // 2430 : 112 - 0x70
      13'h97F: dout  = 8'b00001000; // 2431 :   8 - 0x8
      13'h980: dout  = 8'b00000001; // 2432 :   1 - 0x1 -- Sprite 0x98
      13'h981: dout  = 8'b00000000; // 2433 :   0 - 0x0
      13'h982: dout  = 8'b00000000; // 2434 :   0 - 0x0
      13'h983: dout  = 8'b00000000; // 2435 :   0 - 0x0
      13'h984: dout  = 8'b00000001; // 2436 :   1 - 0x1
      13'h985: dout  = 8'b00000001; // 2437 :   1 - 0x1
      13'h986: dout  = 8'b00000010; // 2438 :   2 - 0x2
      13'h987: dout  = 8'b00000110; // 2439 :   6 - 0x6
      13'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0
      13'h989: dout  = 8'b00000001; // 2441 :   1 - 0x1
      13'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      13'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      13'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      13'h98D: dout  = 8'b00000000; // 2445 :   0 - 0x0
      13'h98E: dout  = 8'b00000001; // 2446 :   1 - 0x1
      13'h98F: dout  = 8'b00000011; // 2447 :   3 - 0x3
      13'h990: dout  = 8'b01111000; // 2448 : 120 - 0x78 -- Sprite 0x99
      13'h991: dout  = 8'b00101010; // 2449 :  42 - 0x2a
      13'h992: dout  = 8'b01010100; // 2450 :  84 - 0x54
      13'h993: dout  = 8'b00101001; // 2451 :  41 - 0x29
      13'h994: dout  = 8'b00101111; // 2452 :  47 - 0x2f
      13'h995: dout  = 8'b00110111; // 2453 :  55 - 0x37
      13'h996: dout  = 8'b00000011; // 2454 :   3 - 0x3
      13'h997: dout  = 8'b00000111; // 2455 :   7 - 0x7
      13'h998: dout  = 8'b00000111; // 2456 :   7 - 0x7
      13'h999: dout  = 8'b00010111; // 2457 :  23 - 0x17
      13'h99A: dout  = 8'b00101111; // 2458 :  47 - 0x2f
      13'h99B: dout  = 8'b00011110; // 2459 :  30 - 0x1e
      13'h99C: dout  = 8'b00010001; // 2460 :  17 - 0x11
      13'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      13'h99E: dout  = 8'b00000001; // 2462 :   1 - 0x1
      13'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout  = 8'b10110000; // 2464 : 176 - 0xb0 -- Sprite 0x9a
      13'h9A1: dout  = 8'b11101000; // 2465 : 232 - 0xe8
      13'h9A2: dout  = 8'b10001100; // 2466 : 140 - 0x8c
      13'h9A3: dout  = 8'b10011110; // 2467 : 158 - 0x9e
      13'h9A4: dout  = 8'b00011111; // 2468 :  31 - 0x1f
      13'h9A5: dout  = 8'b00001111; // 2469 :  15 - 0xf
      13'h9A6: dout  = 8'b10010110; // 2470 : 150 - 0x96
      13'h9A7: dout  = 8'b00011100; // 2471 :  28 - 0x1c
      13'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout  = 8'b00010000; // 2473 :  16 - 0x10
      13'h9AA: dout  = 8'b01111000; // 2474 : 120 - 0x78
      13'h9AB: dout  = 8'b01110100; // 2475 : 116 - 0x74
      13'h9AC: dout  = 8'b11111110; // 2476 : 254 - 0xfe
      13'h9AD: dout  = 8'b11111000; // 2477 : 248 - 0xf8
      13'h9AE: dout  = 8'b11111100; // 2478 : 252 - 0xfc
      13'h9AF: dout  = 8'b11111000; // 2479 : 248 - 0xf8
      13'h9B0: dout  = 8'b00001100; // 2480 :  12 - 0xc -- Sprite 0x9b
      13'h9B1: dout  = 8'b00111000; // 2481 :  56 - 0x38
      13'h9B2: dout  = 8'b11101000; // 2482 : 232 - 0xe8
      13'h9B3: dout  = 8'b11010000; // 2483 : 208 - 0xd0
      13'h9B4: dout  = 8'b11100000; // 2484 : 224 - 0xe0
      13'h9B5: dout  = 8'b10000000; // 2485 : 128 - 0x80
      13'h9B6: dout  = 8'b00000000; // 2486 :   0 - 0x0
      13'h9B7: dout  = 8'b10000000; // 2487 : 128 - 0x80
      13'h9B8: dout  = 8'b11111000; // 2488 : 248 - 0xf8
      13'h9B9: dout  = 8'b11010000; // 2489 : 208 - 0xd0
      13'h9BA: dout  = 8'b00110000; // 2490 :  48 - 0x30
      13'h9BB: dout  = 8'b01100000; // 2491 :  96 - 0x60
      13'h9BC: dout  = 8'b10000000; // 2492 : 128 - 0x80
      13'h9BD: dout  = 8'b00000000; // 2493 :   0 - 0x0
      13'h9BE: dout  = 8'b00000000; // 2494 :   0 - 0x0
      13'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      13'h9C0: dout  = 8'b00000001; // 2496 :   1 - 0x1 -- Sprite 0x9c
      13'h9C1: dout  = 8'b00000000; // 2497 :   0 - 0x0
      13'h9C2: dout  = 8'b00000000; // 2498 :   0 - 0x0
      13'h9C3: dout  = 8'b00000000; // 2499 :   0 - 0x0
      13'h9C4: dout  = 8'b00000001; // 2500 :   1 - 0x1
      13'h9C5: dout  = 8'b00000001; // 2501 :   1 - 0x1
      13'h9C6: dout  = 8'b00000010; // 2502 :   2 - 0x2
      13'h9C7: dout  = 8'b00000110; // 2503 :   6 - 0x6
      13'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0
      13'h9C9: dout  = 8'b00000001; // 2505 :   1 - 0x1
      13'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      13'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      13'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      13'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      13'h9CE: dout  = 8'b00000001; // 2510 :   1 - 0x1
      13'h9CF: dout  = 8'b00000011; // 2511 :   3 - 0x3
      13'h9D0: dout  = 8'b01111000; // 2512 : 120 - 0x78 -- Sprite 0x9d
      13'h9D1: dout  = 8'b00101010; // 2513 :  42 - 0x2a
      13'h9D2: dout  = 8'b01010100; // 2514 :  84 - 0x54
      13'h9D3: dout  = 8'b00101001; // 2515 :  41 - 0x29
      13'h9D4: dout  = 8'b00101111; // 2516 :  47 - 0x2f
      13'h9D5: dout  = 8'b00111100; // 2517 :  60 - 0x3c
      13'h9D6: dout  = 8'b00011110; // 2518 :  30 - 0x1e
      13'h9D7: dout  = 8'b00000000; // 2519 :   0 - 0x0
      13'h9D8: dout  = 8'b00000111; // 2520 :   7 - 0x7
      13'h9D9: dout  = 8'b00010111; // 2521 :  23 - 0x17
      13'h9DA: dout  = 8'b00101111; // 2522 :  47 - 0x2f
      13'h9DB: dout  = 8'b00011110; // 2523 :  30 - 0x1e
      13'h9DC: dout  = 8'b00010000; // 2524 :  16 - 0x10
      13'h9DD: dout  = 8'b00000100; // 2525 :   4 - 0x4
      13'h9DE: dout  = 8'b00000000; // 2526 :   0 - 0x0
      13'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout  = 8'b10110000; // 2528 : 176 - 0xb0 -- Sprite 0x9e
      13'h9E1: dout  = 8'b11101000; // 2529 : 232 - 0xe8
      13'h9E2: dout  = 8'b10001100; // 2530 : 140 - 0x8c
      13'h9E3: dout  = 8'b10011110; // 2531 : 158 - 0x9e
      13'h9E4: dout  = 8'b00011111; // 2532 :  31 - 0x1f
      13'h9E5: dout  = 8'b00001111; // 2533 :  15 - 0xf
      13'h9E6: dout  = 8'b10010110; // 2534 : 150 - 0x96
      13'h9E7: dout  = 8'b00011100; // 2535 :  28 - 0x1c
      13'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout  = 8'b00010000; // 2537 :  16 - 0x10
      13'h9EA: dout  = 8'b01111000; // 2538 : 120 - 0x78
      13'h9EB: dout  = 8'b01110100; // 2539 : 116 - 0x74
      13'h9EC: dout  = 8'b11111110; // 2540 : 254 - 0xfe
      13'h9ED: dout  = 8'b11111000; // 2541 : 248 - 0xf8
      13'h9EE: dout  = 8'b11111100; // 2542 : 252 - 0xfc
      13'h9EF: dout  = 8'b11111000; // 2543 : 248 - 0xf8
      13'h9F0: dout  = 8'b00001100; // 2544 :  12 - 0xc -- Sprite 0x9f
      13'h9F1: dout  = 8'b00111000; // 2545 :  56 - 0x38
      13'h9F2: dout  = 8'b11101000; // 2546 : 232 - 0xe8
      13'h9F3: dout  = 8'b11110000; // 2547 : 240 - 0xf0
      13'h9F4: dout  = 8'b11000000; // 2548 : 192 - 0xc0
      13'h9F5: dout  = 8'b01110000; // 2549 : 112 - 0x70
      13'h9F6: dout  = 8'b11000000; // 2550 : 192 - 0xc0
      13'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      13'h9F8: dout  = 8'b11111000; // 2552 : 248 - 0xf8
      13'h9F9: dout  = 8'b11010000; // 2553 : 208 - 0xd0
      13'h9FA: dout  = 8'b00110000; // 2554 :  48 - 0x30
      13'h9FB: dout  = 8'b11000000; // 2555 : 192 - 0xc0
      13'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      13'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      13'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      13'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout  = 8'b00000011; // 2560 :   3 - 0x3 -- Sprite 0xa0
      13'hA01: dout  = 8'b00001111; // 2561 :  15 - 0xf
      13'hA02: dout  = 8'b00011100; // 2562 :  28 - 0x1c
      13'hA03: dout  = 8'b00110000; // 2563 :  48 - 0x30
      13'hA04: dout  = 8'b01100000; // 2564 :  96 - 0x60
      13'hA05: dout  = 8'b01100000; // 2565 :  96 - 0x60
      13'hA06: dout  = 8'b11000000; // 2566 : 192 - 0xc0
      13'hA07: dout  = 8'b11000000; // 2567 : 192 - 0xc0
      13'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0
      13'hA09: dout  = 8'b00000011; // 2569 :   3 - 0x3
      13'hA0A: dout  = 8'b00001111; // 2570 :  15 - 0xf
      13'hA0B: dout  = 8'b00011111; // 2571 :  31 - 0x1f
      13'hA0C: dout  = 8'b00111111; // 2572 :  63 - 0x3f
      13'hA0D: dout  = 8'b00111111; // 2573 :  63 - 0x3f
      13'hA0E: dout  = 8'b01111111; // 2574 : 127 - 0x7f
      13'hA0F: dout  = 8'b01111111; // 2575 : 127 - 0x7f
      13'hA10: dout  = 8'b11000000; // 2576 : 192 - 0xc0 -- Sprite 0xa1
      13'hA11: dout  = 8'b11000000; // 2577 : 192 - 0xc0
      13'hA12: dout  = 8'b01100000; // 2578 :  96 - 0x60
      13'hA13: dout  = 8'b01100000; // 2579 :  96 - 0x60
      13'hA14: dout  = 8'b00110000; // 2580 :  48 - 0x30
      13'hA15: dout  = 8'b00011010; // 2581 :  26 - 0x1a
      13'hA16: dout  = 8'b00001101; // 2582 :  13 - 0xd
      13'hA17: dout  = 8'b00000011; // 2583 :   3 - 0x3
      13'hA18: dout  = 8'b01111111; // 2584 : 127 - 0x7f
      13'hA19: dout  = 8'b01111111; // 2585 : 127 - 0x7f
      13'hA1A: dout  = 8'b00111111; // 2586 :  63 - 0x3f
      13'hA1B: dout  = 8'b00111111; // 2587 :  63 - 0x3f
      13'hA1C: dout  = 8'b00011111; // 2588 :  31 - 0x1f
      13'hA1D: dout  = 8'b00000101; // 2589 :   5 - 0x5
      13'hA1E: dout  = 8'b00000010; // 2590 :   2 - 0x2
      13'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      13'hA20: dout  = 8'b11000000; // 2592 : 192 - 0xc0 -- Sprite 0xa2
      13'hA21: dout  = 8'b11110000; // 2593 : 240 - 0xf0
      13'hA22: dout  = 8'b00111000; // 2594 :  56 - 0x38
      13'hA23: dout  = 8'b00001100; // 2595 :  12 - 0xc
      13'hA24: dout  = 8'b00000110; // 2596 :   6 - 0x6
      13'hA25: dout  = 8'b00000010; // 2597 :   2 - 0x2
      13'hA26: dout  = 8'b00000101; // 2598 :   5 - 0x5
      13'hA27: dout  = 8'b00000011; // 2599 :   3 - 0x3
      13'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0
      13'hA29: dout  = 8'b11000000; // 2601 : 192 - 0xc0
      13'hA2A: dout  = 8'b11110000; // 2602 : 240 - 0xf0
      13'hA2B: dout  = 8'b11111000; // 2603 : 248 - 0xf8
      13'hA2C: dout  = 8'b11111000; // 2604 : 248 - 0xf8
      13'hA2D: dout  = 8'b11111100; // 2605 : 252 - 0xfc
      13'hA2E: dout  = 8'b11111010; // 2606 : 250 - 0xfa
      13'hA2F: dout  = 8'b11111100; // 2607 : 252 - 0xfc
      13'hA30: dout  = 8'b00000101; // 2608 :   5 - 0x5 -- Sprite 0xa3
      13'hA31: dout  = 8'b00001011; // 2609 :  11 - 0xb
      13'hA32: dout  = 8'b00010110; // 2610 :  22 - 0x16
      13'hA33: dout  = 8'b00101010; // 2611 :  42 - 0x2a
      13'hA34: dout  = 8'b01010100; // 2612 :  84 - 0x54
      13'hA35: dout  = 8'b10101000; // 2613 : 168 - 0xa8
      13'hA36: dout  = 8'b01110000; // 2614 : 112 - 0x70
      13'hA37: dout  = 8'b11000000; // 2615 : 192 - 0xc0
      13'hA38: dout  = 8'b11111010; // 2616 : 250 - 0xfa
      13'hA39: dout  = 8'b11110100; // 2617 : 244 - 0xf4
      13'hA3A: dout  = 8'b11101000; // 2618 : 232 - 0xe8
      13'hA3B: dout  = 8'b11010100; // 2619 : 212 - 0xd4
      13'hA3C: dout  = 8'b10101000; // 2620 : 168 - 0xa8
      13'hA3D: dout  = 8'b01010000; // 2621 :  80 - 0x50
      13'hA3E: dout  = 8'b10000000; // 2622 : 128 - 0x80
      13'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      13'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Sprite 0xa4
      13'hA41: dout  = 8'b00001111; // 2625 :  15 - 0xf
      13'hA42: dout  = 8'b00011111; // 2626 :  31 - 0x1f
      13'hA43: dout  = 8'b00110001; // 2627 :  49 - 0x31
      13'hA44: dout  = 8'b00111111; // 2628 :  63 - 0x3f
      13'hA45: dout  = 8'b01111111; // 2629 : 127 - 0x7f
      13'hA46: dout  = 8'b11111111; // 2630 : 255 - 0xff
      13'hA47: dout  = 8'b11011111; // 2631 : 223 - 0xdf
      13'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0
      13'hA49: dout  = 8'b00000000; // 2633 :   0 - 0x0
      13'hA4A: dout  = 8'b00000000; // 2634 :   0 - 0x0
      13'hA4B: dout  = 8'b00001110; // 2635 :  14 - 0xe
      13'hA4C: dout  = 8'b00000000; // 2636 :   0 - 0x0
      13'hA4D: dout  = 8'b00001010; // 2637 :  10 - 0xa
      13'hA4E: dout  = 8'b01001010; // 2638 :  74 - 0x4a
      13'hA4F: dout  = 8'b01100000; // 2639 :  96 - 0x60
      13'hA50: dout  = 8'b11000000; // 2640 : 192 - 0xc0 -- Sprite 0xa5
      13'hA51: dout  = 8'b11000111; // 2641 : 199 - 0xc7
      13'hA52: dout  = 8'b01101111; // 2642 : 111 - 0x6f
      13'hA53: dout  = 8'b01100111; // 2643 : 103 - 0x67
      13'hA54: dout  = 8'b01100011; // 2644 :  99 - 0x63
      13'hA55: dout  = 8'b00110000; // 2645 :  48 - 0x30
      13'hA56: dout  = 8'b00011000; // 2646 :  24 - 0x18
      13'hA57: dout  = 8'b00000111; // 2647 :   7 - 0x7
      13'hA58: dout  = 8'b01111111; // 2648 : 127 - 0x7f
      13'hA59: dout  = 8'b01111000; // 2649 : 120 - 0x78
      13'hA5A: dout  = 8'b00110111; // 2650 :  55 - 0x37
      13'hA5B: dout  = 8'b00111011; // 2651 :  59 - 0x3b
      13'hA5C: dout  = 8'b00111100; // 2652 :  60 - 0x3c
      13'hA5D: dout  = 8'b00011111; // 2653 :  31 - 0x1f
      13'hA5E: dout  = 8'b00000111; // 2654 :   7 - 0x7
      13'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      13'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Sprite 0xa6
      13'hA61: dout  = 8'b11110000; // 2657 : 240 - 0xf0
      13'hA62: dout  = 8'b11111000; // 2658 : 248 - 0xf8
      13'hA63: dout  = 8'b10001100; // 2659 : 140 - 0x8c
      13'hA64: dout  = 8'b11111100; // 2660 : 252 - 0xfc
      13'hA65: dout  = 8'b11111110; // 2661 : 254 - 0xfe
      13'hA66: dout  = 8'b11111101; // 2662 : 253 - 0xfd
      13'hA67: dout  = 8'b11111001; // 2663 : 249 - 0xf9
      13'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0
      13'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      13'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      13'hA6B: dout  = 8'b01110000; // 2667 : 112 - 0x70
      13'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      13'hA6D: dout  = 8'b01010000; // 2669 :  80 - 0x50
      13'hA6E: dout  = 8'b01010010; // 2670 :  82 - 0x52
      13'hA6F: dout  = 8'b00000110; // 2671 :   6 - 0x6
      13'hA70: dout  = 8'b00000011; // 2672 :   3 - 0x3 -- Sprite 0xa7
      13'hA71: dout  = 8'b11100101; // 2673 : 229 - 0xe5
      13'hA72: dout  = 8'b11110010; // 2674 : 242 - 0xf2
      13'hA73: dout  = 8'b11100110; // 2675 : 230 - 0xe6
      13'hA74: dout  = 8'b11001010; // 2676 : 202 - 0xca
      13'hA75: dout  = 8'b00010100; // 2677 :  20 - 0x14
      13'hA76: dout  = 8'b00111000; // 2678 :  56 - 0x38
      13'hA77: dout  = 8'b11100000; // 2679 : 224 - 0xe0
      13'hA78: dout  = 8'b11111100; // 2680 : 252 - 0xfc
      13'hA79: dout  = 8'b00011010; // 2681 :  26 - 0x1a
      13'hA7A: dout  = 8'b11101100; // 2682 : 236 - 0xec
      13'hA7B: dout  = 8'b11011000; // 2683 : 216 - 0xd8
      13'hA7C: dout  = 8'b00110100; // 2684 :  52 - 0x34
      13'hA7D: dout  = 8'b11101000; // 2685 : 232 - 0xe8
      13'hA7E: dout  = 8'b11000000; // 2686 : 192 - 0xc0
      13'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      13'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      13'hA81: dout  = 8'b00001111; // 2689 :  15 - 0xf
      13'hA82: dout  = 8'b00011111; // 2690 :  31 - 0x1f
      13'hA83: dout  = 8'b00110001; // 2691 :  49 - 0x31
      13'hA84: dout  = 8'b00111111; // 2692 :  63 - 0x3f
      13'hA85: dout  = 8'b01111111; // 2693 : 127 - 0x7f
      13'hA86: dout  = 8'b11111111; // 2694 : 255 - 0xff
      13'hA87: dout  = 8'b11011111; // 2695 : 223 - 0xdf
      13'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0
      13'hA89: dout  = 8'b00000000; // 2697 :   0 - 0x0
      13'hA8A: dout  = 8'b00000000; // 2698 :   0 - 0x0
      13'hA8B: dout  = 8'b00001110; // 2699 :  14 - 0xe
      13'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      13'hA8D: dout  = 8'b00001110; // 2701 :  14 - 0xe
      13'hA8E: dout  = 8'b01001010; // 2702 :  74 - 0x4a
      13'hA8F: dout  = 8'b01100000; // 2703 :  96 - 0x60
      13'hA90: dout  = 8'b11000000; // 2704 : 192 - 0xc0 -- Sprite 0xa9
      13'hA91: dout  = 8'b11000011; // 2705 : 195 - 0xc3
      13'hA92: dout  = 8'b11000111; // 2706 : 199 - 0xc7
      13'hA93: dout  = 8'b11001111; // 2707 : 207 - 0xcf
      13'hA94: dout  = 8'b11000111; // 2708 : 199 - 0xc7
      13'hA95: dout  = 8'b11000000; // 2709 : 192 - 0xc0
      13'hA96: dout  = 8'b11100000; // 2710 : 224 - 0xe0
      13'hA97: dout  = 8'b11111111; // 2711 : 255 - 0xff
      13'hA98: dout  = 8'b01111111; // 2712 : 127 - 0x7f
      13'hA99: dout  = 8'b01111100; // 2713 : 124 - 0x7c
      13'hA9A: dout  = 8'b01111011; // 2714 : 123 - 0x7b
      13'hA9B: dout  = 8'b01110111; // 2715 : 119 - 0x77
      13'hA9C: dout  = 8'b01111000; // 2716 : 120 - 0x78
      13'hA9D: dout  = 8'b01111111; // 2717 : 127 - 0x7f
      13'hA9E: dout  = 8'b01111111; // 2718 : 127 - 0x7f
      13'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Sprite 0xaa
      13'hAA1: dout  = 8'b11110000; // 2721 : 240 - 0xf0
      13'hAA2: dout  = 8'b11111000; // 2722 : 248 - 0xf8
      13'hAA3: dout  = 8'b10001100; // 2723 : 140 - 0x8c
      13'hAA4: dout  = 8'b11111100; // 2724 : 252 - 0xfc
      13'hAA5: dout  = 8'b11111110; // 2725 : 254 - 0xfe
      13'hAA6: dout  = 8'b11111101; // 2726 : 253 - 0xfd
      13'hAA7: dout  = 8'b11111001; // 2727 : 249 - 0xf9
      13'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout  = 8'b01110000; // 2731 : 112 - 0x70
      13'hAAC: dout  = 8'b00000000; // 2732 :   0 - 0x0
      13'hAAD: dout  = 8'b01110000; // 2733 : 112 - 0x70
      13'hAAE: dout  = 8'b01010010; // 2734 :  82 - 0x52
      13'hAAF: dout  = 8'b00000110; // 2735 :   6 - 0x6
      13'hAB0: dout  = 8'b00000011; // 2736 :   3 - 0x3 -- Sprite 0xab
      13'hAB1: dout  = 8'b11000101; // 2737 : 197 - 0xc5
      13'hAB2: dout  = 8'b11100011; // 2738 : 227 - 0xe3
      13'hAB3: dout  = 8'b11110101; // 2739 : 245 - 0xf5
      13'hAB4: dout  = 8'b11100011; // 2740 : 227 - 0xe3
      13'hAB5: dout  = 8'b00000101; // 2741 :   5 - 0x5
      13'hAB6: dout  = 8'b00001011; // 2742 :  11 - 0xb
      13'hAB7: dout  = 8'b11111111; // 2743 : 255 - 0xff
      13'hAB8: dout  = 8'b11111100; // 2744 : 252 - 0xfc
      13'hAB9: dout  = 8'b00111010; // 2745 :  58 - 0x3a
      13'hABA: dout  = 8'b11011100; // 2746 : 220 - 0xdc
      13'hABB: dout  = 8'b11101010; // 2747 : 234 - 0xea
      13'hABC: dout  = 8'b00011100; // 2748 :  28 - 0x1c
      13'hABD: dout  = 8'b11111010; // 2749 : 250 - 0xfa
      13'hABE: dout  = 8'b11110100; // 2750 : 244 - 0xf4
      13'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout  = 8'b10000011; // 2752 : 131 - 0x83 -- Sprite 0xac
      13'hAC1: dout  = 8'b10001100; // 2753 : 140 - 0x8c
      13'hAC2: dout  = 8'b10010000; // 2754 : 144 - 0x90
      13'hAC3: dout  = 8'b10010000; // 2755 : 144 - 0x90
      13'hAC4: dout  = 8'b11100000; // 2756 : 224 - 0xe0
      13'hAC5: dout  = 8'b10100000; // 2757 : 160 - 0xa0
      13'hAC6: dout  = 8'b10101111; // 2758 : 175 - 0xaf
      13'hAC7: dout  = 8'b01101111; // 2759 : 111 - 0x6f
      13'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout  = 8'b00000011; // 2761 :   3 - 0x3
      13'hACA: dout  = 8'b00001111; // 2762 :  15 - 0xf
      13'hACB: dout  = 8'b00001111; // 2763 :  15 - 0xf
      13'hACC: dout  = 8'b00011111; // 2764 :  31 - 0x1f
      13'hACD: dout  = 8'b01011111; // 2765 :  95 - 0x5f
      13'hACE: dout  = 8'b01010000; // 2766 :  80 - 0x50
      13'hACF: dout  = 8'b00010000; // 2767 :  16 - 0x10
      13'hAD0: dout  = 8'b11111011; // 2768 : 251 - 0xfb -- Sprite 0xad
      13'hAD1: dout  = 8'b00000101; // 2769 :   5 - 0x5
      13'hAD2: dout  = 8'b00000101; // 2770 :   5 - 0x5
      13'hAD3: dout  = 8'b00000101; // 2771 :   5 - 0x5
      13'hAD4: dout  = 8'b01000101; // 2772 :  69 - 0x45
      13'hAD5: dout  = 8'b01100101; // 2773 : 101 - 0x65
      13'hAD6: dout  = 8'b11110101; // 2774 : 245 - 0xf5
      13'hAD7: dout  = 8'b11111101; // 2775 : 253 - 0xfd
      13'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0
      13'hAD9: dout  = 8'b11111010; // 2777 : 250 - 0xfa
      13'hADA: dout  = 8'b11111010; // 2778 : 250 - 0xfa
      13'hADB: dout  = 8'b11111010; // 2779 : 250 - 0xfa
      13'hADC: dout  = 8'b10111010; // 2780 : 186 - 0xba
      13'hADD: dout  = 8'b10011010; // 2781 : 154 - 0x9a
      13'hADE: dout  = 8'b00001010; // 2782 :  10 - 0xa
      13'hADF: dout  = 8'b00000010; // 2783 :   2 - 0x2
      13'hAE0: dout  = 8'b10000011; // 2784 : 131 - 0x83 -- Sprite 0xae
      13'hAE1: dout  = 8'b10001100; // 2785 : 140 - 0x8c
      13'hAE2: dout  = 8'b10010000; // 2786 : 144 - 0x90
      13'hAE3: dout  = 8'b10010000; // 2787 : 144 - 0x90
      13'hAE4: dout  = 8'b11100000; // 2788 : 224 - 0xe0
      13'hAE5: dout  = 8'b10100000; // 2789 : 160 - 0xa0
      13'hAE6: dout  = 8'b10101111; // 2790 : 175 - 0xaf
      13'hAE7: dout  = 8'b01101111; // 2791 : 111 - 0x6f
      13'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout  = 8'b00000011; // 2793 :   3 - 0x3
      13'hAEA: dout  = 8'b00001111; // 2794 :  15 - 0xf
      13'hAEB: dout  = 8'b00001111; // 2795 :  15 - 0xf
      13'hAEC: dout  = 8'b00011111; // 2796 :  31 - 0x1f
      13'hAED: dout  = 8'b01011111; // 2797 :  95 - 0x5f
      13'hAEE: dout  = 8'b01010000; // 2798 :  80 - 0x50
      13'hAEF: dout  = 8'b00010111; // 2799 :  23 - 0x17
      13'hAF0: dout  = 8'b11111011; // 2800 : 251 - 0xfb -- Sprite 0xaf
      13'hAF1: dout  = 8'b00000101; // 2801 :   5 - 0x5
      13'hAF2: dout  = 8'b00000101; // 2802 :   5 - 0x5
      13'hAF3: dout  = 8'b00000101; // 2803 :   5 - 0x5
      13'hAF4: dout  = 8'b11000101; // 2804 : 197 - 0xc5
      13'hAF5: dout  = 8'b11100101; // 2805 : 229 - 0xe5
      13'hAF6: dout  = 8'b11110101; // 2806 : 245 - 0xf5
      13'hAF7: dout  = 8'b11111101; // 2807 : 253 - 0xfd
      13'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0
      13'hAF9: dout  = 8'b11111010; // 2809 : 250 - 0xfa
      13'hAFA: dout  = 8'b11111010; // 2810 : 250 - 0xfa
      13'hAFB: dout  = 8'b11111010; // 2811 : 250 - 0xfa
      13'hAFC: dout  = 8'b00111010; // 2812 :  58 - 0x3a
      13'hAFD: dout  = 8'b01011010; // 2813 :  90 - 0x5a
      13'hAFE: dout  = 8'b01101010; // 2814 : 106 - 0x6a
      13'hAFF: dout  = 8'b11110010; // 2815 : 242 - 0xf2
      13'hB00: dout  = 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      13'hB01: dout  = 8'b00000011; // 2817 :   3 - 0x3
      13'hB02: dout  = 8'b00001111; // 2818 :  15 - 0xf
      13'hB03: dout  = 8'b00111111; // 2819 :  63 - 0x3f
      13'hB04: dout  = 8'b01111111; // 2820 : 127 - 0x7f
      13'hB05: dout  = 8'b01111111; // 2821 : 127 - 0x7f
      13'hB06: dout  = 8'b11111111; // 2822 : 255 - 0xff
      13'hB07: dout  = 8'b11111111; // 2823 : 255 - 0xff
      13'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0
      13'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      13'hB0A: dout  = 8'b00000011; // 2826 :   3 - 0x3
      13'hB0B: dout  = 8'b00001111; // 2827 :  15 - 0xf
      13'hB0C: dout  = 8'b00111011; // 2828 :  59 - 0x3b
      13'hB0D: dout  = 8'b00111111; // 2829 :  63 - 0x3f
      13'hB0E: dout  = 8'b01101111; // 2830 : 111 - 0x6f
      13'hB0F: dout  = 8'b01111101; // 2831 : 125 - 0x7d
      13'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Sprite 0xb1
      13'hB11: dout  = 8'b10001111; // 2833 : 143 - 0x8f
      13'hB12: dout  = 8'b10000000; // 2834 : 128 - 0x80
      13'hB13: dout  = 8'b11110000; // 2835 : 240 - 0xf0
      13'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      13'hB15: dout  = 8'b11111111; // 2837 : 255 - 0xff
      13'hB16: dout  = 8'b01111111; // 2838 : 127 - 0x7f
      13'hB17: dout  = 8'b00001111; // 2839 :  15 - 0xf
      13'hB18: dout  = 8'b00001111; // 2840 :  15 - 0xf
      13'hB19: dout  = 8'b01110000; // 2841 : 112 - 0x70
      13'hB1A: dout  = 8'b01111111; // 2842 : 127 - 0x7f
      13'hB1B: dout  = 8'b00001111; // 2843 :  15 - 0xf
      13'hB1C: dout  = 8'b01110000; // 2844 : 112 - 0x70
      13'hB1D: dout  = 8'b01111111; // 2845 : 127 - 0x7f
      13'hB1E: dout  = 8'b00001111; // 2846 :  15 - 0xf
      13'hB1F: dout  = 8'b00000000; // 2847 :   0 - 0x0
      13'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Sprite 0xb2
      13'hB21: dout  = 8'b11000000; // 2849 : 192 - 0xc0
      13'hB22: dout  = 8'b11110000; // 2850 : 240 - 0xf0
      13'hB23: dout  = 8'b11111100; // 2851 : 252 - 0xfc
      13'hB24: dout  = 8'b11111110; // 2852 : 254 - 0xfe
      13'hB25: dout  = 8'b11111110; // 2853 : 254 - 0xfe
      13'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      13'hB27: dout  = 8'b11111111; // 2855 : 255 - 0xff
      13'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0
      13'hB29: dout  = 8'b00000000; // 2857 :   0 - 0x0
      13'hB2A: dout  = 8'b11000000; // 2858 : 192 - 0xc0
      13'hB2B: dout  = 8'b11110000; // 2859 : 240 - 0xf0
      13'hB2C: dout  = 8'b10111100; // 2860 : 188 - 0xbc
      13'hB2D: dout  = 8'b11110100; // 2861 : 244 - 0xf4
      13'hB2E: dout  = 8'b11111110; // 2862 : 254 - 0xfe
      13'hB2F: dout  = 8'b11011110; // 2863 : 222 - 0xde
      13'hB30: dout  = 8'b11111111; // 2864 : 255 - 0xff -- Sprite 0xb3
      13'hB31: dout  = 8'b11110001; // 2865 : 241 - 0xf1
      13'hB32: dout  = 8'b00000001; // 2866 :   1 - 0x1
      13'hB33: dout  = 8'b00001111; // 2867 :  15 - 0xf
      13'hB34: dout  = 8'b11111111; // 2868 : 255 - 0xff
      13'hB35: dout  = 8'b11111111; // 2869 : 255 - 0xff
      13'hB36: dout  = 8'b11111110; // 2870 : 254 - 0xfe
      13'hB37: dout  = 8'b11110000; // 2871 : 240 - 0xf0
      13'hB38: dout  = 8'b11110000; // 2872 : 240 - 0xf0
      13'hB39: dout  = 8'b00001110; // 2873 :  14 - 0xe
      13'hB3A: dout  = 8'b11111110; // 2874 : 254 - 0xfe
      13'hB3B: dout  = 8'b11110000; // 2875 : 240 - 0xf0
      13'hB3C: dout  = 8'b00001110; // 2876 :  14 - 0xe
      13'hB3D: dout  = 8'b11111110; // 2877 : 254 - 0xfe
      13'hB3E: dout  = 8'b11110000; // 2878 : 240 - 0xf0
      13'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Sprite 0xb4
      13'hB41: dout  = 8'b00000011; // 2881 :   3 - 0x3
      13'hB42: dout  = 8'b00001110; // 2882 :  14 - 0xe
      13'hB43: dout  = 8'b00110101; // 2883 :  53 - 0x35
      13'hB44: dout  = 8'b01101110; // 2884 : 110 - 0x6e
      13'hB45: dout  = 8'b01010101; // 2885 :  85 - 0x55
      13'hB46: dout  = 8'b10111010; // 2886 : 186 - 0xba
      13'hB47: dout  = 8'b11010111; // 2887 : 215 - 0xd7
      13'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0
      13'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      13'hB4A: dout  = 8'b00000011; // 2890 :   3 - 0x3
      13'hB4B: dout  = 8'b00001111; // 2891 :  15 - 0xf
      13'hB4C: dout  = 8'b00111011; // 2892 :  59 - 0x3b
      13'hB4D: dout  = 8'b00111111; // 2893 :  63 - 0x3f
      13'hB4E: dout  = 8'b01101111; // 2894 : 111 - 0x6f
      13'hB4F: dout  = 8'b01111101; // 2895 : 125 - 0x7d
      13'hB50: dout  = 8'b11111010; // 2896 : 250 - 0xfa -- Sprite 0xb5
      13'hB51: dout  = 8'b10001111; // 2897 : 143 - 0x8f
      13'hB52: dout  = 8'b10000000; // 2898 : 128 - 0x80
      13'hB53: dout  = 8'b11110000; // 2899 : 240 - 0xf0
      13'hB54: dout  = 8'b10101111; // 2900 : 175 - 0xaf
      13'hB55: dout  = 8'b11010101; // 2901 : 213 - 0xd5
      13'hB56: dout  = 8'b01111010; // 2902 : 122 - 0x7a
      13'hB57: dout  = 8'b00001111; // 2903 :  15 - 0xf
      13'hB58: dout  = 8'b00001111; // 2904 :  15 - 0xf
      13'hB59: dout  = 8'b01110000; // 2905 : 112 - 0x70
      13'hB5A: dout  = 8'b01111111; // 2906 : 127 - 0x7f
      13'hB5B: dout  = 8'b00001111; // 2907 :  15 - 0xf
      13'hB5C: dout  = 8'b01110000; // 2908 : 112 - 0x70
      13'hB5D: dout  = 8'b01111111; // 2909 : 127 - 0x7f
      13'hB5E: dout  = 8'b00001111; // 2910 :  15 - 0xf
      13'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      13'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      13'hB61: dout  = 8'b11000000; // 2913 : 192 - 0xc0
      13'hB62: dout  = 8'b10110000; // 2914 : 176 - 0xb0
      13'hB63: dout  = 8'b01011100; // 2915 :  92 - 0x5c
      13'hB64: dout  = 8'b11101010; // 2916 : 234 - 0xea
      13'hB65: dout  = 8'b01011110; // 2917 :  94 - 0x5e
      13'hB66: dout  = 8'b10101011; // 2918 : 171 - 0xab
      13'hB67: dout  = 8'b01110101; // 2919 : 117 - 0x75
      13'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0
      13'hB69: dout  = 8'b00000000; // 2921 :   0 - 0x0
      13'hB6A: dout  = 8'b11000000; // 2922 : 192 - 0xc0
      13'hB6B: dout  = 8'b11110000; // 2923 : 240 - 0xf0
      13'hB6C: dout  = 8'b10111100; // 2924 : 188 - 0xbc
      13'hB6D: dout  = 8'b11110100; // 2925 : 244 - 0xf4
      13'hB6E: dout  = 8'b11111110; // 2926 : 254 - 0xfe
      13'hB6F: dout  = 8'b11011110; // 2927 : 222 - 0xde
      13'hB70: dout  = 8'b10101111; // 2928 : 175 - 0xaf -- Sprite 0xb7
      13'hB71: dout  = 8'b11110001; // 2929 : 241 - 0xf1
      13'hB72: dout  = 8'b00000001; // 2930 :   1 - 0x1
      13'hB73: dout  = 8'b00001111; // 2931 :  15 - 0xf
      13'hB74: dout  = 8'b11111011; // 2932 : 251 - 0xfb
      13'hB75: dout  = 8'b01010101; // 2933 :  85 - 0x55
      13'hB76: dout  = 8'b10101110; // 2934 : 174 - 0xae
      13'hB77: dout  = 8'b11110000; // 2935 : 240 - 0xf0
      13'hB78: dout  = 8'b11110000; // 2936 : 240 - 0xf0
      13'hB79: dout  = 8'b00001110; // 2937 :  14 - 0xe
      13'hB7A: dout  = 8'b11111110; // 2938 : 254 - 0xfe
      13'hB7B: dout  = 8'b11110000; // 2939 : 240 - 0xf0
      13'hB7C: dout  = 8'b00001110; // 2940 :  14 - 0xe
      13'hB7D: dout  = 8'b11111110; // 2941 : 254 - 0xfe
      13'hB7E: dout  = 8'b11110000; // 2942 : 240 - 0xf0
      13'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Sprite 0xb8
      13'hB81: dout  = 8'b00000011; // 2945 :   3 - 0x3
      13'hB82: dout  = 8'b00001100; // 2946 :  12 - 0xc
      13'hB83: dout  = 8'b00110000; // 2947 :  48 - 0x30
      13'hB84: dout  = 8'b01000100; // 2948 :  68 - 0x44
      13'hB85: dout  = 8'b01000000; // 2949 :  64 - 0x40
      13'hB86: dout  = 8'b10010000; // 2950 : 144 - 0x90
      13'hB87: dout  = 8'b10000010; // 2951 : 130 - 0x82
      13'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0
      13'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      13'hB8A: dout  = 8'b00000011; // 2954 :   3 - 0x3
      13'hB8B: dout  = 8'b00001111; // 2955 :  15 - 0xf
      13'hB8C: dout  = 8'b00111011; // 2956 :  59 - 0x3b
      13'hB8D: dout  = 8'b00111111; // 2957 :  63 - 0x3f
      13'hB8E: dout  = 8'b01101111; // 2958 : 111 - 0x6f
      13'hB8F: dout  = 8'b01111101; // 2959 : 125 - 0x7d
      13'hB90: dout  = 8'b11110000; // 2960 : 240 - 0xf0 -- Sprite 0xb9
      13'hB91: dout  = 8'b11111111; // 2961 : 255 - 0xff
      13'hB92: dout  = 8'b11111111; // 2962 : 255 - 0xff
      13'hB93: dout  = 8'b11111111; // 2963 : 255 - 0xff
      13'hB94: dout  = 8'b10001111; // 2964 : 143 - 0x8f
      13'hB95: dout  = 8'b10000000; // 2965 : 128 - 0x80
      13'hB96: dout  = 8'b01110000; // 2966 : 112 - 0x70
      13'hB97: dout  = 8'b00001111; // 2967 :  15 - 0xf
      13'hB98: dout  = 8'b00001111; // 2968 :  15 - 0xf
      13'hB99: dout  = 8'b00100000; // 2969 :  32 - 0x20
      13'hB9A: dout  = 8'b01010101; // 2970 :  85 - 0x55
      13'hB9B: dout  = 8'b00001010; // 2971 :  10 - 0xa
      13'hB9C: dout  = 8'b01110000; // 2972 : 112 - 0x70
      13'hB9D: dout  = 8'b01111111; // 2973 : 127 - 0x7f
      13'hB9E: dout  = 8'b00001111; // 2974 :  15 - 0xf
      13'hB9F: dout  = 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Sprite 0xba
      13'hBA1: dout  = 8'b11000000; // 2977 : 192 - 0xc0
      13'hBA2: dout  = 8'b00110000; // 2978 :  48 - 0x30
      13'hBA3: dout  = 8'b00001100; // 2979 :  12 - 0xc
      13'hBA4: dout  = 8'b01000010; // 2980 :  66 - 0x42
      13'hBA5: dout  = 8'b00001010; // 2981 :  10 - 0xa
      13'hBA6: dout  = 8'b00000001; // 2982 :   1 - 0x1
      13'hBA7: dout  = 8'b00100001; // 2983 :  33 - 0x21
      13'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0
      13'hBA9: dout  = 8'b00000000; // 2985 :   0 - 0x0
      13'hBAA: dout  = 8'b11000000; // 2986 : 192 - 0xc0
      13'hBAB: dout  = 8'b11110000; // 2987 : 240 - 0xf0
      13'hBAC: dout  = 8'b10111100; // 2988 : 188 - 0xbc
      13'hBAD: dout  = 8'b11110100; // 2989 : 244 - 0xf4
      13'hBAE: dout  = 8'b11111110; // 2990 : 254 - 0xfe
      13'hBAF: dout  = 8'b11011110; // 2991 : 222 - 0xde
      13'hBB0: dout  = 8'b00001111; // 2992 :  15 - 0xf -- Sprite 0xbb
      13'hBB1: dout  = 8'b11111111; // 2993 : 255 - 0xff
      13'hBB2: dout  = 8'b11111111; // 2994 : 255 - 0xff
      13'hBB3: dout  = 8'b11111111; // 2995 : 255 - 0xff
      13'hBB4: dout  = 8'b11110001; // 2996 : 241 - 0xf1
      13'hBB5: dout  = 8'b00000001; // 2997 :   1 - 0x1
      13'hBB6: dout  = 8'b00001110; // 2998 :  14 - 0xe
      13'hBB7: dout  = 8'b11110000; // 2999 : 240 - 0xf0
      13'hBB8: dout  = 8'b11110000; // 3000 : 240 - 0xf0
      13'hBB9: dout  = 8'b00001010; // 3001 :  10 - 0xa
      13'hBBA: dout  = 8'b01010100; // 3002 :  84 - 0x54
      13'hBBB: dout  = 8'b10100000; // 3003 : 160 - 0xa0
      13'hBBC: dout  = 8'b00001110; // 3004 :  14 - 0xe
      13'hBBD: dout  = 8'b11111110; // 3005 : 254 - 0xfe
      13'hBBE: dout  = 8'b11110000; // 3006 : 240 - 0xf0
      13'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout  = 8'b11110011; // 3008 : 243 - 0xf3 -- Sprite 0xbc
      13'hBC1: dout  = 8'b11111111; // 3009 : 255 - 0xff
      13'hBC2: dout  = 8'b11000100; // 3010 : 196 - 0xc4
      13'hBC3: dout  = 8'b11000000; // 3011 : 192 - 0xc0
      13'hBC4: dout  = 8'b01000000; // 3012 :  64 - 0x40
      13'hBC5: dout  = 8'b01100011; // 3013 :  99 - 0x63
      13'hBC6: dout  = 8'b11000111; // 3014 : 199 - 0xc7
      13'hBC7: dout  = 8'b11000110; // 3015 : 198 - 0xc6
      13'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0
      13'hBC9: dout  = 8'b01110011; // 3017 : 115 - 0x73
      13'hBCA: dout  = 8'b01111011; // 3018 : 123 - 0x7b
      13'hBCB: dout  = 8'b01111111; // 3019 : 127 - 0x7f
      13'hBCC: dout  = 8'b00111111; // 3020 :  63 - 0x3f
      13'hBCD: dout  = 8'b00011100; // 3021 :  28 - 0x1c
      13'hBCE: dout  = 8'b01111011; // 3022 : 123 - 0x7b
      13'hBCF: dout  = 8'b01111011; // 3023 : 123 - 0x7b
      13'hBD0: dout  = 8'b11000110; // 3024 : 198 - 0xc6 -- Sprite 0xbd
      13'hBD1: dout  = 8'b11000110; // 3025 : 198 - 0xc6
      13'hBD2: dout  = 8'b01100011; // 3026 :  99 - 0x63
      13'hBD3: dout  = 8'b01000000; // 3027 :  64 - 0x40
      13'hBD4: dout  = 8'b11000000; // 3028 : 192 - 0xc0
      13'hBD5: dout  = 8'b11000100; // 3029 : 196 - 0xc4
      13'hBD6: dout  = 8'b11001100; // 3030 : 204 - 0xcc
      13'hBD7: dout  = 8'b11110011; // 3031 : 243 - 0xf3
      13'hBD8: dout  = 8'b01111011; // 3032 : 123 - 0x7b
      13'hBD9: dout  = 8'b01111011; // 3033 : 123 - 0x7b
      13'hBDA: dout  = 8'b00011100; // 3034 :  28 - 0x1c
      13'hBDB: dout  = 8'b00111111; // 3035 :  63 - 0x3f
      13'hBDC: dout  = 8'b01111111; // 3036 : 127 - 0x7f
      13'hBDD: dout  = 8'b01111011; // 3037 : 123 - 0x7b
      13'hBDE: dout  = 8'b01110011; // 3038 : 115 - 0x73
      13'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout  = 8'b11001111; // 3040 : 207 - 0xcf -- Sprite 0xbe
      13'hBE1: dout  = 8'b11111111; // 3041 : 255 - 0xff
      13'hBE2: dout  = 8'b00100001; // 3042 :  33 - 0x21
      13'hBE3: dout  = 8'b00000001; // 3043 :   1 - 0x1
      13'hBE4: dout  = 8'b00000010; // 3044 :   2 - 0x2
      13'hBE5: dout  = 8'b11000110; // 3045 : 198 - 0xc6
      13'hBE6: dout  = 8'b11100001; // 3046 : 225 - 0xe1
      13'hBE7: dout  = 8'b00100001; // 3047 :  33 - 0x21
      13'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout  = 8'b11001110; // 3049 : 206 - 0xce
      13'hBEA: dout  = 8'b11011110; // 3050 : 222 - 0xde
      13'hBEB: dout  = 8'b11111110; // 3051 : 254 - 0xfe
      13'hBEC: dout  = 8'b11111100; // 3052 : 252 - 0xfc
      13'hBED: dout  = 8'b00111000; // 3053 :  56 - 0x38
      13'hBEE: dout  = 8'b11011110; // 3054 : 222 - 0xde
      13'hBEF: dout  = 8'b11011110; // 3055 : 222 - 0xde
      13'hBF0: dout  = 8'b00100001; // 3056 :  33 - 0x21 -- Sprite 0xbf
      13'hBF1: dout  = 8'b00100001; // 3057 :  33 - 0x21
      13'hBF2: dout  = 8'b11000110; // 3058 : 198 - 0xc6
      13'hBF3: dout  = 8'b00000010; // 3059 :   2 - 0x2
      13'hBF4: dout  = 8'b00000001; // 3060 :   1 - 0x1
      13'hBF5: dout  = 8'b00100001; // 3061 :  33 - 0x21
      13'hBF6: dout  = 8'b00110001; // 3062 :  49 - 0x31
      13'hBF7: dout  = 8'b11001111; // 3063 : 207 - 0xcf
      13'hBF8: dout  = 8'b11011110; // 3064 : 222 - 0xde
      13'hBF9: dout  = 8'b11011110; // 3065 : 222 - 0xde
      13'hBFA: dout  = 8'b00111000; // 3066 :  56 - 0x38
      13'hBFB: dout  = 8'b11111100; // 3067 : 252 - 0xfc
      13'hBFC: dout  = 8'b11111110; // 3068 : 254 - 0xfe
      13'hBFD: dout  = 8'b11011110; // 3069 : 222 - 0xde
      13'hBFE: dout  = 8'b11001110; // 3070 : 206 - 0xce
      13'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      13'hC01: dout  = 8'b01010000; // 3073 :  80 - 0x50
      13'hC02: dout  = 8'b10110011; // 3074 : 179 - 0xb3
      13'hC03: dout  = 8'b10010111; // 3075 : 151 - 0x97
      13'hC04: dout  = 8'b10011111; // 3076 : 159 - 0x9f
      13'hC05: dout  = 8'b01101111; // 3077 : 111 - 0x6f
      13'hC06: dout  = 8'b00011111; // 3078 :  31 - 0x1f
      13'hC07: dout  = 8'b00011111; // 3079 :  31 - 0x1f
      13'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout  = 8'b01000000; // 3082 :  64 - 0x40
      13'hC0B: dout  = 8'b01100000; // 3083 :  96 - 0x60
      13'hC0C: dout  = 8'b01100001; // 3084 :  97 - 0x61
      13'hC0D: dout  = 8'b00000010; // 3085 :   2 - 0x2
      13'hC0E: dout  = 8'b00000010; // 3086 :   2 - 0x2
      13'hC0F: dout  = 8'b00000111; // 3087 :   7 - 0x7
      13'hC10: dout  = 8'b00011111; // 3088 :  31 - 0x1f -- Sprite 0xc1
      13'hC11: dout  = 8'b00011111; // 3089 :  31 - 0x1f
      13'hC12: dout  = 8'b00001111; // 3090 :  15 - 0xf
      13'hC13: dout  = 8'b00000111; // 3091 :   7 - 0x7
      13'hC14: dout  = 8'b00011101; // 3092 :  29 - 0x1d
      13'hC15: dout  = 8'b00101100; // 3093 :  44 - 0x2c
      13'hC16: dout  = 8'b01010100; // 3094 :  84 - 0x54
      13'hC17: dout  = 8'b01111100; // 3095 : 124 - 0x7c
      13'hC18: dout  = 8'b00000111; // 3096 :   7 - 0x7
      13'hC19: dout  = 8'b00000100; // 3097 :   4 - 0x4
      13'hC1A: dout  = 8'b00000111; // 3098 :   7 - 0x7
      13'hC1B: dout  = 8'b00000001; // 3099 :   1 - 0x1
      13'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      13'hC1D: dout  = 8'b00010000; // 3101 :  16 - 0x10
      13'hC1E: dout  = 8'b00101000; // 3102 :  40 - 0x28
      13'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      13'hC21: dout  = 8'b00001010; // 3105 :  10 - 0xa
      13'hC22: dout  = 8'b11001101; // 3106 : 205 - 0xcd
      13'hC23: dout  = 8'b11101001; // 3107 : 233 - 0xe9
      13'hC24: dout  = 8'b11111001; // 3108 : 249 - 0xf9
      13'hC25: dout  = 8'b11110110; // 3109 : 246 - 0xf6
      13'hC26: dout  = 8'b11110000; // 3110 : 240 - 0xf0
      13'hC27: dout  = 8'b11111000; // 3111 : 248 - 0xf8
      13'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout  = 8'b00000010; // 3114 :   2 - 0x2
      13'hC2B: dout  = 8'b00000110; // 3115 :   6 - 0x6
      13'hC2C: dout  = 8'b11100110; // 3116 : 230 - 0xe6
      13'hC2D: dout  = 8'b10100000; // 3117 : 160 - 0xa0
      13'hC2E: dout  = 8'b10100000; // 3118 : 160 - 0xa0
      13'hC2F: dout  = 8'b11110000; // 3119 : 240 - 0xf0
      13'hC30: dout  = 8'b11111000; // 3120 : 248 - 0xf8 -- Sprite 0xc3
      13'hC31: dout  = 8'b11111000; // 3121 : 248 - 0xf8
      13'hC32: dout  = 8'b11110000; // 3122 : 240 - 0xf0
      13'hC33: dout  = 8'b11000000; // 3123 : 192 - 0xc0
      13'hC34: dout  = 8'b10111000; // 3124 : 184 - 0xb8
      13'hC35: dout  = 8'b00110100; // 3125 :  52 - 0x34
      13'hC36: dout  = 8'b00101010; // 3126 :  42 - 0x2a
      13'hC37: dout  = 8'b00111110; // 3127 :  62 - 0x3e
      13'hC38: dout  = 8'b11110000; // 3128 : 240 - 0xf0
      13'hC39: dout  = 8'b00110000; // 3129 :  48 - 0x30
      13'hC3A: dout  = 8'b11000000; // 3130 : 192 - 0xc0
      13'hC3B: dout  = 8'b10000000; // 3131 : 128 - 0x80
      13'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      13'hC3D: dout  = 8'b00001000; // 3133 :   8 - 0x8
      13'hC3E: dout  = 8'b00010100; // 3134 :  20 - 0x14
      13'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout  = 8'b00000101; // 3136 :   5 - 0x5 -- Sprite 0xc4
      13'hC41: dout  = 8'b00001010; // 3137 :  10 - 0xa
      13'hC42: dout  = 8'b00001000; // 3138 :   8 - 0x8
      13'hC43: dout  = 8'b00001111; // 3139 :  15 - 0xf
      13'hC44: dout  = 8'b00000001; // 3140 :   1 - 0x1
      13'hC45: dout  = 8'b00000011; // 3141 :   3 - 0x3
      13'hC46: dout  = 8'b00000111; // 3142 :   7 - 0x7
      13'hC47: dout  = 8'b00001111; // 3143 :  15 - 0xf
      13'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout  = 8'b00000101; // 3145 :   5 - 0x5
      13'hC4A: dout  = 8'b00000111; // 3146 :   7 - 0x7
      13'hC4B: dout  = 8'b00000000; // 3147 :   0 - 0x0
      13'hC4C: dout  = 8'b00000000; // 3148 :   0 - 0x0
      13'hC4D: dout  = 8'b00000000; // 3149 :   0 - 0x0
      13'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout  = 8'b00000001; // 3151 :   1 - 0x1
      13'hC50: dout  = 8'b00001111; // 3152 :  15 - 0xf -- Sprite 0xc5
      13'hC51: dout  = 8'b11101111; // 3153 : 239 - 0xef
      13'hC52: dout  = 8'b11011111; // 3154 : 223 - 0xdf
      13'hC53: dout  = 8'b10101111; // 3155 : 175 - 0xaf
      13'hC54: dout  = 8'b01100111; // 3156 : 103 - 0x67
      13'hC55: dout  = 8'b00001101; // 3157 :  13 - 0xd
      13'hC56: dout  = 8'b00001010; // 3158 :  10 - 0xa
      13'hC57: dout  = 8'b00000111; // 3159 :   7 - 0x7
      13'hC58: dout  = 8'b00000010; // 3160 :   2 - 0x2
      13'hC59: dout  = 8'b00000111; // 3161 :   7 - 0x7
      13'hC5A: dout  = 8'b00100111; // 3162 :  39 - 0x27
      13'hC5B: dout  = 8'b01010011; // 3163 :  83 - 0x53
      13'hC5C: dout  = 8'b00000000; // 3164 :   0 - 0x0
      13'hC5D: dout  = 8'b00000010; // 3165 :   2 - 0x2
      13'hC5E: dout  = 8'b00000101; // 3166 :   5 - 0x5
      13'hC5F: dout  = 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Sprite 0xc6
      13'hC61: dout  = 8'b10000000; // 3169 : 128 - 0x80
      13'hC62: dout  = 8'b10000000; // 3170 : 128 - 0x80
      13'hC63: dout  = 8'b11110000; // 3171 : 240 - 0xf0
      13'hC64: dout  = 8'b11111000; // 3172 : 248 - 0xf8
      13'hC65: dout  = 8'b11111100; // 3173 : 252 - 0xfc
      13'hC66: dout  = 8'b11111100; // 3174 : 252 - 0xfc
      13'hC67: dout  = 8'b11111100; // 3175 : 252 - 0xfc
      13'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0
      13'hC69: dout  = 8'b00000000; // 3177 :   0 - 0x0
      13'hC6A: dout  = 8'b00000000; // 3178 :   0 - 0x0
      13'hC6B: dout  = 8'b00000000; // 3179 :   0 - 0x0
      13'hC6C: dout  = 8'b00000000; // 3180 :   0 - 0x0
      13'hC6D: dout  = 8'b01100000; // 3181 :  96 - 0x60
      13'hC6E: dout  = 8'b11011000; // 3182 : 216 - 0xd8
      13'hC6F: dout  = 8'b10110000; // 3183 : 176 - 0xb0
      13'hC70: dout  = 8'b11111100; // 3184 : 252 - 0xfc -- Sprite 0xc7
      13'hC71: dout  = 8'b11111110; // 3185 : 254 - 0xfe
      13'hC72: dout  = 8'b11111001; // 3186 : 249 - 0xf9
      13'hC73: dout  = 8'b11111010; // 3187 : 250 - 0xfa
      13'hC74: dout  = 8'b11101001; // 3188 : 233 - 0xe9
      13'hC75: dout  = 8'b00001110; // 3189 :  14 - 0xe
      13'hC76: dout  = 8'b10000000; // 3190 : 128 - 0x80
      13'hC77: dout  = 8'b00000000; // 3191 :   0 - 0x0
      13'hC78: dout  = 8'b11101000; // 3192 : 232 - 0xe8
      13'hC79: dout  = 8'b01111000; // 3193 : 120 - 0x78
      13'hC7A: dout  = 8'b10110110; // 3194 : 182 - 0xb6
      13'hC7B: dout  = 8'b11100100; // 3195 : 228 - 0xe4
      13'hC7C: dout  = 8'b00000110; // 3196 :   6 - 0x6
      13'hC7D: dout  = 8'b00000000; // 3197 :   0 - 0x0
      13'hC7E: dout  = 8'b00000000; // 3198 :   0 - 0x0
      13'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      13'hC81: dout  = 8'b11000000; // 3201 : 192 - 0xc0
      13'hC82: dout  = 8'b10100000; // 3202 : 160 - 0xa0
      13'hC83: dout  = 8'b11010011; // 3203 : 211 - 0xd3
      13'hC84: dout  = 8'b10110111; // 3204 : 183 - 0xb7
      13'hC85: dout  = 8'b11111111; // 3205 : 255 - 0xff
      13'hC86: dout  = 8'b00001111; // 3206 :  15 - 0xf
      13'hC87: dout  = 8'b00011111; // 3207 :  31 - 0x1f
      13'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      13'hC8A: dout  = 8'b01000000; // 3210 :  64 - 0x40
      13'hC8B: dout  = 8'b00100000; // 3211 :  32 - 0x20
      13'hC8C: dout  = 8'b01000000; // 3212 :  64 - 0x40
      13'hC8D: dout  = 8'b00000111; // 3213 :   7 - 0x7
      13'hC8E: dout  = 8'b00000101; // 3214 :   5 - 0x5
      13'hC8F: dout  = 8'b00001101; // 3215 :  13 - 0xd
      13'hC90: dout  = 8'b00011111; // 3216 :  31 - 0x1f -- Sprite 0xc9
      13'hC91: dout  = 8'b00001111; // 3217 :  15 - 0xf
      13'hC92: dout  = 8'b11110111; // 3218 : 247 - 0xf7
      13'hC93: dout  = 8'b10110111; // 3219 : 183 - 0xb7
      13'hC94: dout  = 8'b11010011; // 3220 : 211 - 0xd3
      13'hC95: dout  = 8'b10100000; // 3221 : 160 - 0xa0
      13'hC96: dout  = 8'b11000000; // 3222 : 192 - 0xc0
      13'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout  = 8'b00001101; // 3224 :  13 - 0xd
      13'hC99: dout  = 8'b00000101; // 3225 :   5 - 0x5
      13'hC9A: dout  = 8'b00000011; // 3226 :   3 - 0x3
      13'hC9B: dout  = 8'b01000011; // 3227 :  67 - 0x43
      13'hC9C: dout  = 8'b00100000; // 3228 :  32 - 0x20
      13'hC9D: dout  = 8'b01000000; // 3229 :  64 - 0x40
      13'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout  = 8'b00011100; // 3232 :  28 - 0x1c -- Sprite 0xca
      13'hCA1: dout  = 8'b00100010; // 3233 :  34 - 0x22
      13'hCA2: dout  = 8'b00100100; // 3234 :  36 - 0x24
      13'hCA3: dout  = 8'b11011110; // 3235 : 222 - 0xde
      13'hCA4: dout  = 8'b11110000; // 3236 : 240 - 0xf0
      13'hCA5: dout  = 8'b11111000; // 3237 : 248 - 0xf8
      13'hCA6: dout  = 8'b11111100; // 3238 : 252 - 0xfc
      13'hCA7: dout  = 8'b11111100; // 3239 : 252 - 0xfc
      13'hCA8: dout  = 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout  = 8'b00011100; // 3241 :  28 - 0x1c
      13'hCAA: dout  = 8'b00011000; // 3242 :  24 - 0x18
      13'hCAB: dout  = 8'b00000000; // 3243 :   0 - 0x0
      13'hCAC: dout  = 8'b00000000; // 3244 :   0 - 0x0
      13'hCAD: dout  = 8'b10000000; // 3245 : 128 - 0x80
      13'hCAE: dout  = 8'b11100000; // 3246 : 224 - 0xe0
      13'hCAF: dout  = 8'b10010000; // 3247 : 144 - 0x90
      13'hCB0: dout  = 8'b11111100; // 3248 : 252 - 0xfc -- Sprite 0xcb
      13'hCB1: dout  = 8'b11111100; // 3249 : 252 - 0xfc
      13'hCB2: dout  = 8'b11111000; // 3250 : 248 - 0xf8
      13'hCB3: dout  = 8'b11110000; // 3251 : 240 - 0xf0
      13'hCB4: dout  = 8'b10011110; // 3252 : 158 - 0x9e
      13'hCB5: dout  = 8'b00100100; // 3253 :  36 - 0x24
      13'hCB6: dout  = 8'b00100010; // 3254 :  34 - 0x22
      13'hCB7: dout  = 8'b00011100; // 3255 :  28 - 0x1c
      13'hCB8: dout  = 8'b11110000; // 3256 : 240 - 0xf0
      13'hCB9: dout  = 8'b10010000; // 3257 : 144 - 0x90
      13'hCBA: dout  = 8'b11110000; // 3258 : 240 - 0xf0
      13'hCBB: dout  = 8'b10000000; // 3259 : 128 - 0x80
      13'hCBC: dout  = 8'b00000000; // 3260 :   0 - 0x0
      13'hCBD: dout  = 8'b00011000; // 3261 :  24 - 0x18
      13'hCBE: dout  = 8'b00011100; // 3262 :  28 - 0x1c
      13'hCBF: dout  = 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout  = 8'b00001110; // 3264 :  14 - 0xe -- Sprite 0xcc
      13'hCC1: dout  = 8'b00010110; // 3265 :  22 - 0x16
      13'hCC2: dout  = 8'b00011010; // 3266 :  26 - 0x1a
      13'hCC3: dout  = 8'b00000100; // 3267 :   4 - 0x4
      13'hCC4: dout  = 8'b01101111; // 3268 : 111 - 0x6f
      13'hCC5: dout  = 8'b10111111; // 3269 : 191 - 0xbf
      13'hCC6: dout  = 8'b11011111; // 3270 : 223 - 0xdf
      13'hCC7: dout  = 8'b10111111; // 3271 : 191 - 0xbf
      13'hCC8: dout  = 8'b00000000; // 3272 :   0 - 0x0
      13'hCC9: dout  = 8'b00001000; // 3273 :   8 - 0x8
      13'hCCA: dout  = 8'b00000100; // 3274 :   4 - 0x4
      13'hCCB: dout  = 8'b00001000; // 3275 :   8 - 0x8
      13'hCCC: dout  = 8'b00000000; // 3276 :   0 - 0x0
      13'hCCD: dout  = 8'b01000110; // 3277 :  70 - 0x46
      13'hCCE: dout  = 8'b00101111; // 3278 :  47 - 0x2f
      13'hCCF: dout  = 8'b01001110; // 3279 :  78 - 0x4e
      13'hCD0: dout  = 8'b01011111; // 3280 :  95 - 0x5f -- Sprite 0xcd
      13'hCD1: dout  = 8'b00011111; // 3281 :  31 - 0x1f
      13'hCD2: dout  = 8'b00011111; // 3282 :  31 - 0x1f
      13'hCD3: dout  = 8'b00001111; // 3283 :  15 - 0xf
      13'hCD4: dout  = 8'b00111111; // 3284 :  63 - 0x3f
      13'hCD5: dout  = 8'b00100011; // 3285 :  35 - 0x23
      13'hCD6: dout  = 8'b00101010; // 3286 :  42 - 0x2a
      13'hCD7: dout  = 8'b00010100; // 3287 :  20 - 0x14
      13'hCD8: dout  = 8'b00001101; // 3288 :  13 - 0xd
      13'hCD9: dout  = 8'b00001011; // 3289 :  11 - 0xb
      13'hCDA: dout  = 8'b00001111; // 3290 :  15 - 0xf
      13'hCDB: dout  = 8'b00000110; // 3291 :   6 - 0x6
      13'hCDC: dout  = 8'b00000011; // 3292 :   3 - 0x3
      13'hCDD: dout  = 8'b00011100; // 3293 :  28 - 0x1c
      13'hCDE: dout  = 8'b00010100; // 3294 :  20 - 0x14
      13'hCDF: dout  = 8'b00000000; // 3295 :   0 - 0x0
      13'hCE0: dout  = 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      13'hCE1: dout  = 8'b00000000; // 3297 :   0 - 0x0
      13'hCE2: dout  = 8'b00000000; // 3298 :   0 - 0x0
      13'hCE3: dout  = 8'b00000000; // 3299 :   0 - 0x0
      13'hCE4: dout  = 8'b10001110; // 3300 : 142 - 0x8e
      13'hCE5: dout  = 8'b11001001; // 3301 : 201 - 0xc9
      13'hCE6: dout  = 8'b11101010; // 3302 : 234 - 0xea
      13'hCE7: dout  = 8'b11111001; // 3303 : 249 - 0xf9
      13'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout  = 8'b00000000; // 3305 :   0 - 0x0
      13'hCEA: dout  = 8'b00000000; // 3306 :   0 - 0x0
      13'hCEB: dout  = 8'b00000000; // 3307 :   0 - 0x0
      13'hCEC: dout  = 8'b00000000; // 3308 :   0 - 0x0
      13'hCED: dout  = 8'b00000110; // 3309 :   6 - 0x6
      13'hCEE: dout  = 8'b00000100; // 3310 :   4 - 0x4
      13'hCEF: dout  = 8'b10000110; // 3311 : 134 - 0x86
      13'hCF0: dout  = 8'b11111110; // 3312 : 254 - 0xfe -- Sprite 0xcf
      13'hCF1: dout  = 8'b11111000; // 3313 : 248 - 0xf8
      13'hCF2: dout  = 8'b11111000; // 3314 : 248 - 0xf8
      13'hCF3: dout  = 8'b11111000; // 3315 : 248 - 0xf8
      13'hCF4: dout  = 8'b11110000; // 3316 : 240 - 0xf0
      13'hCF5: dout  = 8'b11100000; // 3317 : 224 - 0xe0
      13'hCF6: dout  = 8'b00000000; // 3318 :   0 - 0x0
      13'hCF7: dout  = 8'b00000000; // 3319 :   0 - 0x0
      13'hCF8: dout  = 8'b11000000; // 3320 : 192 - 0xc0
      13'hCF9: dout  = 8'b01100000; // 3321 :  96 - 0x60
      13'hCFA: dout  = 8'b10100000; // 3322 : 160 - 0xa0
      13'hCFB: dout  = 8'b11000000; // 3323 : 192 - 0xc0
      13'hCFC: dout  = 8'b01000000; // 3324 :  64 - 0x40
      13'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      13'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      13'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      13'hD00: dout  = 8'b00000000; // 3328 :   0 - 0x0 -- Sprite 0xd0
      13'hD01: dout  = 8'b00000000; // 3329 :   0 - 0x0
      13'hD02: dout  = 8'b00000100; // 3330 :   4 - 0x4
      13'hD03: dout  = 8'b00100110; // 3331 :  38 - 0x26
      13'hD04: dout  = 8'b00101011; // 3332 :  43 - 0x2b
      13'hD05: dout  = 8'b01110001; // 3333 : 113 - 0x71
      13'hD06: dout  = 8'b01000000; // 3334 :  64 - 0x40
      13'hD07: dout  = 8'b01000111; // 3335 :  71 - 0x47
      13'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout  = 8'b00000000; // 3338 :   0 - 0x0
      13'hD0B: dout  = 8'b00000000; // 3339 :   0 - 0x0
      13'hD0C: dout  = 8'b00000100; // 3340 :   4 - 0x4
      13'hD0D: dout  = 8'b00001110; // 3341 :  14 - 0xe
      13'hD0E: dout  = 8'b00111111; // 3342 :  63 - 0x3f
      13'hD0F: dout  = 8'b00111001; // 3343 :  57 - 0x39
      13'hD10: dout  = 8'b10001111; // 3344 : 143 - 0x8f -- Sprite 0xd1
      13'hD11: dout  = 8'b10001111; // 3345 : 143 - 0x8f
      13'hD12: dout  = 8'b01001111; // 3346 :  79 - 0x4f
      13'hD13: dout  = 8'b01001111; // 3347 :  79 - 0x4f
      13'hD14: dout  = 8'b00111111; // 3348 :  63 - 0x3f
      13'hD15: dout  = 8'b00010011; // 3349 :  19 - 0x13
      13'hD16: dout  = 8'b00010001; // 3350 :  17 - 0x11
      13'hD17: dout  = 8'b00011111; // 3351 :  31 - 0x1f
      13'hD18: dout  = 8'b01110000; // 3352 : 112 - 0x70
      13'hD19: dout  = 8'b01111000; // 3353 : 120 - 0x78
      13'hD1A: dout  = 8'b00111111; // 3354 :  63 - 0x3f
      13'hD1B: dout  = 8'b00111111; // 3355 :  63 - 0x3f
      13'hD1C: dout  = 8'b00000011; // 3356 :   3 - 0x3
      13'hD1D: dout  = 8'b00001100; // 3357 :  12 - 0xc
      13'hD1E: dout  = 8'b00001110; // 3358 :  14 - 0xe
      13'hD1F: dout  = 8'b00000000; // 3359 :   0 - 0x0
      13'hD20: dout  = 8'b00000000; // 3360 :   0 - 0x0 -- Sprite 0xd2
      13'hD21: dout  = 8'b10000000; // 3361 : 128 - 0x80
      13'hD22: dout  = 8'b11001000; // 3362 : 200 - 0xc8
      13'hD23: dout  = 8'b11010100; // 3363 : 212 - 0xd4
      13'hD24: dout  = 8'b00100100; // 3364 :  36 - 0x24
      13'hD25: dout  = 8'b00000010; // 3365 :   2 - 0x2
      13'hD26: dout  = 8'b00000010; // 3366 :   2 - 0x2
      13'hD27: dout  = 8'b11110010; // 3367 : 242 - 0xf2
      13'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0
      13'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      13'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      13'hD2B: dout  = 8'b00001000; // 3371 :   8 - 0x8
      13'hD2C: dout  = 8'b11011000; // 3372 : 216 - 0xd8
      13'hD2D: dout  = 8'b11111100; // 3373 : 252 - 0xfc
      13'hD2E: dout  = 8'b11111100; // 3374 : 252 - 0xfc
      13'hD2F: dout  = 8'b10011100; // 3375 : 156 - 0x9c
      13'hD30: dout  = 8'b11110010; // 3376 : 242 - 0xf2 -- Sprite 0xd3
      13'hD31: dout  = 8'b11110010; // 3377 : 242 - 0xf2
      13'hD32: dout  = 8'b11110100; // 3378 : 244 - 0xf4
      13'hD33: dout  = 8'b11110100; // 3379 : 244 - 0xf4
      13'hD34: dout  = 8'b11110100; // 3380 : 244 - 0xf4
      13'hD35: dout  = 8'b11001000; // 3381 : 200 - 0xc8
      13'hD36: dout  = 8'b01000100; // 3382 :  68 - 0x44
      13'hD37: dout  = 8'b01111100; // 3383 : 124 - 0x7c
      13'hD38: dout  = 8'b00001100; // 3384 :  12 - 0xc
      13'hD39: dout  = 8'b10011100; // 3385 : 156 - 0x9c
      13'hD3A: dout  = 8'b11111000; // 3386 : 248 - 0xf8
      13'hD3B: dout  = 8'b01111000; // 3387 : 120 - 0x78
      13'hD3C: dout  = 8'b10001000; // 3388 : 136 - 0x88
      13'hD3D: dout  = 8'b00110000; // 3389 :  48 - 0x30
      13'hD3E: dout  = 8'b00111000; // 3390 :  56 - 0x38
      13'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      13'hD40: dout  = 8'b00000000; // 3392 :   0 - 0x0 -- Sprite 0xd4
      13'hD41: dout  = 8'b00000000; // 3393 :   0 - 0x0
      13'hD42: dout  = 8'b00000000; // 3394 :   0 - 0x0
      13'hD43: dout  = 8'b00001001; // 3395 :   9 - 0x9
      13'hD44: dout  = 8'b00011010; // 3396 :  26 - 0x1a
      13'hD45: dout  = 8'b00010100; // 3397 :  20 - 0x14
      13'hD46: dout  = 8'b00100000; // 3398 :  32 - 0x20
      13'hD47: dout  = 8'b01000111; // 3399 :  71 - 0x47
      13'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout  = 8'b00000000; // 3401 :   0 - 0x0
      13'hD4A: dout  = 8'b00000000; // 3402 :   0 - 0x0
      13'hD4B: dout  = 8'b00000000; // 3403 :   0 - 0x0
      13'hD4C: dout  = 8'b00000001; // 3404 :   1 - 0x1
      13'hD4D: dout  = 8'b00001011; // 3405 :  11 - 0xb
      13'hD4E: dout  = 8'b00011111; // 3406 :  31 - 0x1f
      13'hD4F: dout  = 8'b00111001; // 3407 :  57 - 0x39
      13'hD50: dout  = 8'b10001111; // 3408 : 143 - 0x8f -- Sprite 0xd5
      13'hD51: dout  = 8'b10001111; // 3409 : 143 - 0x8f
      13'hD52: dout  = 8'b01001111; // 3410 :  79 - 0x4f
      13'hD53: dout  = 8'b01001111; // 3411 :  79 - 0x4f
      13'hD54: dout  = 8'b00111111; // 3412 :  63 - 0x3f
      13'hD55: dout  = 8'b01000111; // 3413 :  71 - 0x47
      13'hD56: dout  = 8'b00100010; // 3414 :  34 - 0x22
      13'hD57: dout  = 8'b00011100; // 3415 :  28 - 0x1c
      13'hD58: dout  = 8'b01110000; // 3416 : 112 - 0x70
      13'hD59: dout  = 8'b01111000; // 3417 : 120 - 0x78
      13'hD5A: dout  = 8'b00111111; // 3418 :  63 - 0x3f
      13'hD5B: dout  = 8'b00111111; // 3419 :  63 - 0x3f
      13'hD5C: dout  = 8'b00000011; // 3420 :   3 - 0x3
      13'hD5D: dout  = 8'b00111000; // 3421 :  56 - 0x38
      13'hD5E: dout  = 8'b00011100; // 3422 :  28 - 0x1c
      13'hD5F: dout  = 8'b00000000; // 3423 :   0 - 0x0
      13'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      13'hD61: dout  = 8'b01000000; // 3425 :  64 - 0x40
      13'hD62: dout  = 8'b11000000; // 3426 : 192 - 0xc0
      13'hD63: dout  = 8'b00101100; // 3427 :  44 - 0x2c
      13'hD64: dout  = 8'b00110100; // 3428 :  52 - 0x34
      13'hD65: dout  = 8'b00000100; // 3429 :   4 - 0x4
      13'hD66: dout  = 8'b00000010; // 3430 :   2 - 0x2
      13'hD67: dout  = 8'b11110010; // 3431 : 242 - 0xf2
      13'hD68: dout  = 8'b00000000; // 3432 :   0 - 0x0
      13'hD69: dout  = 8'b00000000; // 3433 :   0 - 0x0
      13'hD6A: dout  = 8'b00000000; // 3434 :   0 - 0x0
      13'hD6B: dout  = 8'b11000000; // 3435 : 192 - 0xc0
      13'hD6C: dout  = 8'b11001000; // 3436 : 200 - 0xc8
      13'hD6D: dout  = 8'b11111000; // 3437 : 248 - 0xf8
      13'hD6E: dout  = 8'b11111100; // 3438 : 252 - 0xfc
      13'hD6F: dout  = 8'b10011100; // 3439 : 156 - 0x9c
      13'hD70: dout  = 8'b11110010; // 3440 : 242 - 0xf2 -- Sprite 0xd7
      13'hD71: dout  = 8'b11110010; // 3441 : 242 - 0xf2
      13'hD72: dout  = 8'b11110100; // 3442 : 244 - 0xf4
      13'hD73: dout  = 8'b11110111; // 3443 : 247 - 0xf7
      13'hD74: dout  = 8'b11111101; // 3444 : 253 - 0xfd
      13'hD75: dout  = 8'b11100001; // 3445 : 225 - 0xe1
      13'hD76: dout  = 8'b00010010; // 3446 :  18 - 0x12
      13'hD77: dout  = 8'b00001100; // 3447 :  12 - 0xc
      13'hD78: dout  = 8'b00001100; // 3448 :  12 - 0xc
      13'hD79: dout  = 8'b10011100; // 3449 : 156 - 0x9c
      13'hD7A: dout  = 8'b11111000; // 3450 : 248 - 0xf8
      13'hD7B: dout  = 8'b01111000; // 3451 : 120 - 0x78
      13'hD7C: dout  = 8'b11100010; // 3452 : 226 - 0xe2
      13'hD7D: dout  = 8'b00011110; // 3453 :  30 - 0x1e
      13'hD7E: dout  = 8'b00001100; // 3454 :  12 - 0xc
      13'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      13'hD80: dout  = 8'b01111000; // 3456 : 120 - 0x78 -- Sprite 0xd8
      13'hD81: dout  = 8'b01001110; // 3457 :  78 - 0x4e
      13'hD82: dout  = 8'b11000010; // 3458 : 194 - 0xc2
      13'hD83: dout  = 8'b10011010; // 3459 : 154 - 0x9a
      13'hD84: dout  = 8'b10011011; // 3460 : 155 - 0x9b
      13'hD85: dout  = 8'b11011001; // 3461 : 217 - 0xd9
      13'hD86: dout  = 8'b01100011; // 3462 :  99 - 0x63
      13'hD87: dout  = 8'b00111110; // 3463 :  62 - 0x3e
      13'hD88: dout  = 8'b00000000; // 3464 :   0 - 0x0
      13'hD89: dout  = 8'b00110000; // 3465 :  48 - 0x30
      13'hD8A: dout  = 8'b00111100; // 3466 :  60 - 0x3c
      13'hD8B: dout  = 8'b01111100; // 3467 : 124 - 0x7c
      13'hD8C: dout  = 8'b01111100; // 3468 : 124 - 0x7c
      13'hD8D: dout  = 8'b00111110; // 3469 :  62 - 0x3e
      13'hD8E: dout  = 8'b00011100; // 3470 :  28 - 0x1c
      13'hD8F: dout  = 8'b00000000; // 3471 :   0 - 0x0
      13'hD90: dout  = 8'b00011110; // 3472 :  30 - 0x1e -- Sprite 0xd9
      13'hD91: dout  = 8'b01110001; // 3473 : 113 - 0x71
      13'hD92: dout  = 8'b01001001; // 3474 :  73 - 0x49
      13'hD93: dout  = 8'b10111001; // 3475 : 185 - 0xb9
      13'hD94: dout  = 8'b10011101; // 3476 : 157 - 0x9d
      13'hD95: dout  = 8'b01010010; // 3477 :  82 - 0x52
      13'hD96: dout  = 8'b01110010; // 3478 : 114 - 0x72
      13'hD97: dout  = 8'b00011110; // 3479 :  30 - 0x1e
      13'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0
      13'hD99: dout  = 8'b00001110; // 3481 :  14 - 0xe
      13'hD9A: dout  = 8'b00111110; // 3482 :  62 - 0x3e
      13'hD9B: dout  = 8'b01111110; // 3483 : 126 - 0x7e
      13'hD9C: dout  = 8'b01111110; // 3484 : 126 - 0x7e
      13'hD9D: dout  = 8'b00111100; // 3485 :  60 - 0x3c
      13'hD9E: dout  = 8'b00001100; // 3486 :  12 - 0xc
      13'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      13'hDA0: dout  = 8'b01100000; // 3488 :  96 - 0x60 -- Sprite 0xda
      13'hDA1: dout  = 8'b01011110; // 3489 :  94 - 0x5e
      13'hDA2: dout  = 8'b10001001; // 3490 : 137 - 0x89
      13'hDA3: dout  = 8'b10111101; // 3491 : 189 - 0xbd
      13'hDA4: dout  = 8'b10011101; // 3492 : 157 - 0x9d
      13'hDA5: dout  = 8'b11010011; // 3493 : 211 - 0xd3
      13'hDA6: dout  = 8'b01000110; // 3494 :  70 - 0x46
      13'hDA7: dout  = 8'b01111100; // 3495 : 124 - 0x7c
      13'hDA8: dout  = 8'b00000000; // 3496 :   0 - 0x0
      13'hDA9: dout  = 8'b00100000; // 3497 :  32 - 0x20
      13'hDAA: dout  = 8'b01111110; // 3498 : 126 - 0x7e
      13'hDAB: dout  = 8'b01111110; // 3499 : 126 - 0x7e
      13'hDAC: dout  = 8'b01111110; // 3500 : 126 - 0x7e
      13'hDAD: dout  = 8'b00111100; // 3501 :  60 - 0x3c
      13'hDAE: dout  = 8'b00111000; // 3502 :  56 - 0x38
      13'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout  = 8'b00011110; // 3504 :  30 - 0x1e -- Sprite 0xdb
      13'hDB1: dout  = 8'b00100011; // 3505 :  35 - 0x23
      13'hDB2: dout  = 8'b01001001; // 3506 :  73 - 0x49
      13'hDB3: dout  = 8'b10111101; // 3507 : 189 - 0xbd
      13'hDB4: dout  = 8'b10011001; // 3508 : 153 - 0x99
      13'hDB5: dout  = 8'b01000011; // 3509 :  67 - 0x43
      13'hDB6: dout  = 8'b01101110; // 3510 : 110 - 0x6e
      13'hDB7: dout  = 8'b00011000; // 3511 :  24 - 0x18
      13'hDB8: dout  = 8'b00000000; // 3512 :   0 - 0x0
      13'hDB9: dout  = 8'b00011100; // 3513 :  28 - 0x1c
      13'hDBA: dout  = 8'b00111110; // 3514 :  62 - 0x3e
      13'hDBB: dout  = 8'b01111110; // 3515 : 126 - 0x7e
      13'hDBC: dout  = 8'b01111110; // 3516 : 126 - 0x7e
      13'hDBD: dout  = 8'b00111100; // 3517 :  60 - 0x3c
      13'hDBE: dout  = 8'b00010000; // 3518 :  16 - 0x10
      13'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      13'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      13'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      13'hDC2: dout  = 8'b00000001; // 3522 :   1 - 0x1
      13'hDC3: dout  = 8'b00000010; // 3523 :   2 - 0x2
      13'hDC4: dout  = 8'b00000100; // 3524 :   4 - 0x4
      13'hDC5: dout  = 8'b00000010; // 3525 :   2 - 0x2
      13'hDC6: dout  = 8'b00011110; // 3526 :  30 - 0x1e
      13'hDC7: dout  = 8'b00010000; // 3527 :  16 - 0x10
      13'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0
      13'hDC9: dout  = 8'b00000000; // 3529 :   0 - 0x0
      13'hDCA: dout  = 8'b00000000; // 3530 :   0 - 0x0
      13'hDCB: dout  = 8'b00000001; // 3531 :   1 - 0x1
      13'hDCC: dout  = 8'b00000011; // 3532 :   3 - 0x3
      13'hDCD: dout  = 8'b00000001; // 3533 :   1 - 0x1
      13'hDCE: dout  = 8'b00000001; // 3534 :   1 - 0x1
      13'hDCF: dout  = 8'b00001111; // 3535 :  15 - 0xf
      13'hDD0: dout  = 8'b00001000; // 3536 :   8 - 0x8 -- Sprite 0xdd
      13'hDD1: dout  = 8'b00001101; // 3537 :  13 - 0xd
      13'hDD2: dout  = 8'b00111010; // 3538 :  58 - 0x3a
      13'hDD3: dout  = 8'b00100101; // 3539 :  37 - 0x25
      13'hDD4: dout  = 8'b00011011; // 3540 :  27 - 0x1b
      13'hDD5: dout  = 8'b00001111; // 3541 :  15 - 0xf
      13'hDD6: dout  = 8'b00000111; // 3542 :   7 - 0x7
      13'hDD7: dout  = 8'b00000011; // 3543 :   3 - 0x3
      13'hDD8: dout  = 8'b00000111; // 3544 :   7 - 0x7
      13'hDD9: dout  = 8'b00000111; // 3545 :   7 - 0x7
      13'hDDA: dout  = 8'b00000111; // 3546 :   7 - 0x7
      13'hDDB: dout  = 8'b00011111; // 3547 :  31 - 0x1f
      13'hDDC: dout  = 8'b00001111; // 3548 :  15 - 0xf
      13'hDDD: dout  = 8'b00000111; // 3549 :   7 - 0x7
      13'hDDE: dout  = 8'b00000011; // 3550 :   3 - 0x3
      13'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      13'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Sprite 0xde
      13'hDE1: dout  = 8'b00000000; // 3553 :   0 - 0x0
      13'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      13'hDE3: dout  = 8'b11000000; // 3555 : 192 - 0xc0
      13'hDE4: dout  = 8'b01000000; // 3556 :  64 - 0x40
      13'hDE5: dout  = 8'b01011000; // 3557 :  88 - 0x58
      13'hDE6: dout  = 8'b01101000; // 3558 : 104 - 0x68
      13'hDE7: dout  = 8'b00001000; // 3559 :   8 - 0x8
      13'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0
      13'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      13'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      13'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      13'hDEC: dout  = 8'b10000000; // 3564 : 128 - 0x80
      13'hDED: dout  = 8'b10000000; // 3565 : 128 - 0x80
      13'hDEE: dout  = 8'b10010000; // 3566 : 144 - 0x90
      13'hDEF: dout  = 8'b11110000; // 3567 : 240 - 0xf0
      13'hDF0: dout  = 8'b00010000; // 3568 :  16 - 0x10 -- Sprite 0xdf
      13'hDF1: dout  = 8'b01011100; // 3569 :  92 - 0x5c
      13'hDF2: dout  = 8'b10101000; // 3570 : 168 - 0xa8
      13'hDF3: dout  = 8'b11011000; // 3571 : 216 - 0xd8
      13'hDF4: dout  = 8'b10111000; // 3572 : 184 - 0xb8
      13'hDF5: dout  = 8'b11110000; // 3573 : 240 - 0xf0
      13'hDF6: dout  = 8'b11100000; // 3574 : 224 - 0xe0
      13'hDF7: dout  = 8'b11000000; // 3575 : 192 - 0xc0
      13'hDF8: dout  = 8'b11100000; // 3576 : 224 - 0xe0
      13'hDF9: dout  = 8'b11100000; // 3577 : 224 - 0xe0
      13'hDFA: dout  = 8'b11110000; // 3578 : 240 - 0xf0
      13'hDFB: dout  = 8'b11110000; // 3579 : 240 - 0xf0
      13'hDFC: dout  = 8'b11100000; // 3580 : 224 - 0xe0
      13'hDFD: dout  = 8'b11000000; // 3581 : 192 - 0xc0
      13'hDFE: dout  = 8'b11000000; // 3582 : 192 - 0xc0
      13'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      13'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Sprite 0xe0
      13'hE01: dout  = 8'b00000000; // 3585 :   0 - 0x0
      13'hE02: dout  = 8'b00000000; // 3586 :   0 - 0x0
      13'hE03: dout  = 8'b00010011; // 3587 :  19 - 0x13
      13'hE04: dout  = 8'b00010011; // 3588 :  19 - 0x13
      13'hE05: dout  = 8'b00110111; // 3589 :  55 - 0x37
      13'hE06: dout  = 8'b00110111; // 3590 :  55 - 0x37
      13'hE07: dout  = 8'b00000111; // 3591 :   7 - 0x7
      13'hE08: dout  = 8'b00001111; // 3592 :  15 - 0xf
      13'hE09: dout  = 8'b00011111; // 3593 :  31 - 0x1f
      13'hE0A: dout  = 8'b00011111; // 3594 :  31 - 0x1f
      13'hE0B: dout  = 8'b00111111; // 3595 :  63 - 0x3f
      13'hE0C: dout  = 8'b01111111; // 3596 : 127 - 0x7f
      13'hE0D: dout  = 8'b11111111; // 3597 : 255 - 0xff
      13'hE0E: dout  = 8'b11111111; // 3598 : 255 - 0xff
      13'hE0F: dout  = 8'b11111111; // 3599 : 255 - 0xff
      13'hE10: dout  = 8'b00000111; // 3600 :   7 - 0x7 -- Sprite 0xe1
      13'hE11: dout  = 8'b00000100; // 3601 :   4 - 0x4
      13'hE12: dout  = 8'b00000000; // 3602 :   0 - 0x0
      13'hE13: dout  = 8'b00000000; // 3603 :   0 - 0x0
      13'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      13'hE15: dout  = 8'b00100000; // 3605 :  32 - 0x20
      13'hE16: dout  = 8'b01110000; // 3606 : 112 - 0x70
      13'hE17: dout  = 8'b11111000; // 3607 : 248 - 0xf8
      13'hE18: dout  = 8'b11111111; // 3608 : 255 - 0xff
      13'hE19: dout  = 8'b11111111; // 3609 : 255 - 0xff
      13'hE1A: dout  = 8'b01111111; // 3610 : 127 - 0x7f
      13'hE1B: dout  = 8'b00111111; // 3611 :  63 - 0x3f
      13'hE1C: dout  = 8'b00111111; // 3612 :  63 - 0x3f
      13'hE1D: dout  = 8'b00011111; // 3613 :  31 - 0x1f
      13'hE1E: dout  = 8'b00001111; // 3614 :  15 - 0xf
      13'hE1F: dout  = 8'b00000111; // 3615 :   7 - 0x7
      13'hE20: dout  = 8'b00000000; // 3616 :   0 - 0x0 -- Sprite 0xe2
      13'hE21: dout  = 8'b00000000; // 3617 :   0 - 0x0
      13'hE22: dout  = 8'b00000000; // 3618 :   0 - 0x0
      13'hE23: dout  = 8'b11111000; // 3619 : 248 - 0xf8
      13'hE24: dout  = 8'b11111100; // 3620 : 252 - 0xfc
      13'hE25: dout  = 8'b11111100; // 3621 : 252 - 0xfc
      13'hE26: dout  = 8'b11111100; // 3622 : 252 - 0xfc
      13'hE27: dout  = 8'b11111101; // 3623 : 253 - 0xfd
      13'hE28: dout  = 8'b11111110; // 3624 : 254 - 0xfe
      13'hE29: dout  = 8'b11111111; // 3625 : 255 - 0xff
      13'hE2A: dout  = 8'b11111111; // 3626 : 255 - 0xff
      13'hE2B: dout  = 8'b00001111; // 3627 :  15 - 0xf
      13'hE2C: dout  = 8'b10111111; // 3628 : 191 - 0xbf
      13'hE2D: dout  = 8'b10100011; // 3629 : 163 - 0xa3
      13'hE2E: dout  = 8'b11110111; // 3630 : 247 - 0xf7
      13'hE2F: dout  = 8'b11110111; // 3631 : 247 - 0xf7
      13'hE30: dout  = 8'b11111100; // 3632 : 252 - 0xfc -- Sprite 0xe3
      13'hE31: dout  = 8'b00011100; // 3633 :  28 - 0x1c
      13'hE32: dout  = 8'b11000000; // 3634 : 192 - 0xc0
      13'hE33: dout  = 8'b11100000; // 3635 : 224 - 0xe0
      13'hE34: dout  = 8'b00000000; // 3636 :   0 - 0x0
      13'hE35: dout  = 8'b00000000; // 3637 :   0 - 0x0
      13'hE36: dout  = 8'b00000110; // 3638 :   6 - 0x6
      13'hE37: dout  = 8'b00001111; // 3639 :  15 - 0xf
      13'hE38: dout  = 8'b11111111; // 3640 : 255 - 0xff
      13'hE39: dout  = 8'b11111111; // 3641 : 255 - 0xff
      13'hE3A: dout  = 8'b00111111; // 3642 :  63 - 0x3f
      13'hE3B: dout  = 8'b00011111; // 3643 :  31 - 0x1f
      13'hE3C: dout  = 8'b11111110; // 3644 : 254 - 0xfe
      13'hE3D: dout  = 8'b11111100; // 3645 : 252 - 0xfc
      13'hE3E: dout  = 8'b11111000; // 3646 : 248 - 0xf8
      13'hE3F: dout  = 8'b11110000; // 3647 : 240 - 0xf0
      13'hE40: dout  = 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      13'hE41: dout  = 8'b00000000; // 3649 :   0 - 0x0
      13'hE42: dout  = 8'b00000000; // 3650 :   0 - 0x0
      13'hE43: dout  = 8'b00010011; // 3651 :  19 - 0x13
      13'hE44: dout  = 8'b00010011; // 3652 :  19 - 0x13
      13'hE45: dout  = 8'b00110111; // 3653 :  55 - 0x37
      13'hE46: dout  = 8'b00110111; // 3654 :  55 - 0x37
      13'hE47: dout  = 8'b00000111; // 3655 :   7 - 0x7
      13'hE48: dout  = 8'b00001111; // 3656 :  15 - 0xf
      13'hE49: dout  = 8'b00011111; // 3657 :  31 - 0x1f
      13'hE4A: dout  = 8'b00011111; // 3658 :  31 - 0x1f
      13'hE4B: dout  = 8'b00111111; // 3659 :  63 - 0x3f
      13'hE4C: dout  = 8'b01111111; // 3660 : 127 - 0x7f
      13'hE4D: dout  = 8'b11111111; // 3661 : 255 - 0xff
      13'hE4E: dout  = 8'b11111111; // 3662 : 255 - 0xff
      13'hE4F: dout  = 8'b11111111; // 3663 : 255 - 0xff
      13'hE50: dout  = 8'b00000111; // 3664 :   7 - 0x7 -- Sprite 0xe5
      13'hE51: dout  = 8'b00000100; // 3665 :   4 - 0x4
      13'hE52: dout  = 8'b00000001; // 3666 :   1 - 0x1
      13'hE53: dout  = 8'b00000000; // 3667 :   0 - 0x0
      13'hE54: dout  = 8'b00000000; // 3668 :   0 - 0x0
      13'hE55: dout  = 8'b00100000; // 3669 :  32 - 0x20
      13'hE56: dout  = 8'b01110000; // 3670 : 112 - 0x70
      13'hE57: dout  = 8'b11111000; // 3671 : 248 - 0xf8
      13'hE58: dout  = 8'b11111111; // 3672 : 255 - 0xff
      13'hE59: dout  = 8'b11111111; // 3673 : 255 - 0xff
      13'hE5A: dout  = 8'b01111110; // 3674 : 126 - 0x7e
      13'hE5B: dout  = 8'b00111111; // 3675 :  63 - 0x3f
      13'hE5C: dout  = 8'b00111111; // 3676 :  63 - 0x3f
      13'hE5D: dout  = 8'b00011111; // 3677 :  31 - 0x1f
      13'hE5E: dout  = 8'b00001111; // 3678 :  15 - 0xf
      13'hE5F: dout  = 8'b00000111; // 3679 :   7 - 0x7
      13'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Sprite 0xe6
      13'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      13'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      13'hE63: dout  = 8'b11111100; // 3683 : 252 - 0xfc
      13'hE64: dout  = 8'b11111100; // 3684 : 252 - 0xfc
      13'hE65: dout  = 8'b11111100; // 3685 : 252 - 0xfc
      13'hE66: dout  = 8'b11111100; // 3686 : 252 - 0xfc
      13'hE67: dout  = 8'b11111101; // 3687 : 253 - 0xfd
      13'hE68: dout  = 8'b11111110; // 3688 : 254 - 0xfe
      13'hE69: dout  = 8'b11111111; // 3689 : 255 - 0xff
      13'hE6A: dout  = 8'b11111111; // 3690 : 255 - 0xff
      13'hE6B: dout  = 8'b11100011; // 3691 : 227 - 0xe3
      13'hE6C: dout  = 8'b00010111; // 3692 :  23 - 0x17
      13'hE6D: dout  = 8'b10110111; // 3693 : 183 - 0xb7
      13'hE6E: dout  = 8'b10111111; // 3694 : 191 - 0xbf
      13'hE6F: dout  = 8'b11111111; // 3695 : 255 - 0xff
      13'hE70: dout  = 8'b11111100; // 3696 : 252 - 0xfc -- Sprite 0xe7
      13'hE71: dout  = 8'b00001100; // 3697 :  12 - 0xc
      13'hE72: dout  = 8'b11000000; // 3698 : 192 - 0xc0
      13'hE73: dout  = 8'b11110000; // 3699 : 240 - 0xf0
      13'hE74: dout  = 8'b11110000; // 3700 : 240 - 0xf0
      13'hE75: dout  = 8'b00000000; // 3701 :   0 - 0x0
      13'hE76: dout  = 8'b00000110; // 3702 :   6 - 0x6
      13'hE77: dout  = 8'b00001111; // 3703 :  15 - 0xf
      13'hE78: dout  = 8'b11111111; // 3704 : 255 - 0xff
      13'hE79: dout  = 8'b11111111; // 3705 : 255 - 0xff
      13'hE7A: dout  = 8'b00111111; // 3706 :  63 - 0x3f
      13'hE7B: dout  = 8'b00001111; // 3707 :  15 - 0xf
      13'hE7C: dout  = 8'b00001110; // 3708 :  14 - 0xe
      13'hE7D: dout  = 8'b11111100; // 3709 : 252 - 0xfc
      13'hE7E: dout  = 8'b11111000; // 3710 : 248 - 0xf8
      13'hE7F: dout  = 8'b11110000; // 3711 : 240 - 0xf0
      13'hE80: dout  = 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      13'hE81: dout  = 8'b11111111; // 3713 : 255 - 0xff
      13'hE82: dout  = 8'b01111111; // 3714 : 127 - 0x7f
      13'hE83: dout  = 8'b01111111; // 3715 : 127 - 0x7f
      13'hE84: dout  = 8'b01111111; // 3716 : 127 - 0x7f
      13'hE85: dout  = 8'b00111111; // 3717 :  63 - 0x3f
      13'hE86: dout  = 8'b00111111; // 3718 :  63 - 0x3f
      13'hE87: dout  = 8'b00111111; // 3719 :  63 - 0x3f
      13'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0
      13'hE89: dout  = 8'b00000101; // 3721 :   5 - 0x5
      13'hE8A: dout  = 8'b00000111; // 3722 :   7 - 0x7
      13'hE8B: dout  = 8'b00000011; // 3723 :   3 - 0x3
      13'hE8C: dout  = 8'b00000000; // 3724 :   0 - 0x0
      13'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      13'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      13'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      13'hE90: dout  = 8'b00111100; // 3728 :  60 - 0x3c -- Sprite 0xe9
      13'hE91: dout  = 8'b00111110; // 3729 :  62 - 0x3e
      13'hE92: dout  = 8'b00011111; // 3730 :  31 - 0x1f
      13'hE93: dout  = 8'b00001111; // 3731 :  15 - 0xf
      13'hE94: dout  = 8'b00000111; // 3732 :   7 - 0x7
      13'hE95: dout  = 8'b00000000; // 3733 :   0 - 0x0
      13'hE96: dout  = 8'b00000000; // 3734 :   0 - 0x0
      13'hE97: dout  = 8'b00000000; // 3735 :   0 - 0x0
      13'hE98: dout  = 8'b00000000; // 3736 :   0 - 0x0
      13'hE99: dout  = 8'b00000000; // 3737 :   0 - 0x0
      13'hE9A: dout  = 8'b00000000; // 3738 :   0 - 0x0
      13'hE9B: dout  = 8'b00000000; // 3739 :   0 - 0x0
      13'hE9C: dout  = 8'b00000000; // 3740 :   0 - 0x0
      13'hE9D: dout  = 8'b00000000; // 3741 :   0 - 0x0
      13'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      13'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      13'hEA0: dout  = 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      13'hEA1: dout  = 8'b11111110; // 3745 : 254 - 0xfe
      13'hEA2: dout  = 8'b11111110; // 3746 : 254 - 0xfe
      13'hEA3: dout  = 8'b11111100; // 3747 : 252 - 0xfc
      13'hEA4: dout  = 8'b11111000; // 3748 : 248 - 0xf8
      13'hEA5: dout  = 8'b11110000; // 3749 : 240 - 0xf0
      13'hEA6: dout  = 8'b10110000; // 3750 : 176 - 0xb0
      13'hEA7: dout  = 8'b00111001; // 3751 :  57 - 0x39
      13'hEA8: dout  = 8'b00000011; // 3752 :   3 - 0x3
      13'hEA9: dout  = 8'b10011110; // 3753 : 158 - 0x9e
      13'hEAA: dout  = 8'b00001110; // 3754 :  14 - 0xe
      13'hEAB: dout  = 8'b00000000; // 3755 :   0 - 0x0
      13'hEAC: dout  = 8'b00000000; // 3756 :   0 - 0x0
      13'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      13'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      13'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout  = 8'b00011111; // 3760 :  31 - 0x1f -- Sprite 0xeb
      13'hEB1: dout  = 8'b11001111; // 3761 : 207 - 0xcf
      13'hEB2: dout  = 8'b11000110; // 3762 : 198 - 0xc6
      13'hEB3: dout  = 8'b10000000; // 3763 : 128 - 0x80
      13'hEB4: dout  = 8'b00000000; // 3764 :   0 - 0x0
      13'hEB5: dout  = 8'b00000000; // 3765 :   0 - 0x0
      13'hEB6: dout  = 8'b00000000; // 3766 :   0 - 0x0
      13'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      13'hEB8: dout  = 8'b00000000; // 3768 :   0 - 0x0
      13'hEB9: dout  = 8'b00000000; // 3769 :   0 - 0x0
      13'hEBA: dout  = 8'b00000000; // 3770 :   0 - 0x0
      13'hEBB: dout  = 8'b00000000; // 3771 :   0 - 0x0
      13'hEBC: dout  = 8'b00000000; // 3772 :   0 - 0x0
      13'hEBD: dout  = 8'b00000000; // 3773 :   0 - 0x0
      13'hEBE: dout  = 8'b00000000; // 3774 :   0 - 0x0
      13'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      13'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout  = 8'b00000000; // 3777 :   0 - 0x0
      13'hEC2: dout  = 8'b00000000; // 3778 :   0 - 0x0
      13'hEC3: dout  = 8'b00000000; // 3779 :   0 - 0x0
      13'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      13'hEC5: dout  = 8'b00000000; // 3781 :   0 - 0x0
      13'hEC6: dout  = 8'b00001100; // 3782 :  12 - 0xc
      13'hEC7: dout  = 8'b00001100; // 3783 :  12 - 0xc
      13'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout  = 8'b00000000; // 3785 :   0 - 0x0
      13'hECA: dout  = 8'b00000000; // 3786 :   0 - 0x0
      13'hECB: dout  = 8'b00000000; // 3787 :   0 - 0x0
      13'hECC: dout  = 8'b00000100; // 3788 :   4 - 0x4
      13'hECD: dout  = 8'b00001110; // 3789 :  14 - 0xe
      13'hECE: dout  = 8'b00001111; // 3790 :  15 - 0xf
      13'hECF: dout  = 8'b00001011; // 3791 :  11 - 0xb
      13'hED0: dout  = 8'b00110000; // 3792 :  48 - 0x30 -- Sprite 0xed
      13'hED1: dout  = 8'b01000011; // 3793 :  67 - 0x43
      13'hED2: dout  = 8'b01000000; // 3794 :  64 - 0x40
      13'hED3: dout  = 8'b01100000; // 3795 :  96 - 0x60
      13'hED4: dout  = 8'b00000011; // 3796 :   3 - 0x3
      13'hED5: dout  = 8'b00000000; // 3797 :   0 - 0x0
      13'hED6: dout  = 8'b01111111; // 3798 : 127 - 0x7f
      13'hED7: dout  = 8'b00000000; // 3799 :   0 - 0x0
      13'hED8: dout  = 8'b00001111; // 3800 :  15 - 0xf
      13'hED9: dout  = 8'b00001100; // 3801 :  12 - 0xc
      13'hEDA: dout  = 8'b00001111; // 3802 :  15 - 0xf
      13'hEDB: dout  = 8'b00001111; // 3803 :  15 - 0xf
      13'hEDC: dout  = 8'b00000000; // 3804 :   0 - 0x0
      13'hEDD: dout  = 8'b01111111; // 3805 : 127 - 0x7f
      13'hEDE: dout  = 8'b11010101; // 3806 : 213 - 0xd5
      13'hEDF: dout  = 8'b01111111; // 3807 : 127 - 0x7f
      13'hEE0: dout  = 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      13'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      13'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      13'hEE3: dout  = 8'b00000000; // 3811 :   0 - 0x0
      13'hEE4: dout  = 8'b00000000; // 3812 :   0 - 0x0
      13'hEE5: dout  = 8'b00000000; // 3813 :   0 - 0x0
      13'hEE6: dout  = 8'b00110000; // 3814 :  48 - 0x30
      13'hEE7: dout  = 8'b00110000; // 3815 :  48 - 0x30
      13'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0
      13'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout  = 8'b00000000; // 3818 :   0 - 0x0
      13'hEEB: dout  = 8'b00000000; // 3819 :   0 - 0x0
      13'hEEC: dout  = 8'b00100000; // 3820 :  32 - 0x20
      13'hEED: dout  = 8'b01110000; // 3821 : 112 - 0x70
      13'hEEE: dout  = 8'b11110000; // 3822 : 240 - 0xf0
      13'hEEF: dout  = 8'b11100000; // 3823 : 224 - 0xe0
      13'hEF0: dout  = 8'b00001110; // 3824 :  14 - 0xe -- Sprite 0xef
      13'hEF1: dout  = 8'b11001011; // 3825 : 203 - 0xcb
      13'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      13'hEF3: dout  = 8'b00000000; // 3827 :   0 - 0x0
      13'hEF4: dout  = 8'b11000000; // 3828 : 192 - 0xc0
      13'hEF5: dout  = 8'b00000000; // 3829 :   0 - 0x0
      13'hEF6: dout  = 8'b11111110; // 3830 : 254 - 0xfe
      13'hEF7: dout  = 8'b00000000; // 3831 :   0 - 0x0
      13'hEF8: dout  = 8'b11110000; // 3832 : 240 - 0xf0
      13'hEF9: dout  = 8'b00110000; // 3833 :  48 - 0x30
      13'hEFA: dout  = 8'b11110000; // 3834 : 240 - 0xf0
      13'hEFB: dout  = 8'b11110000; // 3835 : 240 - 0xf0
      13'hEFC: dout  = 8'b00000000; // 3836 :   0 - 0x0
      13'hEFD: dout  = 8'b11111110; // 3837 : 254 - 0xfe
      13'hEFE: dout  = 8'b01010101; // 3838 :  85 - 0x55
      13'hEFF: dout  = 8'b11111110; // 3839 : 254 - 0xfe
      13'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      13'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      13'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      13'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      13'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      13'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      13'hF06: dout  = 8'b00001100; // 3846 :  12 - 0xc
      13'hF07: dout  = 8'b00001100; // 3847 :  12 - 0xc
      13'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0
      13'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      13'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      13'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      13'hF0C: dout  = 8'b00000100; // 3852 :   4 - 0x4
      13'hF0D: dout  = 8'b00001110; // 3853 :  14 - 0xe
      13'hF0E: dout  = 8'b00001111; // 3854 :  15 - 0xf
      13'hF0F: dout  = 8'b00001011; // 3855 :  11 - 0xb
      13'hF10: dout  = 8'b00110000; // 3856 :  48 - 0x30 -- Sprite 0xf1
      13'hF11: dout  = 8'b00100011; // 3857 :  35 - 0x23
      13'hF12: dout  = 8'b00100000; // 3858 :  32 - 0x20
      13'hF13: dout  = 8'b01100000; // 3859 :  96 - 0x60
      13'hF14: dout  = 8'b00000011; // 3860 :   3 - 0x3
      13'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      13'hF16: dout  = 8'b01111111; // 3862 : 127 - 0x7f
      13'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout  = 8'b00001111; // 3864 :  15 - 0xf
      13'hF19: dout  = 8'b00001100; // 3865 :  12 - 0xc
      13'hF1A: dout  = 8'b00001111; // 3866 :  15 - 0xf
      13'hF1B: dout  = 8'b00001111; // 3867 :  15 - 0xf
      13'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      13'hF1D: dout  = 8'b01111111; // 3869 : 127 - 0x7f
      13'hF1E: dout  = 8'b10101010; // 3870 : 170 - 0xaa
      13'hF1F: dout  = 8'b01111111; // 3871 : 127 - 0x7f
      13'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      13'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      13'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      13'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      13'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      13'hF26: dout  = 8'b00110000; // 3878 :  48 - 0x30
      13'hF27: dout  = 8'b00110000; // 3879 :  48 - 0x30
      13'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0
      13'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      13'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      13'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      13'hF2C: dout  = 8'b00100000; // 3884 :  32 - 0x20
      13'hF2D: dout  = 8'b01110000; // 3885 : 112 - 0x70
      13'hF2E: dout  = 8'b11110000; // 3886 : 240 - 0xf0
      13'hF2F: dout  = 8'b11100000; // 3887 : 224 - 0xe0
      13'hF30: dout  = 8'b00001001; // 3888 :   9 - 0x9 -- Sprite 0xf3
      13'hF31: dout  = 8'b11001111; // 3889 : 207 - 0xcf
      13'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      13'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      13'hF34: dout  = 8'b11000000; // 3892 : 192 - 0xc0
      13'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      13'hF36: dout  = 8'b11111110; // 3894 : 254 - 0xfe
      13'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      13'hF38: dout  = 8'b11110000; // 3896 : 240 - 0xf0
      13'hF39: dout  = 8'b00110000; // 3897 :  48 - 0x30
      13'hF3A: dout  = 8'b11110000; // 3898 : 240 - 0xf0
      13'hF3B: dout  = 8'b11110000; // 3899 : 240 - 0xf0
      13'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      13'hF3D: dout  = 8'b11111110; // 3901 : 254 - 0xfe
      13'hF3E: dout  = 8'b10101011; // 3902 : 171 - 0xab
      13'hF3F: dout  = 8'b11111110; // 3903 : 254 - 0xfe
      13'hF40: dout  = 8'b00111111; // 3904 :  63 - 0x3f -- Sprite 0xf4
      13'hF41: dout  = 8'b00110101; // 3905 :  53 - 0x35
      13'hF42: dout  = 8'b00011010; // 3906 :  26 - 0x1a
      13'hF43: dout  = 8'b00001101; // 3907 :  13 - 0xd
      13'hF44: dout  = 8'b00001010; // 3908 :  10 - 0xa
      13'hF45: dout  = 8'b00001101; // 3909 :  13 - 0xd
      13'hF46: dout  = 8'b00001000; // 3910 :   8 - 0x8
      13'hF47: dout  = 8'b00111000; // 3911 :  56 - 0x38
      13'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0
      13'hF49: dout  = 8'b00010101; // 3913 :  21 - 0x15
      13'hF4A: dout  = 8'b00001010; // 3914 :  10 - 0xa
      13'hF4B: dout  = 8'b00000101; // 3915 :   5 - 0x5
      13'hF4C: dout  = 8'b00000010; // 3916 :   2 - 0x2
      13'hF4D: dout  = 8'b00000101; // 3917 :   5 - 0x5
      13'hF4E: dout  = 8'b00000111; // 3918 :   7 - 0x7
      13'hF4F: dout  = 8'b00000111; // 3919 :   7 - 0x7
      13'hF50: dout  = 8'b01110011; // 3920 : 115 - 0x73 -- Sprite 0xf5
      13'hF51: dout  = 8'b11000100; // 3921 : 196 - 0xc4
      13'hF52: dout  = 8'b11000100; // 3922 : 196 - 0xc4
      13'hF53: dout  = 8'b11000000; // 3923 : 192 - 0xc0
      13'hF54: dout  = 8'b11000001; // 3924 : 193 - 0xc1
      13'hF55: dout  = 8'b11000000; // 3925 : 192 - 0xc0
      13'hF56: dout  = 8'b01100001; // 3926 :  97 - 0x61
      13'hF57: dout  = 8'b00111111; // 3927 :  63 - 0x3f
      13'hF58: dout  = 8'b00111100; // 3928 :  60 - 0x3c
      13'hF59: dout  = 8'b01111011; // 3929 : 123 - 0x7b
      13'hF5A: dout  = 8'b01111011; // 3930 : 123 - 0x7b
      13'hF5B: dout  = 8'b01111111; // 3931 : 127 - 0x7f
      13'hF5C: dout  = 8'b01111110; // 3932 : 126 - 0x7e
      13'hF5D: dout  = 8'b01111111; // 3933 : 127 - 0x7f
      13'hF5E: dout  = 8'b00111110; // 3934 :  62 - 0x3e
      13'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout  = 8'b11111100; // 3936 : 252 - 0xfc -- Sprite 0xf6
      13'hF61: dout  = 8'b01010100; // 3937 :  84 - 0x54
      13'hF62: dout  = 8'b10101000; // 3938 : 168 - 0xa8
      13'hF63: dout  = 8'b01010000; // 3939 :  80 - 0x50
      13'hF64: dout  = 8'b10110000; // 3940 : 176 - 0xb0
      13'hF65: dout  = 8'b01010000; // 3941 :  80 - 0x50
      13'hF66: dout  = 8'b10010000; // 3942 : 144 - 0x90
      13'hF67: dout  = 8'b00011100; // 3943 :  28 - 0x1c
      13'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0
      13'hF69: dout  = 8'b01010000; // 3945 :  80 - 0x50
      13'hF6A: dout  = 8'b10100000; // 3946 : 160 - 0xa0
      13'hF6B: dout  = 8'b01000000; // 3947 :  64 - 0x40
      13'hF6C: dout  = 8'b10100000; // 3948 : 160 - 0xa0
      13'hF6D: dout  = 8'b01000000; // 3949 :  64 - 0x40
      13'hF6E: dout  = 8'b11100000; // 3950 : 224 - 0xe0
      13'hF6F: dout  = 8'b11100000; // 3951 : 224 - 0xe0
      13'hF70: dout  = 8'b10000110; // 3952 : 134 - 0x86 -- Sprite 0xf7
      13'hF71: dout  = 8'b01000010; // 3953 :  66 - 0x42
      13'hF72: dout  = 8'b01000111; // 3954 :  71 - 0x47
      13'hF73: dout  = 8'b01000001; // 3955 :  65 - 0x41
      13'hF74: dout  = 8'b10000011; // 3956 : 131 - 0x83
      13'hF75: dout  = 8'b00000001; // 3957 :   1 - 0x1
      13'hF76: dout  = 8'b10000110; // 3958 : 134 - 0x86
      13'hF77: dout  = 8'b11111100; // 3959 : 252 - 0xfc
      13'hF78: dout  = 8'b01111000; // 3960 : 120 - 0x78
      13'hF79: dout  = 8'b10111100; // 3961 : 188 - 0xbc
      13'hF7A: dout  = 8'b10111000; // 3962 : 184 - 0xb8
      13'hF7B: dout  = 8'b10111110; // 3963 : 190 - 0xbe
      13'hF7C: dout  = 8'b01111100; // 3964 : 124 - 0x7c
      13'hF7D: dout  = 8'b11111110; // 3965 : 254 - 0xfe
      13'hF7E: dout  = 8'b01111000; // 3966 : 120 - 0x78
      13'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      13'hF80: dout  = 8'b11100100; // 3968 : 228 - 0xe4 -- Sprite 0xf8
      13'hF81: dout  = 8'b11100100; // 3969 : 228 - 0xe4
      13'hF82: dout  = 8'b11101111; // 3970 : 239 - 0xef
      13'hF83: dout  = 8'b11101111; // 3971 : 239 - 0xef
      13'hF84: dout  = 8'b11111111; // 3972 : 255 - 0xff
      13'hF85: dout  = 8'b11111111; // 3973 : 255 - 0xff
      13'hF86: dout  = 8'b01111111; // 3974 : 127 - 0x7f
      13'hF87: dout  = 8'b01111111; // 3975 : 127 - 0x7f
      13'hF88: dout  = 8'b00000011; // 3976 :   3 - 0x3
      13'hF89: dout  = 8'b00000011; // 3977 :   3 - 0x3
      13'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      13'hF8B: dout  = 8'b00000011; // 3979 :   3 - 0x3
      13'hF8C: dout  = 8'b00000111; // 3980 :   7 - 0x7
      13'hF8D: dout  = 8'b00000110; // 3981 :   6 - 0x6
      13'hF8E: dout  = 8'b00000111; // 3982 :   7 - 0x7
      13'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      13'hF90: dout  = 8'b00111111; // 3984 :  63 - 0x3f -- Sprite 0xf9
      13'hF91: dout  = 8'b01111111; // 3985 : 127 - 0x7f
      13'hF92: dout  = 8'b01111111; // 3986 : 127 - 0x7f
      13'hF93: dout  = 8'b11111111; // 3987 : 255 - 0xff
      13'hF94: dout  = 8'b11111111; // 3988 : 255 - 0xff
      13'hF95: dout  = 8'b11111111; // 3989 : 255 - 0xff
      13'hF96: dout  = 8'b11111111; // 3990 : 255 - 0xff
      13'hF97: dout  = 8'b11111111; // 3991 : 255 - 0xff
      13'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0
      13'hF99: dout  = 8'b00011111; // 3993 :  31 - 0x1f
      13'hF9A: dout  = 8'b00011111; // 3994 :  31 - 0x1f
      13'hF9B: dout  = 8'b00001111; // 3995 :  15 - 0xf
      13'hF9C: dout  = 8'b00000011; // 3996 :   3 - 0x3
      13'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      13'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      13'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      13'hFA0: dout  = 8'b00010011; // 4000 :  19 - 0x13 -- Sprite 0xfa
      13'hFA1: dout  = 8'b00010011; // 4001 :  19 - 0x13
      13'hFA2: dout  = 8'b11111011; // 4002 : 251 - 0xfb
      13'hFA3: dout  = 8'b11111011; // 4003 : 251 - 0xfb
      13'hFA4: dout  = 8'b11111111; // 4004 : 255 - 0xff
      13'hFA5: dout  = 8'b11111111; // 4005 : 255 - 0xff
      13'hFA6: dout  = 8'b11111110; // 4006 : 254 - 0xfe
      13'hFA7: dout  = 8'b11111110; // 4007 : 254 - 0xfe
      13'hFA8: dout  = 8'b11100000; // 4008 : 224 - 0xe0
      13'hFA9: dout  = 8'b11100000; // 4009 : 224 - 0xe0
      13'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      13'hFAB: dout  = 8'b00110000; // 4011 :  48 - 0x30
      13'hFAC: dout  = 8'b01110000; // 4012 : 112 - 0x70
      13'hFAD: dout  = 8'b01100000; // 4013 :  96 - 0x60
      13'hFAE: dout  = 8'b01110000; // 4014 : 112 - 0x70
      13'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      13'hFB0: dout  = 8'b11111110; // 4016 : 254 - 0xfe -- Sprite 0xfb
      13'hFB1: dout  = 8'b11111111; // 4017 : 255 - 0xff
      13'hFB2: dout  = 8'b11111111; // 4018 : 255 - 0xff
      13'hFB3: dout  = 8'b11111111; // 4019 : 255 - 0xff
      13'hFB4: dout  = 8'b11111111; // 4020 : 255 - 0xff
      13'hFB5: dout  = 8'b11111111; // 4021 : 255 - 0xff
      13'hFB6: dout  = 8'b11111111; // 4022 : 255 - 0xff
      13'hFB7: dout  = 8'b11111111; // 4023 : 255 - 0xff
      13'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0
      13'hFB9: dout  = 8'b11111000; // 4025 : 248 - 0xf8
      13'hFBA: dout  = 8'b11111000; // 4026 : 248 - 0xf8
      13'hFBB: dout  = 8'b11110000; // 4027 : 240 - 0xf0
      13'hFBC: dout  = 8'b11000000; // 4028 : 192 - 0xc0
      13'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      13'hFBE: dout  = 8'b00000000; // 4030 :   0 - 0x0
      13'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      13'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      13'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      13'hFC2: dout  = 8'b01111100; // 4034 : 124 - 0x7c
      13'hFC3: dout  = 8'b11111110; // 4035 : 254 - 0xfe
      13'hFC4: dout  = 8'b11111110; // 4036 : 254 - 0xfe
      13'hFC5: dout  = 8'b01111100; // 4037 : 124 - 0x7c
      13'hFC6: dout  = 8'b01000100; // 4038 :  68 - 0x44
      13'hFC7: dout  = 8'b10000010; // 4039 : 130 - 0x82
      13'hFC8: dout  = 8'b00111000; // 4040 :  56 - 0x38
      13'hFC9: dout  = 8'b00111000; // 4041 :  56 - 0x38
      13'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      13'hFCB: dout  = 8'b01111100; // 4043 : 124 - 0x7c
      13'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      13'hFCD: dout  = 8'b00111000; // 4045 :  56 - 0x38
      13'hFCE: dout  = 8'b00111000; // 4046 :  56 - 0x38
      13'hFCF: dout  = 8'b01111100; // 4047 : 124 - 0x7c
      13'hFD0: dout  = 8'b10000010; // 4048 : 130 - 0x82 -- Sprite 0xfd
      13'hFD1: dout  = 8'b10000010; // 4049 : 130 - 0x82
      13'hFD2: dout  = 8'b10000010; // 4050 : 130 - 0x82
      13'hFD3: dout  = 8'b11000110; // 4051 : 198 - 0xc6
      13'hFD4: dout  = 8'b11111110; // 4052 : 254 - 0xfe
      13'hFD5: dout  = 8'b11111110; // 4053 : 254 - 0xfe
      13'hFD6: dout  = 8'b10111010; // 4054 : 186 - 0xba
      13'hFD7: dout  = 8'b01111100; // 4055 : 124 - 0x7c
      13'hFD8: dout  = 8'b01111100; // 4056 : 124 - 0x7c
      13'hFD9: dout  = 8'b01111100; // 4057 : 124 - 0x7c
      13'hFDA: dout  = 8'b01111100; // 4058 : 124 - 0x7c
      13'hFDB: dout  = 8'b00111000; // 4059 :  56 - 0x38
      13'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      13'hFDD: dout  = 8'b01111100; // 4061 : 124 - 0x7c
      13'hFDE: dout  = 8'b01111100; // 4062 : 124 - 0x7c
      13'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      13'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      13'hFE1: dout  = 8'b00011001; // 4065 :  25 - 0x19
      13'hFE2: dout  = 8'b00111110; // 4066 :  62 - 0x3e
      13'hFE3: dout  = 8'b00111100; // 4067 :  60 - 0x3c
      13'hFE4: dout  = 8'b00111100; // 4068 :  60 - 0x3c
      13'hFE5: dout  = 8'b00111100; // 4069 :  60 - 0x3c
      13'hFE6: dout  = 8'b00111110; // 4070 :  62 - 0x3e
      13'hFE7: dout  = 8'b00011001; // 4071 :  25 - 0x19
      13'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0
      13'hFE9: dout  = 8'b00000000; // 4073 :   0 - 0x0
      13'hFEA: dout  = 8'b00010001; // 4074 :  17 - 0x11
      13'hFEB: dout  = 8'b11010111; // 4075 : 215 - 0xd7
      13'hFEC: dout  = 8'b11010111; // 4076 : 215 - 0xd7
      13'hFED: dout  = 8'b11010111; // 4077 : 215 - 0xd7
      13'hFEE: dout  = 8'b00010001; // 4078 :  17 - 0x11
      13'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      13'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      13'hFF1: dout  = 8'b11111110; // 4081 : 254 - 0xfe
      13'hFF2: dout  = 8'b00011101; // 4082 :  29 - 0x1d
      13'hFF3: dout  = 8'b00001111; // 4083 :  15 - 0xf
      13'hFF4: dout  = 8'b00001111; // 4084 :  15 - 0xf
      13'hFF5: dout  = 8'b00001111; // 4085 :  15 - 0xf
      13'hFF6: dout  = 8'b00011101; // 4086 :  29 - 0x1d
      13'hFF7: dout  = 8'b11111110; // 4087 : 254 - 0xfe
      13'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      13'hFFA: dout  = 8'b11100110; // 4090 : 230 - 0xe6
      13'hFFB: dout  = 8'b11110110; // 4091 : 246 - 0xf6
      13'hFFC: dout  = 8'b11110110; // 4092 : 246 - 0xf6
      13'hFFD: dout  = 8'b11110110; // 4093 : 246 - 0xf6
      13'hFFE: dout  = 8'b11100110; // 4094 : 230 - 0xe6
      13'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
          // Pattern Table 1---------
      13'h1000: dout  = 8'b11111111; // 4096 : 255 - 0xff -- Background 0x0
      13'h1001: dout  = 8'b11111111; // 4097 : 255 - 0xff
      13'h1002: dout  = 8'b11000000; // 4098 : 192 - 0xc0
      13'h1003: dout  = 8'b11000000; // 4099 : 192 - 0xc0
      13'h1004: dout  = 8'b11000000; // 4100 : 192 - 0xc0
      13'h1005: dout  = 8'b11000000; // 4101 : 192 - 0xc0
      13'h1006: dout  = 8'b11010101; // 4102 : 213 - 0xd5
      13'h1007: dout  = 8'b11111111; // 4103 : 255 - 0xff
      13'h1008: dout  = 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout  = 8'b01111111; // 4105 : 127 - 0x7f
      13'h100A: dout  = 8'b01111111; // 4106 : 127 - 0x7f
      13'h100B: dout  = 8'b01111111; // 4107 : 127 - 0x7f
      13'h100C: dout  = 8'b01111111; // 4108 : 127 - 0x7f
      13'h100D: dout  = 8'b01111111; // 4109 : 127 - 0x7f
      13'h100E: dout  = 8'b01101010; // 4110 : 106 - 0x6a
      13'h100F: dout  = 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout  = 8'b11111111; // 4112 : 255 - 0xff -- Background 0x1
      13'h1011: dout  = 8'b11111111; // 4113 : 255 - 0xff
      13'h1012: dout  = 8'b11001110; // 4114 : 206 - 0xce
      13'h1013: dout  = 8'b11000110; // 4115 : 198 - 0xc6
      13'h1014: dout  = 8'b11001110; // 4116 : 206 - 0xce
      13'h1015: dout  = 8'b11000110; // 4117 : 198 - 0xc6
      13'h1016: dout  = 8'b11101110; // 4118 : 238 - 0xee
      13'h1017: dout  = 8'b11111111; // 4119 : 255 - 0xff
      13'h1018: dout  = 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout  = 8'b01111011; // 4121 : 123 - 0x7b
      13'h101A: dout  = 8'b01110011; // 4122 : 115 - 0x73
      13'h101B: dout  = 8'b01111011; // 4123 : 123 - 0x7b
      13'h101C: dout  = 8'b01110011; // 4124 : 115 - 0x73
      13'h101D: dout  = 8'b01111011; // 4125 : 123 - 0x7b
      13'h101E: dout  = 8'b01010011; // 4126 :  83 - 0x53
      13'h101F: dout  = 8'b00000000; // 4127 :   0 - 0x0
      13'h1020: dout  = 8'b11111111; // 4128 : 255 - 0xff -- Background 0x2
      13'h1021: dout  = 8'b11111111; // 4129 : 255 - 0xff
      13'h1022: dout  = 8'b01110001; // 4130 : 113 - 0x71
      13'h1023: dout  = 8'b00110011; // 4131 :  51 - 0x33
      13'h1024: dout  = 8'b01110001; // 4132 : 113 - 0x71
      13'h1025: dout  = 8'b00110011; // 4133 :  51 - 0x33
      13'h1026: dout  = 8'b01110101; // 4134 : 117 - 0x75
      13'h1027: dout  = 8'b11111111; // 4135 : 255 - 0xff
      13'h1028: dout  = 8'b00000000; // 4136 :   0 - 0x0
      13'h1029: dout  = 8'b11011110; // 4137 : 222 - 0xde
      13'h102A: dout  = 8'b10011110; // 4138 : 158 - 0x9e
      13'h102B: dout  = 8'b11011100; // 4139 : 220 - 0xdc
      13'h102C: dout  = 8'b10011110; // 4140 : 158 - 0x9e
      13'h102D: dout  = 8'b11011100; // 4141 : 220 - 0xdc
      13'h102E: dout  = 8'b10011010; // 4142 : 154 - 0x9a
      13'h102F: dout  = 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout  = 8'b11111111; // 4144 : 255 - 0xff -- Background 0x3
      13'h1031: dout  = 8'b11111111; // 4145 : 255 - 0xff
      13'h1032: dout  = 8'b00000011; // 4146 :   3 - 0x3
      13'h1033: dout  = 8'b00000001; // 4147 :   1 - 0x1
      13'h1034: dout  = 8'b00000011; // 4148 :   3 - 0x3
      13'h1035: dout  = 8'b00000001; // 4149 :   1 - 0x1
      13'h1036: dout  = 8'b10101011; // 4150 : 171 - 0xab
      13'h1037: dout  = 8'b11111111; // 4151 : 255 - 0xff
      13'h1038: dout  = 8'b00000000; // 4152 :   0 - 0x0
      13'h1039: dout  = 8'b11111110; // 4153 : 254 - 0xfe
      13'h103A: dout  = 8'b11111100; // 4154 : 252 - 0xfc
      13'h103B: dout  = 8'b11111110; // 4155 : 254 - 0xfe
      13'h103C: dout  = 8'b11111100; // 4156 : 252 - 0xfc
      13'h103D: dout  = 8'b11111110; // 4157 : 254 - 0xfe
      13'h103E: dout  = 8'b01010100; // 4158 :  84 - 0x54
      13'h103F: dout  = 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout  = 8'b11111111; // 4160 : 255 - 0xff -- Background 0x4
      13'h1041: dout  = 8'b11111111; // 4161 : 255 - 0xff
      13'h1042: dout  = 8'b11100000; // 4162 : 224 - 0xe0
      13'h1043: dout  = 8'b11000110; // 4163 : 198 - 0xc6
      13'h1044: dout  = 8'b11000110; // 4164 : 198 - 0xc6
      13'h1045: dout  = 8'b11110110; // 4165 : 246 - 0xf6
      13'h1046: dout  = 8'b11110000; // 4166 : 240 - 0xf0
      13'h1047: dout  = 8'b11110001; // 4167 : 241 - 0xf1
      13'h1048: dout  = 8'b00000000; // 4168 :   0 - 0x0
      13'h1049: dout  = 8'b01111111; // 4169 : 127 - 0x7f
      13'h104A: dout  = 8'b01011111; // 4170 :  95 - 0x5f
      13'h104B: dout  = 8'b01111001; // 4171 : 121 - 0x79
      13'h104C: dout  = 8'b01111001; // 4172 : 121 - 0x79
      13'h104D: dout  = 8'b01001001; // 4173 :  73 - 0x49
      13'h104E: dout  = 8'b01001111; // 4174 :  79 - 0x4f
      13'h104F: dout  = 8'b01001110; // 4175 :  78 - 0x4e
      13'h1050: dout  = 8'b11000111; // 4176 : 199 - 0xc7 -- Background 0x5
      13'h1051: dout  = 8'b11001111; // 4177 : 207 - 0xcf
      13'h1052: dout  = 8'b11011111; // 4178 : 223 - 0xdf
      13'h1053: dout  = 8'b11011111; // 4179 : 223 - 0xdf
      13'h1054: dout  = 8'b11001110; // 4180 : 206 - 0xce
      13'h1055: dout  = 8'b11100000; // 4181 : 224 - 0xe0
      13'h1056: dout  = 8'b11111111; // 4182 : 255 - 0xff
      13'h1057: dout  = 8'b11111111; // 4183 : 255 - 0xff
      13'h1058: dout  = 8'b01111000; // 4184 : 120 - 0x78
      13'h1059: dout  = 8'b01110000; // 4185 : 112 - 0x70
      13'h105A: dout  = 8'b01100000; // 4186 :  96 - 0x60
      13'h105B: dout  = 8'b01100000; // 4187 :  96 - 0x60
      13'h105C: dout  = 8'b01110001; // 4188 : 113 - 0x71
      13'h105D: dout  = 8'b01011111; // 4189 :  95 - 0x5f
      13'h105E: dout  = 8'b01111111; // 4190 : 127 - 0x7f
      13'h105F: dout  = 8'b00000000; // 4191 :   0 - 0x0
      13'h1060: dout  = 8'b11111111; // 4192 : 255 - 0xff -- Background 0x6
      13'h1061: dout  = 8'b11111111; // 4193 : 255 - 0xff
      13'h1062: dout  = 8'b00000111; // 4194 :   7 - 0x7
      13'h1063: dout  = 8'b01100011; // 4195 :  99 - 0x63
      13'h1064: dout  = 8'b01100011; // 4196 :  99 - 0x63
      13'h1065: dout  = 8'b01101111; // 4197 : 111 - 0x6f
      13'h1066: dout  = 8'b00001111; // 4198 :  15 - 0xf
      13'h1067: dout  = 8'b10001111; // 4199 : 143 - 0x8f
      13'h1068: dout  = 8'b00000000; // 4200 :   0 - 0x0
      13'h1069: dout  = 8'b11111110; // 4201 : 254 - 0xfe
      13'h106A: dout  = 8'b11111010; // 4202 : 250 - 0xfa
      13'h106B: dout  = 8'b10011110; // 4203 : 158 - 0x9e
      13'h106C: dout  = 8'b10011110; // 4204 : 158 - 0x9e
      13'h106D: dout  = 8'b10010010; // 4205 : 146 - 0x92
      13'h106E: dout  = 8'b11110010; // 4206 : 242 - 0xf2
      13'h106F: dout  = 8'b01110010; // 4207 : 114 - 0x72
      13'h1070: dout  = 8'b11100011; // 4208 : 227 - 0xe3 -- Background 0x7
      13'h1071: dout  = 8'b11110011; // 4209 : 243 - 0xf3
      13'h1072: dout  = 8'b11111011; // 4210 : 251 - 0xfb
      13'h1073: dout  = 8'b11111011; // 4211 : 251 - 0xfb
      13'h1074: dout  = 8'b01110011; // 4212 : 115 - 0x73
      13'h1075: dout  = 8'b00000111; // 4213 :   7 - 0x7
      13'h1076: dout  = 8'b11111111; // 4214 : 255 - 0xff
      13'h1077: dout  = 8'b11111111; // 4215 : 255 - 0xff
      13'h1078: dout  = 8'b00011110; // 4216 :  30 - 0x1e
      13'h1079: dout  = 8'b00001110; // 4217 :  14 - 0xe
      13'h107A: dout  = 8'b00000110; // 4218 :   6 - 0x6
      13'h107B: dout  = 8'b00000110; // 4219 :   6 - 0x6
      13'h107C: dout  = 8'b10001110; // 4220 : 142 - 0x8e
      13'h107D: dout  = 8'b11111010; // 4221 : 250 - 0xfa
      13'h107E: dout  = 8'b11111110; // 4222 : 254 - 0xfe
      13'h107F: dout  = 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout  = 8'b11111111; // 4224 : 255 - 0xff -- Background 0x8
      13'h1081: dout  = 8'b11010101; // 4225 : 213 - 0xd5
      13'h1082: dout  = 8'b10101010; // 4226 : 170 - 0xaa
      13'h1083: dout  = 8'b11010101; // 4227 : 213 - 0xd5
      13'h1084: dout  = 8'b10101010; // 4228 : 170 - 0xaa
      13'h1085: dout  = 8'b11010101; // 4229 : 213 - 0xd5
      13'h1086: dout  = 8'b10101010; // 4230 : 170 - 0xaa
      13'h1087: dout  = 8'b11010101; // 4231 : 213 - 0xd5
      13'h1088: dout  = 8'b00000000; // 4232 :   0 - 0x0
      13'h1089: dout  = 8'b01111111; // 4233 : 127 - 0x7f
      13'h108A: dout  = 8'b01011111; // 4234 :  95 - 0x5f
      13'h108B: dout  = 8'b01111111; // 4235 : 127 - 0x7f
      13'h108C: dout  = 8'b01111111; // 4236 : 127 - 0x7f
      13'h108D: dout  = 8'b01111111; // 4237 : 127 - 0x7f
      13'h108E: dout  = 8'b01111111; // 4238 : 127 - 0x7f
      13'h108F: dout  = 8'b01111111; // 4239 : 127 - 0x7f
      13'h1090: dout  = 8'b10101010; // 4240 : 170 - 0xaa -- Background 0x9
      13'h1091: dout  = 8'b11010101; // 4241 : 213 - 0xd5
      13'h1092: dout  = 8'b10101010; // 4242 : 170 - 0xaa
      13'h1093: dout  = 8'b11010101; // 4243 : 213 - 0xd5
      13'h1094: dout  = 8'b10101010; // 4244 : 170 - 0xaa
      13'h1095: dout  = 8'b11110101; // 4245 : 245 - 0xf5
      13'h1096: dout  = 8'b10101010; // 4246 : 170 - 0xaa
      13'h1097: dout  = 8'b11111111; // 4247 : 255 - 0xff
      13'h1098: dout  = 8'b01111111; // 4248 : 127 - 0x7f
      13'h1099: dout  = 8'b01111111; // 4249 : 127 - 0x7f
      13'h109A: dout  = 8'b01111111; // 4250 : 127 - 0x7f
      13'h109B: dout  = 8'b01111111; // 4251 : 127 - 0x7f
      13'h109C: dout  = 8'b01111111; // 4252 : 127 - 0x7f
      13'h109D: dout  = 8'b01011111; // 4253 :  95 - 0x5f
      13'h109E: dout  = 8'b01111111; // 4254 : 127 - 0x7f
      13'h109F: dout  = 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout  = 8'b11111111; // 4256 : 255 - 0xff -- Background 0xa
      13'h10A1: dout  = 8'b01010101; // 4257 :  85 - 0x55
      13'h10A2: dout  = 8'b10101111; // 4258 : 175 - 0xaf
      13'h10A3: dout  = 8'b01010101; // 4259 :  85 - 0x55
      13'h10A4: dout  = 8'b10101011; // 4260 : 171 - 0xab
      13'h10A5: dout  = 8'b01010101; // 4261 :  85 - 0x55
      13'h10A6: dout  = 8'b10101011; // 4262 : 171 - 0xab
      13'h10A7: dout  = 8'b01010101; // 4263 :  85 - 0x55
      13'h10A8: dout  = 8'b00000000; // 4264 :   0 - 0x0
      13'h10A9: dout  = 8'b11111110; // 4265 : 254 - 0xfe
      13'h10AA: dout  = 8'b11111010; // 4266 : 250 - 0xfa
      13'h10AB: dout  = 8'b11111110; // 4267 : 254 - 0xfe
      13'h10AC: dout  = 8'b11111110; // 4268 : 254 - 0xfe
      13'h10AD: dout  = 8'b11111110; // 4269 : 254 - 0xfe
      13'h10AE: dout  = 8'b11111110; // 4270 : 254 - 0xfe
      13'h10AF: dout  = 8'b11111110; // 4271 : 254 - 0xfe
      13'h10B0: dout  = 8'b10101011; // 4272 : 171 - 0xab -- Background 0xb
      13'h10B1: dout  = 8'b01010101; // 4273 :  85 - 0x55
      13'h10B2: dout  = 8'b10101011; // 4274 : 171 - 0xab
      13'h10B3: dout  = 8'b01010101; // 4275 :  85 - 0x55
      13'h10B4: dout  = 8'b10101011; // 4276 : 171 - 0xab
      13'h10B5: dout  = 8'b01010101; // 4277 :  85 - 0x55
      13'h10B6: dout  = 8'b10101011; // 4278 : 171 - 0xab
      13'h10B7: dout  = 8'b11111111; // 4279 : 255 - 0xff
      13'h10B8: dout  = 8'b11111110; // 4280 : 254 - 0xfe
      13'h10B9: dout  = 8'b11111110; // 4281 : 254 - 0xfe
      13'h10BA: dout  = 8'b11111110; // 4282 : 254 - 0xfe
      13'h10BB: dout  = 8'b11111110; // 4283 : 254 - 0xfe
      13'h10BC: dout  = 8'b11111110; // 4284 : 254 - 0xfe
      13'h10BD: dout  = 8'b11111010; // 4285 : 250 - 0xfa
      13'h10BE: dout  = 8'b11111110; // 4286 : 254 - 0xfe
      13'h10BF: dout  = 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout  = 8'b11111111; // 4288 : 255 - 0xff -- Background 0xc
      13'h10C1: dout  = 8'b11010101; // 4289 : 213 - 0xd5
      13'h10C2: dout  = 8'b10100000; // 4290 : 160 - 0xa0
      13'h10C3: dout  = 8'b11010000; // 4291 : 208 - 0xd0
      13'h10C4: dout  = 8'b10001111; // 4292 : 143 - 0x8f
      13'h10C5: dout  = 8'b11001000; // 4293 : 200 - 0xc8
      13'h10C6: dout  = 8'b10001000; // 4294 : 136 - 0x88
      13'h10C7: dout  = 8'b11001000; // 4295 : 200 - 0xc8
      13'h10C8: dout  = 8'b00000000; // 4296 :   0 - 0x0
      13'h10C9: dout  = 8'b00111111; // 4297 :  63 - 0x3f
      13'h10CA: dout  = 8'b01011111; // 4298 :  95 - 0x5f
      13'h10CB: dout  = 8'b01101111; // 4299 : 111 - 0x6f
      13'h10CC: dout  = 8'b01110000; // 4300 : 112 - 0x70
      13'h10CD: dout  = 8'b01110111; // 4301 : 119 - 0x77
      13'h10CE: dout  = 8'b01110111; // 4302 : 119 - 0x77
      13'h10CF: dout  = 8'b01110111; // 4303 : 119 - 0x77
      13'h10D0: dout  = 8'b10001000; // 4304 : 136 - 0x88 -- Background 0xd
      13'h10D1: dout  = 8'b11001000; // 4305 : 200 - 0xc8
      13'h10D2: dout  = 8'b10001000; // 4306 : 136 - 0x88
      13'h10D3: dout  = 8'b11001111; // 4307 : 207 - 0xcf
      13'h10D4: dout  = 8'b10010000; // 4308 : 144 - 0x90
      13'h10D5: dout  = 8'b11100000; // 4309 : 224 - 0xe0
      13'h10D6: dout  = 8'b11101010; // 4310 : 234 - 0xea
      13'h10D7: dout  = 8'b11111111; // 4311 : 255 - 0xff
      13'h10D8: dout  = 8'b01110111; // 4312 : 119 - 0x77
      13'h10D9: dout  = 8'b01110111; // 4313 : 119 - 0x77
      13'h10DA: dout  = 8'b01110111; // 4314 : 119 - 0x77
      13'h10DB: dout  = 8'b01110000; // 4315 : 112 - 0x70
      13'h10DC: dout  = 8'b01101111; // 4316 : 111 - 0x6f
      13'h10DD: dout  = 8'b01011111; // 4317 :  95 - 0x5f
      13'h10DE: dout  = 8'b00010101; // 4318 :  21 - 0x15
      13'h10DF: dout  = 8'b00000000; // 4319 :   0 - 0x0
      13'h10E0: dout  = 8'b11111111; // 4320 : 255 - 0xff -- Background 0xe
      13'h10E1: dout  = 8'b01011011; // 4321 :  91 - 0x5b
      13'h10E2: dout  = 8'b00000111; // 4322 :   7 - 0x7
      13'h10E3: dout  = 8'b00001001; // 4323 :   9 - 0x9
      13'h10E4: dout  = 8'b11110011; // 4324 : 243 - 0xf3
      13'h10E5: dout  = 8'b00010001; // 4325 :  17 - 0x11
      13'h10E6: dout  = 8'b00010011; // 4326 :  19 - 0x13
      13'h10E7: dout  = 8'b00010001; // 4327 :  17 - 0x11
      13'h10E8: dout  = 8'b00000000; // 4328 :   0 - 0x0
      13'h10E9: dout  = 8'b11111100; // 4329 : 252 - 0xfc
      13'h10EA: dout  = 8'b11111000; // 4330 : 248 - 0xf8
      13'h10EB: dout  = 8'b11110110; // 4331 : 246 - 0xf6
      13'h10EC: dout  = 8'b00001100; // 4332 :  12 - 0xc
      13'h10ED: dout  = 8'b11101110; // 4333 : 238 - 0xee
      13'h10EE: dout  = 8'b11101100; // 4334 : 236 - 0xec
      13'h10EF: dout  = 8'b11101110; // 4335 : 238 - 0xee
      13'h10F0: dout  = 8'b00010011; // 4336 :  19 - 0x13 -- Background 0xf
      13'h10F1: dout  = 8'b00010001; // 4337 :  17 - 0x11
      13'h10F2: dout  = 8'b00010011; // 4338 :  19 - 0x13
      13'h10F3: dout  = 8'b11110001; // 4339 : 241 - 0xf1
      13'h10F4: dout  = 8'b00001011; // 4340 :  11 - 0xb
      13'h10F5: dout  = 8'b00000101; // 4341 :   5 - 0x5
      13'h10F6: dout  = 8'b10101011; // 4342 : 171 - 0xab
      13'h10F7: dout  = 8'b11111111; // 4343 : 255 - 0xff
      13'h10F8: dout  = 8'b11101100; // 4344 : 236 - 0xec
      13'h10F9: dout  = 8'b11101110; // 4345 : 238 - 0xee
      13'h10FA: dout  = 8'b11101100; // 4346 : 236 - 0xec
      13'h10FB: dout  = 8'b00001110; // 4347 :  14 - 0xe
      13'h10FC: dout  = 8'b11110100; // 4348 : 244 - 0xf4
      13'h10FD: dout  = 8'b11111010; // 4349 : 250 - 0xfa
      13'h10FE: dout  = 8'b01010100; // 4350 :  84 - 0x54
      13'h10FF: dout  = 8'b00000000; // 4351 :   0 - 0x0
      13'h1100: dout  = 8'b11010000; // 4352 : 208 - 0xd0 -- Background 0x10
      13'h1101: dout  = 8'b10010000; // 4353 : 144 - 0x90
      13'h1102: dout  = 8'b11011111; // 4354 : 223 - 0xdf
      13'h1103: dout  = 8'b10011010; // 4355 : 154 - 0x9a
      13'h1104: dout  = 8'b11010101; // 4356 : 213 - 0xd5
      13'h1105: dout  = 8'b10011111; // 4357 : 159 - 0x9f
      13'h1106: dout  = 8'b11010000; // 4358 : 208 - 0xd0
      13'h1107: dout  = 8'b10010000; // 4359 : 144 - 0x90
      13'h1108: dout  = 8'b01100000; // 4360 :  96 - 0x60
      13'h1109: dout  = 8'b01100000; // 4361 :  96 - 0x60
      13'h110A: dout  = 8'b01100000; // 4362 :  96 - 0x60
      13'h110B: dout  = 8'b01101111; // 4363 : 111 - 0x6f
      13'h110C: dout  = 8'b01101010; // 4364 : 106 - 0x6a
      13'h110D: dout  = 8'b01100000; // 4365 :  96 - 0x60
      13'h110E: dout  = 8'b01100000; // 4366 :  96 - 0x60
      13'h110F: dout  = 8'b01100000; // 4367 :  96 - 0x60
      13'h1110: dout  = 8'b00001001; // 4368 :   9 - 0x9 -- Background 0x11
      13'h1111: dout  = 8'b00001011; // 4369 :  11 - 0xb
      13'h1112: dout  = 8'b11111001; // 4370 : 249 - 0xf9
      13'h1113: dout  = 8'b10101011; // 4371 : 171 - 0xab
      13'h1114: dout  = 8'b01011001; // 4372 :  89 - 0x59
      13'h1115: dout  = 8'b11111011; // 4373 : 251 - 0xfb
      13'h1116: dout  = 8'b00001001; // 4374 :   9 - 0x9
      13'h1117: dout  = 8'b00001011; // 4375 :  11 - 0xb
      13'h1118: dout  = 8'b00000110; // 4376 :   6 - 0x6
      13'h1119: dout  = 8'b00000100; // 4377 :   4 - 0x4
      13'h111A: dout  = 8'b00000110; // 4378 :   6 - 0x6
      13'h111B: dout  = 8'b11110100; // 4379 : 244 - 0xf4
      13'h111C: dout  = 8'b10100110; // 4380 : 166 - 0xa6
      13'h111D: dout  = 8'b00000100; // 4381 :   4 - 0x4
      13'h111E: dout  = 8'b00000110; // 4382 :   6 - 0x6
      13'h111F: dout  = 8'b00000100; // 4383 :   4 - 0x4
      13'h1120: dout  = 8'b00011000; // 4384 :  24 - 0x18 -- Background 0x12
      13'h1121: dout  = 8'b00010100; // 4385 :  20 - 0x14
      13'h1122: dout  = 8'b00010100; // 4386 :  20 - 0x14
      13'h1123: dout  = 8'b00111010; // 4387 :  58 - 0x3a
      13'h1124: dout  = 8'b00111010; // 4388 :  58 - 0x3a
      13'h1125: dout  = 8'b01111010; // 4389 : 122 - 0x7a
      13'h1126: dout  = 8'b01111010; // 4390 : 122 - 0x7a
      13'h1127: dout  = 8'b01111010; // 4391 : 122 - 0x7a
      13'h1128: dout  = 8'b00000000; // 4392 :   0 - 0x0
      13'h1129: dout  = 8'b00001000; // 4393 :   8 - 0x8
      13'h112A: dout  = 8'b00001000; // 4394 :   8 - 0x8
      13'h112B: dout  = 8'b00011100; // 4395 :  28 - 0x1c
      13'h112C: dout  = 8'b00011100; // 4396 :  28 - 0x1c
      13'h112D: dout  = 8'b00111100; // 4397 :  60 - 0x3c
      13'h112E: dout  = 8'b00111100; // 4398 :  60 - 0x3c
      13'h112F: dout  = 8'b00111100; // 4399 :  60 - 0x3c
      13'h1130: dout  = 8'b11111011; // 4400 : 251 - 0xfb -- Background 0x13
      13'h1131: dout  = 8'b11111101; // 4401 : 253 - 0xfd
      13'h1132: dout  = 8'b11111101; // 4402 : 253 - 0xfd
      13'h1133: dout  = 8'b11111101; // 4403 : 253 - 0xfd
      13'h1134: dout  = 8'b11111101; // 4404 : 253 - 0xfd
      13'h1135: dout  = 8'b11111101; // 4405 : 253 - 0xfd
      13'h1136: dout  = 8'b10000001; // 4406 : 129 - 0x81
      13'h1137: dout  = 8'b11111111; // 4407 : 255 - 0xff
      13'h1138: dout  = 8'b00111100; // 4408 :  60 - 0x3c
      13'h1139: dout  = 8'b01111110; // 4409 : 126 - 0x7e
      13'h113A: dout  = 8'b01111110; // 4410 : 126 - 0x7e
      13'h113B: dout  = 8'b01111110; // 4411 : 126 - 0x7e
      13'h113C: dout  = 8'b01111110; // 4412 : 126 - 0x7e
      13'h113D: dout  = 8'b01111110; // 4413 : 126 - 0x7e
      13'h113E: dout  = 8'b01111110; // 4414 : 126 - 0x7e
      13'h113F: dout  = 8'b00000000; // 4415 :   0 - 0x0
      13'h1140: dout  = 8'b00000000; // 4416 :   0 - 0x0 -- Background 0x14
      13'h1141: dout  = 8'b00000111; // 4417 :   7 - 0x7
      13'h1142: dout  = 8'b00000010; // 4418 :   2 - 0x2
      13'h1143: dout  = 8'b00000100; // 4419 :   4 - 0x4
      13'h1144: dout  = 8'b00000011; // 4420 :   3 - 0x3
      13'h1145: dout  = 8'b00000011; // 4421 :   3 - 0x3
      13'h1146: dout  = 8'b00001101; // 4422 :  13 - 0xd
      13'h1147: dout  = 8'b00010111; // 4423 :  23 - 0x17
      13'h1148: dout  = 8'b00000000; // 4424 :   0 - 0x0
      13'h1149: dout  = 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout  = 8'b00000101; // 4426 :   5 - 0x5
      13'h114B: dout  = 8'b00000011; // 4427 :   3 - 0x3
      13'h114C: dout  = 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout  = 8'b00000000; // 4429 :   0 - 0x0
      13'h114E: dout  = 8'b00000010; // 4430 :   2 - 0x2
      13'h114F: dout  = 8'b00001111; // 4431 :  15 - 0xf
      13'h1150: dout  = 8'b00101111; // 4432 :  47 - 0x2f -- Background 0x15
      13'h1151: dout  = 8'b01001111; // 4433 :  79 - 0x4f
      13'h1152: dout  = 8'b01001111; // 4434 :  79 - 0x4f
      13'h1153: dout  = 8'b01001111; // 4435 :  79 - 0x4f
      13'h1154: dout  = 8'b01001111; // 4436 :  79 - 0x4f
      13'h1155: dout  = 8'b00100111; // 4437 :  39 - 0x27
      13'h1156: dout  = 8'b00010000; // 4438 :  16 - 0x10
      13'h1157: dout  = 8'b00001111; // 4439 :  15 - 0xf
      13'h1158: dout  = 8'b00011100; // 4440 :  28 - 0x1c
      13'h1159: dout  = 8'b00111010; // 4441 :  58 - 0x3a
      13'h115A: dout  = 8'b00111100; // 4442 :  60 - 0x3c
      13'h115B: dout  = 8'b00111111; // 4443 :  63 - 0x3f
      13'h115C: dout  = 8'b00111000; // 4444 :  56 - 0x38
      13'h115D: dout  = 8'b00011110; // 4445 :  30 - 0x1e
      13'h115E: dout  = 8'b00001111; // 4446 :  15 - 0xf
      13'h115F: dout  = 8'b00000000; // 4447 :   0 - 0x0
      13'h1160: dout  = 8'b00000000; // 4448 :   0 - 0x0 -- Background 0x16
      13'h1161: dout  = 8'b11100000; // 4449 : 224 - 0xe0
      13'h1162: dout  = 8'b10100000; // 4450 : 160 - 0xa0
      13'h1163: dout  = 8'b00100000; // 4451 :  32 - 0x20
      13'h1164: dout  = 8'b11000000; // 4452 : 192 - 0xc0
      13'h1165: dout  = 8'b01000000; // 4453 :  64 - 0x40
      13'h1166: dout  = 8'b00110000; // 4454 :  48 - 0x30
      13'h1167: dout  = 8'b11101000; // 4455 : 232 - 0xe8
      13'h1168: dout  = 8'b00000000; // 4456 :   0 - 0x0
      13'h1169: dout  = 8'b00000000; // 4457 :   0 - 0x0
      13'h116A: dout  = 8'b01000000; // 4458 :  64 - 0x40
      13'h116B: dout  = 8'b11000000; // 4459 : 192 - 0xc0
      13'h116C: dout  = 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout  = 8'b10000000; // 4461 : 128 - 0x80
      13'h116E: dout  = 8'b11000000; // 4462 : 192 - 0xc0
      13'h116F: dout  = 8'b01110000; // 4463 : 112 - 0x70
      13'h1170: dout  = 8'b11110100; // 4464 : 244 - 0xf4 -- Background 0x17
      13'h1171: dout  = 8'b11110010; // 4465 : 242 - 0xf2
      13'h1172: dout  = 8'b11110010; // 4466 : 242 - 0xf2
      13'h1173: dout  = 8'b11110010; // 4467 : 242 - 0xf2
      13'h1174: dout  = 8'b11110010; // 4468 : 242 - 0xf2
      13'h1175: dout  = 8'b11100100; // 4469 : 228 - 0xe4
      13'h1176: dout  = 8'b00001000; // 4470 :   8 - 0x8
      13'h1177: dout  = 8'b11110000; // 4471 : 240 - 0xf0
      13'h1178: dout  = 8'b00011000; // 4472 :  24 - 0x18
      13'h1179: dout  = 8'b11111100; // 4473 : 252 - 0xfc
      13'h117A: dout  = 8'b00111100; // 4474 :  60 - 0x3c
      13'h117B: dout  = 8'b01011100; // 4475 :  92 - 0x5c
      13'h117C: dout  = 8'b00111100; // 4476 :  60 - 0x3c
      13'h117D: dout  = 8'b11111000; // 4477 : 248 - 0xf8
      13'h117E: dout  = 8'b11110000; // 4478 : 240 - 0xf0
      13'h117F: dout  = 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout  = 8'b00111111; // 4480 :  63 - 0x3f -- Background 0x18
      13'h1181: dout  = 8'b01000000; // 4481 :  64 - 0x40
      13'h1182: dout  = 8'b01000000; // 4482 :  64 - 0x40
      13'h1183: dout  = 8'b10000000; // 4483 : 128 - 0x80
      13'h1184: dout  = 8'b10000000; // 4484 : 128 - 0x80
      13'h1185: dout  = 8'b01111111; // 4485 : 127 - 0x7f
      13'h1186: dout  = 8'b00000001; // 4486 :   1 - 0x1
      13'h1187: dout  = 8'b01111111; // 4487 : 127 - 0x7f
      13'h1188: dout  = 8'b00000000; // 4488 :   0 - 0x0
      13'h1189: dout  = 8'b00111111; // 4489 :  63 - 0x3f
      13'h118A: dout  = 8'b00111111; // 4490 :  63 - 0x3f
      13'h118B: dout  = 8'b01111111; // 4491 : 127 - 0x7f
      13'h118C: dout  = 8'b01111111; // 4492 : 127 - 0x7f
      13'h118D: dout  = 8'b00000000; // 4493 :   0 - 0x0
      13'h118E: dout  = 8'b00000000; // 4494 :   0 - 0x0
      13'h118F: dout  = 8'b00000000; // 4495 :   0 - 0x0
      13'h1190: dout  = 8'b11111100; // 4496 : 252 - 0xfc -- Background 0x19
      13'h1191: dout  = 8'b00000010; // 4497 :   2 - 0x2
      13'h1192: dout  = 8'b00000010; // 4498 :   2 - 0x2
      13'h1193: dout  = 8'b00000001; // 4499 :   1 - 0x1
      13'h1194: dout  = 8'b00000001; // 4500 :   1 - 0x1
      13'h1195: dout  = 8'b11111110; // 4501 : 254 - 0xfe
      13'h1196: dout  = 8'b10000000; // 4502 : 128 - 0x80
      13'h1197: dout  = 8'b11111110; // 4503 : 254 - 0xfe
      13'h1198: dout  = 8'b00000000; // 4504 :   0 - 0x0
      13'h1199: dout  = 8'b11111100; // 4505 : 252 - 0xfc
      13'h119A: dout  = 8'b11111100; // 4506 : 252 - 0xfc
      13'h119B: dout  = 8'b11111110; // 4507 : 254 - 0xfe
      13'h119C: dout  = 8'b11111110; // 4508 : 254 - 0xfe
      13'h119D: dout  = 8'b00000000; // 4509 :   0 - 0x0
      13'h119E: dout  = 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout  = 8'b00000000; // 4511 :   0 - 0x0
      13'h11A0: dout  = 8'b00000000; // 4512 :   0 - 0x0 -- Background 0x1a
      13'h11A1: dout  = 8'b00000000; // 4513 :   0 - 0x0
      13'h11A2: dout  = 8'b00111111; // 4514 :  63 - 0x3f
      13'h11A3: dout  = 8'b01000000; // 4515 :  64 - 0x40
      13'h11A4: dout  = 8'b01000000; // 4516 :  64 - 0x40
      13'h11A5: dout  = 8'b10000000; // 4517 : 128 - 0x80
      13'h11A6: dout  = 8'b10000000; // 4518 : 128 - 0x80
      13'h11A7: dout  = 8'b01111111; // 4519 : 127 - 0x7f
      13'h11A8: dout  = 8'b00000000; // 4520 :   0 - 0x0
      13'h11A9: dout  = 8'b00000000; // 4521 :   0 - 0x0
      13'h11AA: dout  = 8'b00000000; // 4522 :   0 - 0x0
      13'h11AB: dout  = 8'b00111111; // 4523 :  63 - 0x3f
      13'h11AC: dout  = 8'b00111111; // 4524 :  63 - 0x3f
      13'h11AD: dout  = 8'b01111111; // 4525 : 127 - 0x7f
      13'h11AE: dout  = 8'b01111111; // 4526 : 127 - 0x7f
      13'h11AF: dout  = 8'b00000000; // 4527 :   0 - 0x0
      13'h11B0: dout  = 8'b00000000; // 4528 :   0 - 0x0 -- Background 0x1b
      13'h11B1: dout  = 8'b00000000; // 4529 :   0 - 0x0
      13'h11B2: dout  = 8'b11111100; // 4530 : 252 - 0xfc
      13'h11B3: dout  = 8'b00000010; // 4531 :   2 - 0x2
      13'h11B4: dout  = 8'b00000010; // 4532 :   2 - 0x2
      13'h11B5: dout  = 8'b00000001; // 4533 :   1 - 0x1
      13'h11B6: dout  = 8'b00000001; // 4534 :   1 - 0x1
      13'h11B7: dout  = 8'b11111110; // 4535 : 254 - 0xfe
      13'h11B8: dout  = 8'b00000000; // 4536 :   0 - 0x0
      13'h11B9: dout  = 8'b00000000; // 4537 :   0 - 0x0
      13'h11BA: dout  = 8'b00000000; // 4538 :   0 - 0x0
      13'h11BB: dout  = 8'b11111100; // 4539 : 252 - 0xfc
      13'h11BC: dout  = 8'b11111100; // 4540 : 252 - 0xfc
      13'h11BD: dout  = 8'b11111110; // 4541 : 254 - 0xfe
      13'h11BE: dout  = 8'b11111110; // 4542 : 254 - 0xfe
      13'h11BF: dout  = 8'b00000000; // 4543 :   0 - 0x0
      13'h11C0: dout  = 8'b01111111; // 4544 : 127 - 0x7f -- Background 0x1c
      13'h11C1: dout  = 8'b10000000; // 4545 : 128 - 0x80
      13'h11C2: dout  = 8'b10000000; // 4546 : 128 - 0x80
      13'h11C3: dout  = 8'b10000000; // 4547 : 128 - 0x80
      13'h11C4: dout  = 8'b10011011; // 4548 : 155 - 0x9b
      13'h11C5: dout  = 8'b10100100; // 4549 : 164 - 0xa4
      13'h11C6: dout  = 8'b10100110; // 4550 : 166 - 0xa6
      13'h11C7: dout  = 8'b10000000; // 4551 : 128 - 0x80
      13'h11C8: dout  = 8'b00000000; // 4552 :   0 - 0x0
      13'h11C9: dout  = 8'b01111111; // 4553 : 127 - 0x7f
      13'h11CA: dout  = 8'b01111111; // 4554 : 127 - 0x7f
      13'h11CB: dout  = 8'b01111111; // 4555 : 127 - 0x7f
      13'h11CC: dout  = 8'b01100100; // 4556 : 100 - 0x64
      13'h11CD: dout  = 8'b01011011; // 4557 :  91 - 0x5b
      13'h11CE: dout  = 8'b01011001; // 4558 :  89 - 0x59
      13'h11CF: dout  = 8'b01111111; // 4559 : 127 - 0x7f
      13'h11D0: dout  = 8'b10000000; // 4560 : 128 - 0x80 -- Background 0x1d
      13'h11D1: dout  = 8'b01111111; // 4561 : 127 - 0x7f
      13'h11D2: dout  = 8'b00000010; // 4562 :   2 - 0x2
      13'h11D3: dout  = 8'b00000010; // 4563 :   2 - 0x2
      13'h11D4: dout  = 8'b00000010; // 4564 :   2 - 0x2
      13'h11D5: dout  = 8'b00000010; // 4565 :   2 - 0x2
      13'h11D6: dout  = 8'b00000010; // 4566 :   2 - 0x2
      13'h11D7: dout  = 8'b00001111; // 4567 :  15 - 0xf
      13'h11D8: dout  = 8'b01111111; // 4568 : 127 - 0x7f
      13'h11D9: dout  = 8'b00000000; // 4569 :   0 - 0x0
      13'h11DA: dout  = 8'b00000001; // 4570 :   1 - 0x1
      13'h11DB: dout  = 8'b00000001; // 4571 :   1 - 0x1
      13'h11DC: dout  = 8'b00000001; // 4572 :   1 - 0x1
      13'h11DD: dout  = 8'b00000001; // 4573 :   1 - 0x1
      13'h11DE: dout  = 8'b00000001; // 4574 :   1 - 0x1
      13'h11DF: dout  = 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout  = 8'b11111110; // 4576 : 254 - 0xfe -- Background 0x1e
      13'h11E1: dout  = 8'b00000001; // 4577 :   1 - 0x1
      13'h11E2: dout  = 8'b00000001; // 4578 :   1 - 0x1
      13'h11E3: dout  = 8'b00000001; // 4579 :   1 - 0x1
      13'h11E4: dout  = 8'b01000001; // 4580 :  65 - 0x41
      13'h11E5: dout  = 8'b11110101; // 4581 : 245 - 0xf5
      13'h11E6: dout  = 8'b00011101; // 4582 :  29 - 0x1d
      13'h11E7: dout  = 8'b00000001; // 4583 :   1 - 0x1
      13'h11E8: dout  = 8'b00000000; // 4584 :   0 - 0x0
      13'h11E9: dout  = 8'b11111110; // 4585 : 254 - 0xfe
      13'h11EA: dout  = 8'b11111110; // 4586 : 254 - 0xfe
      13'h11EB: dout  = 8'b11111110; // 4587 : 254 - 0xfe
      13'h11EC: dout  = 8'b10111110; // 4588 : 190 - 0xbe
      13'h11ED: dout  = 8'b00001010; // 4589 :  10 - 0xa
      13'h11EE: dout  = 8'b11100010; // 4590 : 226 - 0xe2
      13'h11EF: dout  = 8'b11111110; // 4591 : 254 - 0xfe
      13'h11F0: dout  = 8'b00000001; // 4592 :   1 - 0x1 -- Background 0x1f
      13'h11F1: dout  = 8'b11111110; // 4593 : 254 - 0xfe
      13'h11F2: dout  = 8'b01000000; // 4594 :  64 - 0x40
      13'h11F3: dout  = 8'b01000000; // 4595 :  64 - 0x40
      13'h11F4: dout  = 8'b01000000; // 4596 :  64 - 0x40
      13'h11F5: dout  = 8'b01000000; // 4597 :  64 - 0x40
      13'h11F6: dout  = 8'b01000000; // 4598 :  64 - 0x40
      13'h11F7: dout  = 8'b11110000; // 4599 : 240 - 0xf0
      13'h11F8: dout  = 8'b11111110; // 4600 : 254 - 0xfe
      13'h11F9: dout  = 8'b00000000; // 4601 :   0 - 0x0
      13'h11FA: dout  = 8'b10000000; // 4602 : 128 - 0x80
      13'h11FB: dout  = 8'b10000000; // 4603 : 128 - 0x80
      13'h11FC: dout  = 8'b10000000; // 4604 : 128 - 0x80
      13'h11FD: dout  = 8'b10000000; // 4605 : 128 - 0x80
      13'h11FE: dout  = 8'b10000000; // 4606 : 128 - 0x80
      13'h11FF: dout  = 8'b00000000; // 4607 :   0 - 0x0
      13'h1200: dout  = 8'b00000111; // 4608 :   7 - 0x7 -- Background 0x20
      13'h1201: dout  = 8'b00011111; // 4609 :  31 - 0x1f
      13'h1202: dout  = 8'b00111111; // 4610 :  63 - 0x3f
      13'h1203: dout  = 8'b01111111; // 4611 : 127 - 0x7f
      13'h1204: dout  = 8'b01111111; // 4612 : 127 - 0x7f
      13'h1205: dout  = 8'b11111111; // 4613 : 255 - 0xff
      13'h1206: dout  = 8'b11111111; // 4614 : 255 - 0xff
      13'h1207: dout  = 8'b11111111; // 4615 : 255 - 0xff
      13'h1208: dout  = 8'b00000000; // 4616 :   0 - 0x0
      13'h1209: dout  = 8'b00000000; // 4617 :   0 - 0x0
      13'h120A: dout  = 8'b00000000; // 4618 :   0 - 0x0
      13'h120B: dout  = 8'b00000000; // 4619 :   0 - 0x0
      13'h120C: dout  = 8'b00000000; // 4620 :   0 - 0x0
      13'h120D: dout  = 8'b00000000; // 4621 :   0 - 0x0
      13'h120E: dout  = 8'b00000000; // 4622 :   0 - 0x0
      13'h120F: dout  = 8'b00000000; // 4623 :   0 - 0x0
      13'h1210: dout  = 8'b11100000; // 4624 : 224 - 0xe0 -- Background 0x21
      13'h1211: dout  = 8'b11111000; // 4625 : 248 - 0xf8
      13'h1212: dout  = 8'b11111100; // 4626 : 252 - 0xfc
      13'h1213: dout  = 8'b11111110; // 4627 : 254 - 0xfe
      13'h1214: dout  = 8'b11111110; // 4628 : 254 - 0xfe
      13'h1215: dout  = 8'b11111111; // 4629 : 255 - 0xff
      13'h1216: dout  = 8'b11111111; // 4630 : 255 - 0xff
      13'h1217: dout  = 8'b11111111; // 4631 : 255 - 0xff
      13'h1218: dout  = 8'b00000000; // 4632 :   0 - 0x0
      13'h1219: dout  = 8'b00000000; // 4633 :   0 - 0x0
      13'h121A: dout  = 8'b00000000; // 4634 :   0 - 0x0
      13'h121B: dout  = 8'b00000000; // 4635 :   0 - 0x0
      13'h121C: dout  = 8'b00000000; // 4636 :   0 - 0x0
      13'h121D: dout  = 8'b00000000; // 4637 :   0 - 0x0
      13'h121E: dout  = 8'b00000000; // 4638 :   0 - 0x0
      13'h121F: dout  = 8'b00000000; // 4639 :   0 - 0x0
      13'h1220: dout  = 8'b00000111; // 4640 :   7 - 0x7 -- Background 0x22
      13'h1221: dout  = 8'b00011111; // 4641 :  31 - 0x1f
      13'h1222: dout  = 8'b00111111; // 4642 :  63 - 0x3f
      13'h1223: dout  = 8'b01111111; // 4643 : 127 - 0x7f
      13'h1224: dout  = 8'b01111111; // 4644 : 127 - 0x7f
      13'h1225: dout  = 8'b11111111; // 4645 : 255 - 0xff
      13'h1226: dout  = 8'b11111111; // 4646 : 255 - 0xff
      13'h1227: dout  = 8'b11111111; // 4647 : 255 - 0xff
      13'h1228: dout  = 8'b00000000; // 4648 :   0 - 0x0
      13'h1229: dout  = 8'b00000000; // 4649 :   0 - 0x0
      13'h122A: dout  = 8'b00011000; // 4650 :  24 - 0x18
      13'h122B: dout  = 8'b00010000; // 4651 :  16 - 0x10
      13'h122C: dout  = 8'b00011010; // 4652 :  26 - 0x1a
      13'h122D: dout  = 8'b00010001; // 4653 :  17 - 0x11
      13'h122E: dout  = 8'b00011010; // 4654 :  26 - 0x1a
      13'h122F: dout  = 8'b00000000; // 4655 :   0 - 0x0
      13'h1230: dout  = 8'b11100000; // 4656 : 224 - 0xe0 -- Background 0x23
      13'h1231: dout  = 8'b11111000; // 4657 : 248 - 0xf8
      13'h1232: dout  = 8'b11111100; // 4658 : 252 - 0xfc
      13'h1233: dout  = 8'b11111110; // 4659 : 254 - 0xfe
      13'h1234: dout  = 8'b11111110; // 4660 : 254 - 0xfe
      13'h1235: dout  = 8'b11111111; // 4661 : 255 - 0xff
      13'h1236: dout  = 8'b11111111; // 4662 : 255 - 0xff
      13'h1237: dout  = 8'b11111111; // 4663 : 255 - 0xff
      13'h1238: dout  = 8'b00000000; // 4664 :   0 - 0x0
      13'h1239: dout  = 8'b00000000; // 4665 :   0 - 0x0
      13'h123A: dout  = 8'b00000000; // 4666 :   0 - 0x0
      13'h123B: dout  = 8'b00101000; // 4667 :  40 - 0x28
      13'h123C: dout  = 8'b10001100; // 4668 : 140 - 0x8c
      13'h123D: dout  = 8'b00101000; // 4669 :  40 - 0x28
      13'h123E: dout  = 8'b10101100; // 4670 : 172 - 0xac
      13'h123F: dout  = 8'b00000000; // 4671 :   0 - 0x0
      13'h1240: dout  = 8'b00000000; // 4672 :   0 - 0x0 -- Background 0x24
      13'h1241: dout  = 8'b00000000; // 4673 :   0 - 0x0
      13'h1242: dout  = 8'b00000000; // 4674 :   0 - 0x0
      13'h1243: dout  = 8'b00000000; // 4675 :   0 - 0x0
      13'h1244: dout  = 8'b00000000; // 4676 :   0 - 0x0
      13'h1245: dout  = 8'b00000000; // 4677 :   0 - 0x0
      13'h1246: dout  = 8'b00000000; // 4678 :   0 - 0x0
      13'h1247: dout  = 8'b00000000; // 4679 :   0 - 0x0
      13'h1248: dout  = 8'b00000000; // 4680 :   0 - 0x0
      13'h1249: dout  = 8'b00000000; // 4681 :   0 - 0x0
      13'h124A: dout  = 8'b00000000; // 4682 :   0 - 0x0
      13'h124B: dout  = 8'b00000000; // 4683 :   0 - 0x0
      13'h124C: dout  = 8'b00000000; // 4684 :   0 - 0x0
      13'h124D: dout  = 8'b00000000; // 4685 :   0 - 0x0
      13'h124E: dout  = 8'b00000000; // 4686 :   0 - 0x0
      13'h124F: dout  = 8'b00000000; // 4687 :   0 - 0x0
      13'h1250: dout  = 8'b00101111; // 4688 :  47 - 0x2f -- Background 0x25
      13'h1251: dout  = 8'b01001111; // 4689 :  79 - 0x4f
      13'h1252: dout  = 8'b01001111; // 4690 :  79 - 0x4f
      13'h1253: dout  = 8'b01001111; // 4691 :  79 - 0x4f
      13'h1254: dout  = 8'b01001111; // 4692 :  79 - 0x4f
      13'h1255: dout  = 8'b00100111; // 4693 :  39 - 0x27
      13'h1256: dout  = 8'b00010000; // 4694 :  16 - 0x10
      13'h1257: dout  = 8'b00001111; // 4695 :  15 - 0xf
      13'h1258: dout  = 8'b00011100; // 4696 :  28 - 0x1c
      13'h1259: dout  = 8'b00111001; // 4697 :  57 - 0x39
      13'h125A: dout  = 8'b00111111; // 4698 :  63 - 0x3f
      13'h125B: dout  = 8'b00111110; // 4699 :  62 - 0x3e
      13'h125C: dout  = 8'b00111111; // 4700 :  63 - 0x3f
      13'h125D: dout  = 8'b00011110; // 4701 :  30 - 0x1e
      13'h125E: dout  = 8'b00001111; // 4702 :  15 - 0xf
      13'h125F: dout  = 8'b00000000; // 4703 :   0 - 0x0
      13'h1260: dout  = 8'b00000000; // 4704 :   0 - 0x0 -- Background 0x26
      13'h1261: dout  = 8'b11100000; // 4705 : 224 - 0xe0
      13'h1262: dout  = 8'b10100000; // 4706 : 160 - 0xa0
      13'h1263: dout  = 8'b00100000; // 4707 :  32 - 0x20
      13'h1264: dout  = 8'b11000000; // 4708 : 192 - 0xc0
      13'h1265: dout  = 8'b01000000; // 4709 :  64 - 0x40
      13'h1266: dout  = 8'b00110000; // 4710 :  48 - 0x30
      13'h1267: dout  = 8'b11101000; // 4711 : 232 - 0xe8
      13'h1268: dout  = 8'b00000000; // 4712 :   0 - 0x0
      13'h1269: dout  = 8'b00000000; // 4713 :   0 - 0x0
      13'h126A: dout  = 8'b01000000; // 4714 :  64 - 0x40
      13'h126B: dout  = 8'b11000000; // 4715 : 192 - 0xc0
      13'h126C: dout  = 8'b00000000; // 4716 :   0 - 0x0
      13'h126D: dout  = 8'b10000000; // 4717 : 128 - 0x80
      13'h126E: dout  = 8'b11000000; // 4718 : 192 - 0xc0
      13'h126F: dout  = 8'b11110000; // 4719 : 240 - 0xf0
      13'h1270: dout  = 8'b11110100; // 4720 : 244 - 0xf4 -- Background 0x27
      13'h1271: dout  = 8'b11110010; // 4721 : 242 - 0xf2
      13'h1272: dout  = 8'b11110010; // 4722 : 242 - 0xf2
      13'h1273: dout  = 8'b11110010; // 4723 : 242 - 0xf2
      13'h1274: dout  = 8'b11110010; // 4724 : 242 - 0xf2
      13'h1275: dout  = 8'b11100100; // 4725 : 228 - 0xe4
      13'h1276: dout  = 8'b00001000; // 4726 :   8 - 0x8
      13'h1277: dout  = 8'b11110000; // 4727 : 240 - 0xf0
      13'h1278: dout  = 8'b00111000; // 4728 :  56 - 0x38
      13'h1279: dout  = 8'b10011100; // 4729 : 156 - 0x9c
      13'h127A: dout  = 8'b10011100; // 4730 : 156 - 0x9c
      13'h127B: dout  = 8'b00111100; // 4731 :  60 - 0x3c
      13'h127C: dout  = 8'b11111100; // 4732 : 252 - 0xfc
      13'h127D: dout  = 8'b01111000; // 4733 : 120 - 0x78
      13'h127E: dout  = 8'b11110000; // 4734 : 240 - 0xf0
      13'h127F: dout  = 8'b00000000; // 4735 :   0 - 0x0
      13'h1280: dout  = 8'b11111111; // 4736 : 255 - 0xff -- Background 0x28
      13'h1281: dout  = 8'b11010101; // 4737 : 213 - 0xd5
      13'h1282: dout  = 8'b10100011; // 4738 : 163 - 0xa3
      13'h1283: dout  = 8'b11010111; // 4739 : 215 - 0xd7
      13'h1284: dout  = 8'b10001111; // 4740 : 143 - 0x8f
      13'h1285: dout  = 8'b11001111; // 4741 : 207 - 0xcf
      13'h1286: dout  = 8'b10001011; // 4742 : 139 - 0x8b
      13'h1287: dout  = 8'b11001011; // 4743 : 203 - 0xcb
      13'h1288: dout  = 8'b00000000; // 4744 :   0 - 0x0
      13'h1289: dout  = 8'b00111110; // 4745 :  62 - 0x3e
      13'h128A: dout  = 8'b01011101; // 4746 :  93 - 0x5d
      13'h128B: dout  = 8'b01101011; // 4747 : 107 - 0x6b
      13'h128C: dout  = 8'b01110101; // 4748 : 117 - 0x75
      13'h128D: dout  = 8'b01110001; // 4749 : 113 - 0x71
      13'h128E: dout  = 8'b01110101; // 4750 : 117 - 0x75
      13'h128F: dout  = 8'b01110100; // 4751 : 116 - 0x74
      13'h1290: dout  = 8'b10001111; // 4752 : 143 - 0x8f -- Background 0x29
      13'h1291: dout  = 8'b11001111; // 4753 : 207 - 0xcf
      13'h1292: dout  = 8'b10001111; // 4754 : 143 - 0x8f
      13'h1293: dout  = 8'b11001111; // 4755 : 207 - 0xcf
      13'h1294: dout  = 8'b10010000; // 4756 : 144 - 0x90
      13'h1295: dout  = 8'b11100000; // 4757 : 224 - 0xe0
      13'h1296: dout  = 8'b11101010; // 4758 : 234 - 0xea
      13'h1297: dout  = 8'b11111111; // 4759 : 255 - 0xff
      13'h1298: dout  = 8'b01110000; // 4760 : 112 - 0x70
      13'h1299: dout  = 8'b01110111; // 4761 : 119 - 0x77
      13'h129A: dout  = 8'b01110111; // 4762 : 119 - 0x77
      13'h129B: dout  = 8'b01110000; // 4763 : 112 - 0x70
      13'h129C: dout  = 8'b01101111; // 4764 : 111 - 0x6f
      13'h129D: dout  = 8'b01011111; // 4765 :  95 - 0x5f
      13'h129E: dout  = 8'b00010101; // 4766 :  21 - 0x15
      13'h129F: dout  = 8'b00000000; // 4767 :   0 - 0x0
      13'h12A0: dout  = 8'b11111111; // 4768 : 255 - 0xff -- Background 0x2a
      13'h12A1: dout  = 8'b11011011; // 4769 : 219 - 0xdb
      13'h12A2: dout  = 8'b11000111; // 4770 : 199 - 0xc7
      13'h12A3: dout  = 8'b11101001; // 4771 : 233 - 0xe9
      13'h12A4: dout  = 8'b11110011; // 4772 : 243 - 0xf3
      13'h12A5: dout  = 8'b11110001; // 4773 : 241 - 0xf1
      13'h12A6: dout  = 8'b11010011; // 4774 : 211 - 0xd3
      13'h12A7: dout  = 8'b11010001; // 4775 : 209 - 0xd1
      13'h12A8: dout  = 8'b00000000; // 4776 :   0 - 0x0
      13'h12A9: dout  = 8'b01111100; // 4777 : 124 - 0x7c
      13'h12AA: dout  = 8'b10111000; // 4778 : 184 - 0xb8
      13'h12AB: dout  = 8'b11010110; // 4779 : 214 - 0xd6
      13'h12AC: dout  = 8'b10101100; // 4780 : 172 - 0xac
      13'h12AD: dout  = 8'b10001110; // 4781 : 142 - 0x8e
      13'h12AE: dout  = 8'b10101100; // 4782 : 172 - 0xac
      13'h12AF: dout  = 8'b00101110; // 4783 :  46 - 0x2e
      13'h12B0: dout  = 8'b11110011; // 4784 : 243 - 0xf3 -- Background 0x2b
      13'h12B1: dout  = 8'b11110001; // 4785 : 241 - 0xf1
      13'h12B2: dout  = 8'b11110011; // 4786 : 243 - 0xf3
      13'h12B3: dout  = 8'b11110001; // 4787 : 241 - 0xf1
      13'h12B4: dout  = 8'b00001011; // 4788 :  11 - 0xb
      13'h12B5: dout  = 8'b00000101; // 4789 :   5 - 0x5
      13'h12B6: dout  = 8'b10101011; // 4790 : 171 - 0xab
      13'h12B7: dout  = 8'b11111111; // 4791 : 255 - 0xff
      13'h12B8: dout  = 8'b00001100; // 4792 :  12 - 0xc
      13'h12B9: dout  = 8'b11101110; // 4793 : 238 - 0xee
      13'h12BA: dout  = 8'b11101100; // 4794 : 236 - 0xec
      13'h12BB: dout  = 8'b00001110; // 4795 :  14 - 0xe
      13'h12BC: dout  = 8'b11110100; // 4796 : 244 - 0xf4
      13'h12BD: dout  = 8'b11111010; // 4797 : 250 - 0xfa
      13'h12BE: dout  = 8'b01010100; // 4798 :  84 - 0x54
      13'h12BF: dout  = 8'b00000000; // 4799 :   0 - 0x0
      13'h12C0: dout  = 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout  = 8'b00000000; // 4801 :   0 - 0x0
      13'h12C2: dout  = 8'b00000000; // 4802 :   0 - 0x0
      13'h12C3: dout  = 8'b00000000; // 4803 :   0 - 0x0
      13'h12C4: dout  = 8'b00000000; // 4804 :   0 - 0x0
      13'h12C5: dout  = 8'b00000000; // 4805 :   0 - 0x0
      13'h12C6: dout  = 8'b00000000; // 4806 :   0 - 0x0
      13'h12C7: dout  = 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout  = 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout  = 8'b00000000; // 4809 :   0 - 0x0
      13'h12CA: dout  = 8'b00000000; // 4810 :   0 - 0x0
      13'h12CB: dout  = 8'b00000000; // 4811 :   0 - 0x0
      13'h12CC: dout  = 8'b00000000; // 4812 :   0 - 0x0
      13'h12CD: dout  = 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout  = 8'b00000000; // 4814 :   0 - 0x0
      13'h12CF: dout  = 8'b00000000; // 4815 :   0 - 0x0
      13'h12D0: dout  = 8'b00101111; // 4816 :  47 - 0x2f -- Background 0x2d
      13'h12D1: dout  = 8'b01001111; // 4817 :  79 - 0x4f
      13'h12D2: dout  = 8'b01001111; // 4818 :  79 - 0x4f
      13'h12D3: dout  = 8'b01001111; // 4819 :  79 - 0x4f
      13'h12D4: dout  = 8'b01001111; // 4820 :  79 - 0x4f
      13'h12D5: dout  = 8'b00100111; // 4821 :  39 - 0x27
      13'h12D6: dout  = 8'b00010000; // 4822 :  16 - 0x10
      13'h12D7: dout  = 8'b00001111; // 4823 :  15 - 0xf
      13'h12D8: dout  = 8'b00011110; // 4824 :  30 - 0x1e
      13'h12D9: dout  = 8'b00111110; // 4825 :  62 - 0x3e
      13'h12DA: dout  = 8'b00111110; // 4826 :  62 - 0x3e
      13'h12DB: dout  = 8'b00111110; // 4827 :  62 - 0x3e
      13'h12DC: dout  = 8'b00111111; // 4828 :  63 - 0x3f
      13'h12DD: dout  = 8'b00011110; // 4829 :  30 - 0x1e
      13'h12DE: dout  = 8'b00001111; // 4830 :  15 - 0xf
      13'h12DF: dout  = 8'b00000000; // 4831 :   0 - 0x0
      13'h12E0: dout  = 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout  = 8'b00000000; // 4833 :   0 - 0x0
      13'h12E2: dout  = 8'b00000000; // 4834 :   0 - 0x0
      13'h12E3: dout  = 8'b00000000; // 4835 :   0 - 0x0
      13'h12E4: dout  = 8'b00000000; // 4836 :   0 - 0x0
      13'h12E5: dout  = 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout  = 8'b00000000; // 4838 :   0 - 0x0
      13'h12E7: dout  = 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout  = 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout  = 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout  = 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout  = 8'b00000000; // 4843 :   0 - 0x0
      13'h12EC: dout  = 8'b00000000; // 4844 :   0 - 0x0
      13'h12ED: dout  = 8'b00000000; // 4845 :   0 - 0x0
      13'h12EE: dout  = 8'b00000000; // 4846 :   0 - 0x0
      13'h12EF: dout  = 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout  = 8'b11110100; // 4848 : 244 - 0xf4 -- Background 0x2f
      13'h12F1: dout  = 8'b11110010; // 4849 : 242 - 0xf2
      13'h12F2: dout  = 8'b11110010; // 4850 : 242 - 0xf2
      13'h12F3: dout  = 8'b11110010; // 4851 : 242 - 0xf2
      13'h12F4: dout  = 8'b11110010; // 4852 : 242 - 0xf2
      13'h12F5: dout  = 8'b11100100; // 4853 : 228 - 0xe4
      13'h12F6: dout  = 8'b00001000; // 4854 :   8 - 0x8
      13'h12F7: dout  = 8'b11110000; // 4855 : 240 - 0xf0
      13'h12F8: dout  = 8'b01111000; // 4856 : 120 - 0x78
      13'h12F9: dout  = 8'b01111100; // 4857 : 124 - 0x7c
      13'h12FA: dout  = 8'b01111100; // 4858 : 124 - 0x7c
      13'h12FB: dout  = 8'b01111100; // 4859 : 124 - 0x7c
      13'h12FC: dout  = 8'b11111100; // 4860 : 252 - 0xfc
      13'h12FD: dout  = 8'b01111000; // 4861 : 120 - 0x78
      13'h12FE: dout  = 8'b11110000; // 4862 : 240 - 0xf0
      13'h12FF: dout  = 8'b00000000; // 4863 :   0 - 0x0
      13'h1300: dout  = 8'b00011000; // 4864 :  24 - 0x18 -- Background 0x30
      13'h1301: dout  = 8'b00100100; // 4865 :  36 - 0x24
      13'h1302: dout  = 8'b01000010; // 4866 :  66 - 0x42
      13'h1303: dout  = 8'b10100101; // 4867 : 165 - 0xa5
      13'h1304: dout  = 8'b11100111; // 4868 : 231 - 0xe7
      13'h1305: dout  = 8'b00100100; // 4869 :  36 - 0x24
      13'h1306: dout  = 8'b00100100; // 4870 :  36 - 0x24
      13'h1307: dout  = 8'b00111100; // 4871 :  60 - 0x3c
      13'h1308: dout  = 8'b00000000; // 4872 :   0 - 0x0
      13'h1309: dout  = 8'b00011000; // 4873 :  24 - 0x18
      13'h130A: dout  = 8'b00111100; // 4874 :  60 - 0x3c
      13'h130B: dout  = 8'b01011010; // 4875 :  90 - 0x5a
      13'h130C: dout  = 8'b00011000; // 4876 :  24 - 0x18
      13'h130D: dout  = 8'b00011000; // 4877 :  24 - 0x18
      13'h130E: dout  = 8'b00011000; // 4878 :  24 - 0x18
      13'h130F: dout  = 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout  = 8'b00111100; // 4880 :  60 - 0x3c -- Background 0x31
      13'h1311: dout  = 8'b00100100; // 4881 :  36 - 0x24
      13'h1312: dout  = 8'b00100100; // 4882 :  36 - 0x24
      13'h1313: dout  = 8'b01100110; // 4883 : 102 - 0x66
      13'h1314: dout  = 8'b10100101; // 4884 : 165 - 0xa5
      13'h1315: dout  = 8'b01000010; // 4885 :  66 - 0x42
      13'h1316: dout  = 8'b00100100; // 4886 :  36 - 0x24
      13'h1317: dout  = 8'b00011000; // 4887 :  24 - 0x18
      13'h1318: dout  = 8'b00000000; // 4888 :   0 - 0x0
      13'h1319: dout  = 8'b00011000; // 4889 :  24 - 0x18
      13'h131A: dout  = 8'b00011000; // 4890 :  24 - 0x18
      13'h131B: dout  = 8'b00011000; // 4891 :  24 - 0x18
      13'h131C: dout  = 8'b01011010; // 4892 :  90 - 0x5a
      13'h131D: dout  = 8'b00111100; // 4893 :  60 - 0x3c
      13'h131E: dout  = 8'b00011000; // 4894 :  24 - 0x18
      13'h131F: dout  = 8'b00000000; // 4895 :   0 - 0x0
      13'h1320: dout  = 8'b00000010; // 4896 :   2 - 0x2 -- Background 0x32
      13'h1321: dout  = 8'b00000010; // 4897 :   2 - 0x2
      13'h1322: dout  = 8'b00000011; // 4898 :   3 - 0x3
      13'h1323: dout  = 8'b00000010; // 4899 :   2 - 0x2
      13'h1324: dout  = 8'b00000010; // 4900 :   2 - 0x2
      13'h1325: dout  = 8'b00000010; // 4901 :   2 - 0x2
      13'h1326: dout  = 8'b00000011; // 4902 :   3 - 0x3
      13'h1327: dout  = 8'b00000010; // 4903 :   2 - 0x2
      13'h1328: dout  = 8'b00000001; // 4904 :   1 - 0x1
      13'h1329: dout  = 8'b00000001; // 4905 :   1 - 0x1
      13'h132A: dout  = 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout  = 8'b00000001; // 4907 :   1 - 0x1
      13'h132C: dout  = 8'b00000001; // 4908 :   1 - 0x1
      13'h132D: dout  = 8'b00000001; // 4909 :   1 - 0x1
      13'h132E: dout  = 8'b00000000; // 4910 :   0 - 0x0
      13'h132F: dout  = 8'b00000001; // 4911 :   1 - 0x1
      13'h1330: dout  = 8'b01000000; // 4912 :  64 - 0x40 -- Background 0x33
      13'h1331: dout  = 8'b11000000; // 4913 : 192 - 0xc0
      13'h1332: dout  = 8'b01000000; // 4914 :  64 - 0x40
      13'h1333: dout  = 8'b01000000; // 4915 :  64 - 0x40
      13'h1334: dout  = 8'b01000000; // 4916 :  64 - 0x40
      13'h1335: dout  = 8'b11000000; // 4917 : 192 - 0xc0
      13'h1336: dout  = 8'b01000000; // 4918 :  64 - 0x40
      13'h1337: dout  = 8'b01000000; // 4919 :  64 - 0x40
      13'h1338: dout  = 8'b10000000; // 4920 : 128 - 0x80
      13'h1339: dout  = 8'b00000000; // 4921 :   0 - 0x0
      13'h133A: dout  = 8'b10000000; // 4922 : 128 - 0x80
      13'h133B: dout  = 8'b10000000; // 4923 : 128 - 0x80
      13'h133C: dout  = 8'b10000000; // 4924 : 128 - 0x80
      13'h133D: dout  = 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout  = 8'b10000000; // 4926 : 128 - 0x80
      13'h133F: dout  = 8'b10000000; // 4927 : 128 - 0x80
      13'h1340: dout  = 8'b00000000; // 4928 :   0 - 0x0 -- Background 0x34
      13'h1341: dout  = 8'b00011000; // 4929 :  24 - 0x18
      13'h1342: dout  = 8'b00111100; // 4930 :  60 - 0x3c
      13'h1343: dout  = 8'b01100010; // 4931 :  98 - 0x62
      13'h1344: dout  = 8'b01100001; // 4932 :  97 - 0x61
      13'h1345: dout  = 8'b11000000; // 4933 : 192 - 0xc0
      13'h1346: dout  = 8'b11000000; // 4934 : 192 - 0xc0
      13'h1347: dout  = 8'b11000000; // 4935 : 192 - 0xc0
      13'h1348: dout  = 8'b00000000; // 4936 :   0 - 0x0
      13'h1349: dout  = 8'b00000000; // 4937 :   0 - 0x0
      13'h134A: dout  = 8'b00011000; // 4938 :  24 - 0x18
      13'h134B: dout  = 8'b00111100; // 4939 :  60 - 0x3c
      13'h134C: dout  = 8'b00111110; // 4940 :  62 - 0x3e
      13'h134D: dout  = 8'b01111111; // 4941 : 127 - 0x7f
      13'h134E: dout  = 8'b01111111; // 4942 : 127 - 0x7f
      13'h134F: dout  = 8'b01111111; // 4943 : 127 - 0x7f
      13'h1350: dout  = 8'b01100000; // 4944 :  96 - 0x60 -- Background 0x35
      13'h1351: dout  = 8'b01100000; // 4945 :  96 - 0x60
      13'h1352: dout  = 8'b00110000; // 4946 :  48 - 0x30
      13'h1353: dout  = 8'b00011000; // 4947 :  24 - 0x18
      13'h1354: dout  = 8'b00001100; // 4948 :  12 - 0xc
      13'h1355: dout  = 8'b00000110; // 4949 :   6 - 0x6
      13'h1356: dout  = 8'b00000010; // 4950 :   2 - 0x2
      13'h1357: dout  = 8'b00000001; // 4951 :   1 - 0x1
      13'h1358: dout  = 8'b00111111; // 4952 :  63 - 0x3f
      13'h1359: dout  = 8'b00111111; // 4953 :  63 - 0x3f
      13'h135A: dout  = 8'b00011111; // 4954 :  31 - 0x1f
      13'h135B: dout  = 8'b00001111; // 4955 :  15 - 0xf
      13'h135C: dout  = 8'b00000111; // 4956 :   7 - 0x7
      13'h135D: dout  = 8'b00000011; // 4957 :   3 - 0x3
      13'h135E: dout  = 8'b00000001; // 4958 :   1 - 0x1
      13'h135F: dout  = 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout  = 8'b00000000; // 4960 :   0 - 0x0 -- Background 0x36
      13'h1361: dout  = 8'b00011000; // 4961 :  24 - 0x18
      13'h1362: dout  = 8'b00100100; // 4962 :  36 - 0x24
      13'h1363: dout  = 8'b01000010; // 4963 :  66 - 0x42
      13'h1364: dout  = 8'b10000010; // 4964 : 130 - 0x82
      13'h1365: dout  = 8'b00000001; // 4965 :   1 - 0x1
      13'h1366: dout  = 8'b00000001; // 4966 :   1 - 0x1
      13'h1367: dout  = 8'b00000001; // 4967 :   1 - 0x1
      13'h1368: dout  = 8'b00000000; // 4968 :   0 - 0x0
      13'h1369: dout  = 8'b00000000; // 4969 :   0 - 0x0
      13'h136A: dout  = 8'b00011000; // 4970 :  24 - 0x18
      13'h136B: dout  = 8'b00111100; // 4971 :  60 - 0x3c
      13'h136C: dout  = 8'b01111100; // 4972 : 124 - 0x7c
      13'h136D: dout  = 8'b11111110; // 4973 : 254 - 0xfe
      13'h136E: dout  = 8'b11111110; // 4974 : 254 - 0xfe
      13'h136F: dout  = 8'b11111110; // 4975 : 254 - 0xfe
      13'h1370: dout  = 8'b00000010; // 4976 :   2 - 0x2 -- Background 0x37
      13'h1371: dout  = 8'b00000010; // 4977 :   2 - 0x2
      13'h1372: dout  = 8'b00000100; // 4978 :   4 - 0x4
      13'h1373: dout  = 8'b00001000; // 4979 :   8 - 0x8
      13'h1374: dout  = 8'b00010000; // 4980 :  16 - 0x10
      13'h1375: dout  = 8'b00100000; // 4981 :  32 - 0x20
      13'h1376: dout  = 8'b01000000; // 4982 :  64 - 0x40
      13'h1377: dout  = 8'b10000000; // 4983 : 128 - 0x80
      13'h1378: dout  = 8'b11111100; // 4984 : 252 - 0xfc
      13'h1379: dout  = 8'b11111100; // 4985 : 252 - 0xfc
      13'h137A: dout  = 8'b11111000; // 4986 : 248 - 0xf8
      13'h137B: dout  = 8'b11110000; // 4987 : 240 - 0xf0
      13'h137C: dout  = 8'b11100000; // 4988 : 224 - 0xe0
      13'h137D: dout  = 8'b11000000; // 4989 : 192 - 0xc0
      13'h137E: dout  = 8'b10000000; // 4990 : 128 - 0x80
      13'h137F: dout  = 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout  = 8'b00000000; // 4992 :   0 - 0x0 -- Background 0x38
      13'h1381: dout  = 8'b00000110; // 4993 :   6 - 0x6
      13'h1382: dout  = 8'b00001101; // 4994 :  13 - 0xd
      13'h1383: dout  = 8'b00001100; // 4995 :  12 - 0xc
      13'h1384: dout  = 8'b00001100; // 4996 :  12 - 0xc
      13'h1385: dout  = 8'b00000110; // 4997 :   6 - 0x6
      13'h1386: dout  = 8'b00000010; // 4998 :   2 - 0x2
      13'h1387: dout  = 8'b00000001; // 4999 :   1 - 0x1
      13'h1388: dout  = 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout  = 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout  = 8'b00000110; // 5002 :   6 - 0x6
      13'h138B: dout  = 8'b00000111; // 5003 :   7 - 0x7
      13'h138C: dout  = 8'b00000111; // 5004 :   7 - 0x7
      13'h138D: dout  = 8'b00000011; // 5005 :   3 - 0x3
      13'h138E: dout  = 8'b00000001; // 5006 :   1 - 0x1
      13'h138F: dout  = 8'b00000000; // 5007 :   0 - 0x0
      13'h1390: dout  = 8'b11111111; // 5008 : 255 - 0xff -- Background 0x39
      13'h1391: dout  = 8'b00000000; // 5009 :   0 - 0x0
      13'h1392: dout  = 8'b00000000; // 5010 :   0 - 0x0
      13'h1393: dout  = 8'b00000000; // 5011 :   0 - 0x0
      13'h1394: dout  = 8'b00000000; // 5012 :   0 - 0x0
      13'h1395: dout  = 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout  = 8'b00000000; // 5014 :   0 - 0x0
      13'h1397: dout  = 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout  = 8'b00000000; // 5016 :   0 - 0x0
      13'h1399: dout  = 8'b00000000; // 5017 :   0 - 0x0
      13'h139A: dout  = 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout  = 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout  = 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout  = 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout  = 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout  = 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout  = 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout  = 8'b01100000; // 5025 :  96 - 0x60
      13'h13A2: dout  = 8'b10010000; // 5026 : 144 - 0x90
      13'h13A3: dout  = 8'b00010000; // 5027 :  16 - 0x10
      13'h13A4: dout  = 8'b00010000; // 5028 :  16 - 0x10
      13'h13A5: dout  = 8'b00100000; // 5029 :  32 - 0x20
      13'h13A6: dout  = 8'b01000000; // 5030 :  64 - 0x40
      13'h13A7: dout  = 8'b10000000; // 5031 : 128 - 0x80
      13'h13A8: dout  = 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout  = 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout  = 8'b01100000; // 5034 :  96 - 0x60
      13'h13AB: dout  = 8'b11100000; // 5035 : 224 - 0xe0
      13'h13AC: dout  = 8'b11100000; // 5036 : 224 - 0xe0
      13'h13AD: dout  = 8'b11000000; // 5037 : 192 - 0xc0
      13'h13AE: dout  = 8'b10000000; // 5038 : 128 - 0x80
      13'h13AF: dout  = 8'b00000000; // 5039 :   0 - 0x0
      13'h13B0: dout  = 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout  = 8'b01010100; // 5041 :  84 - 0x54
      13'h13B2: dout  = 8'b00000010; // 5042 :   2 - 0x2
      13'h13B3: dout  = 8'b01000000; // 5043 :  64 - 0x40
      13'h13B4: dout  = 8'b00000010; // 5044 :   2 - 0x2
      13'h13B5: dout  = 8'b01000000; // 5045 :  64 - 0x40
      13'h13B6: dout  = 8'b00101010; // 5046 :  42 - 0x2a
      13'h13B7: dout  = 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout  = 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout  = 8'b00101010; // 5049 :  42 - 0x2a
      13'h13BA: dout  = 8'b01000000; // 5050 :  64 - 0x40
      13'h13BB: dout  = 8'b00000010; // 5051 :   2 - 0x2
      13'h13BC: dout  = 8'b01000000; // 5052 :  64 - 0x40
      13'h13BD: dout  = 8'b00000010; // 5053 :   2 - 0x2
      13'h13BE: dout  = 8'b01010100; // 5054 :  84 - 0x54
      13'h13BF: dout  = 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout  = 8'b11111111; // 5056 : 255 - 0xff -- Background 0x3c
      13'h13C1: dout  = 8'b11111111; // 5057 : 255 - 0xff
      13'h13C2: dout  = 8'b11111111; // 5058 : 255 - 0xff
      13'h13C3: dout  = 8'b11111111; // 5059 : 255 - 0xff
      13'h13C4: dout  = 8'b11111111; // 5060 : 255 - 0xff
      13'h13C5: dout  = 8'b11111111; // 5061 : 255 - 0xff
      13'h13C6: dout  = 8'b11111111; // 5062 : 255 - 0xff
      13'h13C7: dout  = 8'b11111111; // 5063 : 255 - 0xff
      13'h13C8: dout  = 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout  = 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout  = 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout  = 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout  = 8'b00000000; // 5068 :   0 - 0x0
      13'h13CD: dout  = 8'b00000000; // 5069 :   0 - 0x0
      13'h13CE: dout  = 8'b00000000; // 5070 :   0 - 0x0
      13'h13CF: dout  = 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout  = 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout  = 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout  = 8'b00000000; // 5074 :   0 - 0x0
      13'h13D3: dout  = 8'b00000000; // 5075 :   0 - 0x0
      13'h13D4: dout  = 8'b00000000; // 5076 :   0 - 0x0
      13'h13D5: dout  = 8'b00000000; // 5077 :   0 - 0x0
      13'h13D6: dout  = 8'b00000000; // 5078 :   0 - 0x0
      13'h13D7: dout  = 8'b00000000; // 5079 :   0 - 0x0
      13'h13D8: dout  = 8'b11111111; // 5080 : 255 - 0xff
      13'h13D9: dout  = 8'b11111111; // 5081 : 255 - 0xff
      13'h13DA: dout  = 8'b11111111; // 5082 : 255 - 0xff
      13'h13DB: dout  = 8'b11111111; // 5083 : 255 - 0xff
      13'h13DC: dout  = 8'b11111111; // 5084 : 255 - 0xff
      13'h13DD: dout  = 8'b11111111; // 5085 : 255 - 0xff
      13'h13DE: dout  = 8'b11111111; // 5086 : 255 - 0xff
      13'h13DF: dout  = 8'b11111111; // 5087 : 255 - 0xff
      13'h13E0: dout  = 8'b11111111; // 5088 : 255 - 0xff -- Background 0x3e
      13'h13E1: dout  = 8'b11111111; // 5089 : 255 - 0xff
      13'h13E2: dout  = 8'b11111111; // 5090 : 255 - 0xff
      13'h13E3: dout  = 8'b11111111; // 5091 : 255 - 0xff
      13'h13E4: dout  = 8'b11111111; // 5092 : 255 - 0xff
      13'h13E5: dout  = 8'b11111111; // 5093 : 255 - 0xff
      13'h13E6: dout  = 8'b11111111; // 5094 : 255 - 0xff
      13'h13E7: dout  = 8'b11111111; // 5095 : 255 - 0xff
      13'h13E8: dout  = 8'b11111111; // 5096 : 255 - 0xff
      13'h13E9: dout  = 8'b11111111; // 5097 : 255 - 0xff
      13'h13EA: dout  = 8'b11111111; // 5098 : 255 - 0xff
      13'h13EB: dout  = 8'b11111111; // 5099 : 255 - 0xff
      13'h13EC: dout  = 8'b11111111; // 5100 : 255 - 0xff
      13'h13ED: dout  = 8'b11111111; // 5101 : 255 - 0xff
      13'h13EE: dout  = 8'b11111111; // 5102 : 255 - 0xff
      13'h13EF: dout  = 8'b11111111; // 5103 : 255 - 0xff
      13'h13F0: dout  = 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout  = 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout  = 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout  = 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout  = 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout  = 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout  = 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout  = 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout  = 8'b00000000; // 5112 :   0 - 0x0
      13'h13F9: dout  = 8'b00000000; // 5113 :   0 - 0x0
      13'h13FA: dout  = 8'b00000000; // 5114 :   0 - 0x0
      13'h13FB: dout  = 8'b00000000; // 5115 :   0 - 0x0
      13'h13FC: dout  = 8'b00000000; // 5116 :   0 - 0x0
      13'h13FD: dout  = 8'b00000000; // 5117 :   0 - 0x0
      13'h13FE: dout  = 8'b00000000; // 5118 :   0 - 0x0
      13'h13FF: dout  = 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout  = 8'b00111100; // 5120 :  60 - 0x3c -- Background 0x40
      13'h1401: dout  = 8'b01000010; // 5121 :  66 - 0x42
      13'h1402: dout  = 8'b10011001; // 5122 : 153 - 0x99
      13'h1403: dout  = 8'b10100101; // 5123 : 165 - 0xa5
      13'h1404: dout  = 8'b10100101; // 5124 : 165 - 0xa5
      13'h1405: dout  = 8'b10011010; // 5125 : 154 - 0x9a
      13'h1406: dout  = 8'b01000000; // 5126 :  64 - 0x40
      13'h1407: dout  = 8'b00111100; // 5127 :  60 - 0x3c
      13'h1408: dout  = 8'b00000000; // 5128 :   0 - 0x0
      13'h1409: dout  = 8'b00000000; // 5129 :   0 - 0x0
      13'h140A: dout  = 8'b00000000; // 5130 :   0 - 0x0
      13'h140B: dout  = 8'b00000000; // 5131 :   0 - 0x0
      13'h140C: dout  = 8'b00000000; // 5132 :   0 - 0x0
      13'h140D: dout  = 8'b00000000; // 5133 :   0 - 0x0
      13'h140E: dout  = 8'b00000000; // 5134 :   0 - 0x0
      13'h140F: dout  = 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout  = 8'b00001100; // 5136 :  12 - 0xc -- Background 0x41
      13'h1411: dout  = 8'b00010010; // 5137 :  18 - 0x12
      13'h1412: dout  = 8'b00100010; // 5138 :  34 - 0x22
      13'h1413: dout  = 8'b00100010; // 5139 :  34 - 0x22
      13'h1414: dout  = 8'b01111110; // 5140 : 126 - 0x7e
      13'h1415: dout  = 8'b00100010; // 5141 :  34 - 0x22
      13'h1416: dout  = 8'b00100100; // 5142 :  36 - 0x24
      13'h1417: dout  = 8'b00000000; // 5143 :   0 - 0x0
      13'h1418: dout  = 8'b00000000; // 5144 :   0 - 0x0
      13'h1419: dout  = 8'b00000000; // 5145 :   0 - 0x0
      13'h141A: dout  = 8'b00000000; // 5146 :   0 - 0x0
      13'h141B: dout  = 8'b00000000; // 5147 :   0 - 0x0
      13'h141C: dout  = 8'b00000000; // 5148 :   0 - 0x0
      13'h141D: dout  = 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout  = 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout  = 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout  = 8'b00111100; // 5152 :  60 - 0x3c -- Background 0x42
      13'h1421: dout  = 8'b01000010; // 5153 :  66 - 0x42
      13'h1422: dout  = 8'b01010010; // 5154 :  82 - 0x52
      13'h1423: dout  = 8'b00011100; // 5155 :  28 - 0x1c
      13'h1424: dout  = 8'b00010010; // 5156 :  18 - 0x12
      13'h1425: dout  = 8'b00110010; // 5157 :  50 - 0x32
      13'h1426: dout  = 8'b00011100; // 5158 :  28 - 0x1c
      13'h1427: dout  = 8'b00000000; // 5159 :   0 - 0x0
      13'h1428: dout  = 8'b00000000; // 5160 :   0 - 0x0
      13'h1429: dout  = 8'b00000000; // 5161 :   0 - 0x0
      13'h142A: dout  = 8'b00000000; // 5162 :   0 - 0x0
      13'h142B: dout  = 8'b00000000; // 5163 :   0 - 0x0
      13'h142C: dout  = 8'b00000000; // 5164 :   0 - 0x0
      13'h142D: dout  = 8'b00000000; // 5165 :   0 - 0x0
      13'h142E: dout  = 8'b00000000; // 5166 :   0 - 0x0
      13'h142F: dout  = 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout  = 8'b00011000; // 5168 :  24 - 0x18 -- Background 0x43
      13'h1431: dout  = 8'b00100100; // 5169 :  36 - 0x24
      13'h1432: dout  = 8'b01010100; // 5170 :  84 - 0x54
      13'h1433: dout  = 8'b01001000; // 5171 :  72 - 0x48
      13'h1434: dout  = 8'b01000010; // 5172 :  66 - 0x42
      13'h1435: dout  = 8'b00100100; // 5173 :  36 - 0x24
      13'h1436: dout  = 8'b00011000; // 5174 :  24 - 0x18
      13'h1437: dout  = 8'b00000000; // 5175 :   0 - 0x0
      13'h1438: dout  = 8'b00000000; // 5176 :   0 - 0x0
      13'h1439: dout  = 8'b00000000; // 5177 :   0 - 0x0
      13'h143A: dout  = 8'b00000000; // 5178 :   0 - 0x0
      13'h143B: dout  = 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout  = 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout  = 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout  = 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout  = 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout  = 8'b01011000; // 5184 :  88 - 0x58 -- Background 0x44
      13'h1441: dout  = 8'b11100100; // 5185 : 228 - 0xe4
      13'h1442: dout  = 8'b01000010; // 5186 :  66 - 0x42
      13'h1443: dout  = 8'b01000010; // 5187 :  66 - 0x42
      13'h1444: dout  = 8'b00100010; // 5188 :  34 - 0x22
      13'h1445: dout  = 8'b01100100; // 5189 : 100 - 0x64
      13'h1446: dout  = 8'b00111000; // 5190 :  56 - 0x38
      13'h1447: dout  = 8'b00000000; // 5191 :   0 - 0x0
      13'h1448: dout  = 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout  = 8'b00000000; // 5193 :   0 - 0x0
      13'h144A: dout  = 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout  = 8'b00000000; // 5195 :   0 - 0x0
      13'h144C: dout  = 8'b00000000; // 5196 :   0 - 0x0
      13'h144D: dout  = 8'b00000000; // 5197 :   0 - 0x0
      13'h144E: dout  = 8'b00000000; // 5198 :   0 - 0x0
      13'h144F: dout  = 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout  = 8'b00011100; // 5200 :  28 - 0x1c -- Background 0x45
      13'h1451: dout  = 8'b00100000; // 5201 :  32 - 0x20
      13'h1452: dout  = 8'b00100000; // 5202 :  32 - 0x20
      13'h1453: dout  = 8'b00101100; // 5203 :  44 - 0x2c
      13'h1454: dout  = 8'b01110000; // 5204 : 112 - 0x70
      13'h1455: dout  = 8'b00100010; // 5205 :  34 - 0x22
      13'h1456: dout  = 8'b00011100; // 5206 :  28 - 0x1c
      13'h1457: dout  = 8'b00000000; // 5207 :   0 - 0x0
      13'h1458: dout  = 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout  = 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout  = 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout  = 8'b00000000; // 5211 :   0 - 0x0
      13'h145C: dout  = 8'b00000000; // 5212 :   0 - 0x0
      13'h145D: dout  = 8'b00000000; // 5213 :   0 - 0x0
      13'h145E: dout  = 8'b00000000; // 5214 :   0 - 0x0
      13'h145F: dout  = 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout  = 8'b00011100; // 5216 :  28 - 0x1c -- Background 0x46
      13'h1461: dout  = 8'b00100000; // 5217 :  32 - 0x20
      13'h1462: dout  = 8'b00100000; // 5218 :  32 - 0x20
      13'h1463: dout  = 8'b00101100; // 5219 :  44 - 0x2c
      13'h1464: dout  = 8'b01110000; // 5220 : 112 - 0x70
      13'h1465: dout  = 8'b00010000; // 5221 :  16 - 0x10
      13'h1466: dout  = 8'b00010000; // 5222 :  16 - 0x10
      13'h1467: dout  = 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout  = 8'b00000000; // 5224 :   0 - 0x0
      13'h1469: dout  = 8'b00000000; // 5225 :   0 - 0x0
      13'h146A: dout  = 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout  = 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout  = 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout  = 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout  = 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout  = 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout  = 8'b00011000; // 5232 :  24 - 0x18 -- Background 0x47
      13'h1471: dout  = 8'b00100100; // 5233 :  36 - 0x24
      13'h1472: dout  = 8'b01000000; // 5234 :  64 - 0x40
      13'h1473: dout  = 8'b01001110; // 5235 :  78 - 0x4e
      13'h1474: dout  = 8'b01000010; // 5236 :  66 - 0x42
      13'h1475: dout  = 8'b00100100; // 5237 :  36 - 0x24
      13'h1476: dout  = 8'b00011000; // 5238 :  24 - 0x18
      13'h1477: dout  = 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout  = 8'b00000000; // 5240 :   0 - 0x0
      13'h1479: dout  = 8'b00000000; // 5241 :   0 - 0x0
      13'h147A: dout  = 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout  = 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout  = 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout  = 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout  = 8'b00000000; // 5246 :   0 - 0x0
      13'h147F: dout  = 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout  = 8'b00100000; // 5248 :  32 - 0x20 -- Background 0x48
      13'h1481: dout  = 8'b01000100; // 5249 :  68 - 0x44
      13'h1482: dout  = 8'b01000100; // 5250 :  68 - 0x44
      13'h1483: dout  = 8'b01000100; // 5251 :  68 - 0x44
      13'h1484: dout  = 8'b11111100; // 5252 : 252 - 0xfc
      13'h1485: dout  = 8'b01000100; // 5253 :  68 - 0x44
      13'h1486: dout  = 8'b01001000; // 5254 :  72 - 0x48
      13'h1487: dout  = 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout  = 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout  = 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout  = 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout  = 8'b00000000; // 5259 :   0 - 0x0
      13'h148C: dout  = 8'b00000000; // 5260 :   0 - 0x0
      13'h148D: dout  = 8'b00000000; // 5261 :   0 - 0x0
      13'h148E: dout  = 8'b00000000; // 5262 :   0 - 0x0
      13'h148F: dout  = 8'b00000000; // 5263 :   0 - 0x0
      13'h1490: dout  = 8'b00010000; // 5264 :  16 - 0x10 -- Background 0x49
      13'h1491: dout  = 8'b00010000; // 5265 :  16 - 0x10
      13'h1492: dout  = 8'b00010000; // 5266 :  16 - 0x10
      13'h1493: dout  = 8'b00010000; // 5267 :  16 - 0x10
      13'h1494: dout  = 8'b00010000; // 5268 :  16 - 0x10
      13'h1495: dout  = 8'b00001000; // 5269 :   8 - 0x8
      13'h1496: dout  = 8'b00001000; // 5270 :   8 - 0x8
      13'h1497: dout  = 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout  = 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout  = 8'b00000000; // 5273 :   0 - 0x0
      13'h149A: dout  = 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout  = 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout  = 8'b00000000; // 5276 :   0 - 0x0
      13'h149D: dout  = 8'b00000000; // 5277 :   0 - 0x0
      13'h149E: dout  = 8'b00000000; // 5278 :   0 - 0x0
      13'h149F: dout  = 8'b00000000; // 5279 :   0 - 0x0
      13'h14A0: dout  = 8'b00001000; // 5280 :   8 - 0x8 -- Background 0x4a
      13'h14A1: dout  = 8'b00001000; // 5281 :   8 - 0x8
      13'h14A2: dout  = 8'b00000100; // 5282 :   4 - 0x4
      13'h14A3: dout  = 8'b00000100; // 5283 :   4 - 0x4
      13'h14A4: dout  = 8'b01000100; // 5284 :  68 - 0x44
      13'h14A5: dout  = 8'b01001000; // 5285 :  72 - 0x48
      13'h14A6: dout  = 8'b00110000; // 5286 :  48 - 0x30
      13'h14A7: dout  = 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout  = 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout  = 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout  = 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout  = 8'b00000000; // 5291 :   0 - 0x0
      13'h14AC: dout  = 8'b00000000; // 5292 :   0 - 0x0
      13'h14AD: dout  = 8'b00000000; // 5293 :   0 - 0x0
      13'h14AE: dout  = 8'b00000000; // 5294 :   0 - 0x0
      13'h14AF: dout  = 8'b00000000; // 5295 :   0 - 0x0
      13'h14B0: dout  = 8'b01000100; // 5296 :  68 - 0x44 -- Background 0x4b
      13'h14B1: dout  = 8'b01000100; // 5297 :  68 - 0x44
      13'h14B2: dout  = 8'b01001000; // 5298 :  72 - 0x48
      13'h14B3: dout  = 8'b01110000; // 5299 : 112 - 0x70
      13'h14B4: dout  = 8'b01001000; // 5300 :  72 - 0x48
      13'h14B5: dout  = 8'b00100100; // 5301 :  36 - 0x24
      13'h14B6: dout  = 8'b00100010; // 5302 :  34 - 0x22
      13'h14B7: dout  = 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout  = 8'b00000000; // 5304 :   0 - 0x0
      13'h14B9: dout  = 8'b00000000; // 5305 :   0 - 0x0
      13'h14BA: dout  = 8'b00000000; // 5306 :   0 - 0x0
      13'h14BB: dout  = 8'b00000000; // 5307 :   0 - 0x0
      13'h14BC: dout  = 8'b00000000; // 5308 :   0 - 0x0
      13'h14BD: dout  = 8'b00000000; // 5309 :   0 - 0x0
      13'h14BE: dout  = 8'b00000000; // 5310 :   0 - 0x0
      13'h14BF: dout  = 8'b00000000; // 5311 :   0 - 0x0
      13'h14C0: dout  = 8'b00010000; // 5312 :  16 - 0x10 -- Background 0x4c
      13'h14C1: dout  = 8'b00100000; // 5313 :  32 - 0x20
      13'h14C2: dout  = 8'b00100000; // 5314 :  32 - 0x20
      13'h14C3: dout  = 8'b00100000; // 5315 :  32 - 0x20
      13'h14C4: dout  = 8'b01000000; // 5316 :  64 - 0x40
      13'h14C5: dout  = 8'b01000000; // 5317 :  64 - 0x40
      13'h14C6: dout  = 8'b01000110; // 5318 :  70 - 0x46
      13'h14C7: dout  = 8'b00111000; // 5319 :  56 - 0x38
      13'h14C8: dout  = 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout  = 8'b00000000; // 5321 :   0 - 0x0
      13'h14CA: dout  = 8'b00000000; // 5322 :   0 - 0x0
      13'h14CB: dout  = 8'b00000000; // 5323 :   0 - 0x0
      13'h14CC: dout  = 8'b00000000; // 5324 :   0 - 0x0
      13'h14CD: dout  = 8'b00000000; // 5325 :   0 - 0x0
      13'h14CE: dout  = 8'b00000000; // 5326 :   0 - 0x0
      13'h14CF: dout  = 8'b00000000; // 5327 :   0 - 0x0
      13'h14D0: dout  = 8'b00100100; // 5328 :  36 - 0x24 -- Background 0x4d
      13'h14D1: dout  = 8'b01011010; // 5329 :  90 - 0x5a
      13'h14D2: dout  = 8'b01011010; // 5330 :  90 - 0x5a
      13'h14D3: dout  = 8'b01011010; // 5331 :  90 - 0x5a
      13'h14D4: dout  = 8'b01000010; // 5332 :  66 - 0x42
      13'h14D5: dout  = 8'b01000010; // 5333 :  66 - 0x42
      13'h14D6: dout  = 8'b00100010; // 5334 :  34 - 0x22
      13'h14D7: dout  = 8'b00000000; // 5335 :   0 - 0x0
      13'h14D8: dout  = 8'b00000000; // 5336 :   0 - 0x0
      13'h14D9: dout  = 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout  = 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout  = 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout  = 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout  = 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout  = 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout  = 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout  = 8'b00100100; // 5344 :  36 - 0x24 -- Background 0x4e
      13'h14E1: dout  = 8'b01010010; // 5345 :  82 - 0x52
      13'h14E2: dout  = 8'b01010010; // 5346 :  82 - 0x52
      13'h14E3: dout  = 8'b01010010; // 5347 :  82 - 0x52
      13'h14E4: dout  = 8'b01010010; // 5348 :  82 - 0x52
      13'h14E5: dout  = 8'b01010010; // 5349 :  82 - 0x52
      13'h14E6: dout  = 8'b01001100; // 5350 :  76 - 0x4c
      13'h14E7: dout  = 8'b00000000; // 5351 :   0 - 0x0
      13'h14E8: dout  = 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout  = 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout  = 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout  = 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout  = 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout  = 8'b00000000; // 5357 :   0 - 0x0
      13'h14EE: dout  = 8'b00000000; // 5358 :   0 - 0x0
      13'h14EF: dout  = 8'b00000000; // 5359 :   0 - 0x0
      13'h14F0: dout  = 8'b00111000; // 5360 :  56 - 0x38 -- Background 0x4f
      13'h14F1: dout  = 8'b01000100; // 5361 :  68 - 0x44
      13'h14F2: dout  = 8'b10000010; // 5362 : 130 - 0x82
      13'h14F3: dout  = 8'b10000010; // 5363 : 130 - 0x82
      13'h14F4: dout  = 8'b10000010; // 5364 : 130 - 0x82
      13'h14F5: dout  = 8'b01000100; // 5365 :  68 - 0x44
      13'h14F6: dout  = 8'b00111000; // 5366 :  56 - 0x38
      13'h14F7: dout  = 8'b00000000; // 5367 :   0 - 0x0
      13'h14F8: dout  = 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout  = 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout  = 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout  = 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout  = 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout  = 8'b00000000; // 5373 :   0 - 0x0
      13'h14FE: dout  = 8'b00000000; // 5374 :   0 - 0x0
      13'h14FF: dout  = 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout  = 8'b01111111; // 5376 : 127 - 0x7f -- Background 0x50
      13'h1501: dout  = 8'b11000000; // 5377 : 192 - 0xc0
      13'h1502: dout  = 8'b10000000; // 5378 : 128 - 0x80
      13'h1503: dout  = 8'b10000000; // 5379 : 128 - 0x80
      13'h1504: dout  = 8'b10000000; // 5380 : 128 - 0x80
      13'h1505: dout  = 8'b11000011; // 5381 : 195 - 0xc3
      13'h1506: dout  = 8'b11111111; // 5382 : 255 - 0xff
      13'h1507: dout  = 8'b11111111; // 5383 : 255 - 0xff
      13'h1508: dout  = 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout  = 8'b00111111; // 5385 :  63 - 0x3f
      13'h150A: dout  = 8'b01111111; // 5386 : 127 - 0x7f
      13'h150B: dout  = 8'b01111111; // 5387 : 127 - 0x7f
      13'h150C: dout  = 8'b01111111; // 5388 : 127 - 0x7f
      13'h150D: dout  = 8'b00111100; // 5389 :  60 - 0x3c
      13'h150E: dout  = 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout  = 8'b01000000; // 5391 :  64 - 0x40
      13'h1510: dout  = 8'b11111110; // 5392 : 254 - 0xfe -- Background 0x51
      13'h1511: dout  = 8'b00000011; // 5393 :   3 - 0x3
      13'h1512: dout  = 8'b00000001; // 5394 :   1 - 0x1
      13'h1513: dout  = 8'b00000001; // 5395 :   1 - 0x1
      13'h1514: dout  = 8'b00000001; // 5396 :   1 - 0x1
      13'h1515: dout  = 8'b11000011; // 5397 : 195 - 0xc3
      13'h1516: dout  = 8'b11111111; // 5398 : 255 - 0xff
      13'h1517: dout  = 8'b11111111; // 5399 : 255 - 0xff
      13'h1518: dout  = 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout  = 8'b11111100; // 5401 : 252 - 0xfc
      13'h151A: dout  = 8'b11111110; // 5402 : 254 - 0xfe
      13'h151B: dout  = 8'b11111110; // 5403 : 254 - 0xfe
      13'h151C: dout  = 8'b11111110; // 5404 : 254 - 0xfe
      13'h151D: dout  = 8'b00111100; // 5405 :  60 - 0x3c
      13'h151E: dout  = 8'b00000000; // 5406 :   0 - 0x0
      13'h151F: dout  = 8'b00000010; // 5407 :   2 - 0x2
      13'h1520: dout  = 8'b00000000; // 5408 :   0 - 0x0 -- Background 0x52
      13'h1521: dout  = 8'b00000111; // 5409 :   7 - 0x7
      13'h1522: dout  = 8'b00001100; // 5410 :  12 - 0xc
      13'h1523: dout  = 8'b00011000; // 5411 :  24 - 0x18
      13'h1524: dout  = 8'b00110000; // 5412 :  48 - 0x30
      13'h1525: dout  = 8'b01100000; // 5413 :  96 - 0x60
      13'h1526: dout  = 8'b01000000; // 5414 :  64 - 0x40
      13'h1527: dout  = 8'b01001111; // 5415 :  79 - 0x4f
      13'h1528: dout  = 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout  = 8'b00000000; // 5417 :   0 - 0x0
      13'h152A: dout  = 8'b00000011; // 5418 :   3 - 0x3
      13'h152B: dout  = 8'b00000111; // 5419 :   7 - 0x7
      13'h152C: dout  = 8'b00001111; // 5420 :  15 - 0xf
      13'h152D: dout  = 8'b00011111; // 5421 :  31 - 0x1f
      13'h152E: dout  = 8'b00111111; // 5422 :  63 - 0x3f
      13'h152F: dout  = 8'b00110000; // 5423 :  48 - 0x30
      13'h1530: dout  = 8'b00000000; // 5424 :   0 - 0x0 -- Background 0x53
      13'h1531: dout  = 8'b11110000; // 5425 : 240 - 0xf0
      13'h1532: dout  = 8'b01010000; // 5426 :  80 - 0x50
      13'h1533: dout  = 8'b01001000; // 5427 :  72 - 0x48
      13'h1534: dout  = 8'b01001100; // 5428 :  76 - 0x4c
      13'h1535: dout  = 8'b01000100; // 5429 :  68 - 0x44
      13'h1536: dout  = 8'b10000010; // 5430 : 130 - 0x82
      13'h1537: dout  = 8'b10000011; // 5431 : 131 - 0x83
      13'h1538: dout  = 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout  = 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout  = 8'b10100000; // 5434 : 160 - 0xa0
      13'h153B: dout  = 8'b10110000; // 5435 : 176 - 0xb0
      13'h153C: dout  = 8'b10110000; // 5436 : 176 - 0xb0
      13'h153D: dout  = 8'b10111000; // 5437 : 184 - 0xb8
      13'h153E: dout  = 8'b01111100; // 5438 : 124 - 0x7c
      13'h153F: dout  = 8'b01111100; // 5439 : 124 - 0x7c
      13'h1540: dout  = 8'b01111111; // 5440 : 127 - 0x7f -- Background 0x54
      13'h1541: dout  = 8'b11011110; // 5441 : 222 - 0xde
      13'h1542: dout  = 8'b10001110; // 5442 : 142 - 0x8e
      13'h1543: dout  = 8'b11000101; // 5443 : 197 - 0xc5
      13'h1544: dout  = 8'b10010010; // 5444 : 146 - 0x92
      13'h1545: dout  = 8'b11000111; // 5445 : 199 - 0xc7
      13'h1546: dout  = 8'b11100010; // 5446 : 226 - 0xe2
      13'h1547: dout  = 8'b11010000; // 5447 : 208 - 0xd0
      13'h1548: dout  = 8'b00000000; // 5448 :   0 - 0x0
      13'h1549: dout  = 8'b00100001; // 5449 :  33 - 0x21
      13'h154A: dout  = 8'b01110001; // 5450 : 113 - 0x71
      13'h154B: dout  = 8'b00111010; // 5451 :  58 - 0x3a
      13'h154C: dout  = 8'b01101101; // 5452 : 109 - 0x6d
      13'h154D: dout  = 8'b00111000; // 5453 :  56 - 0x38
      13'h154E: dout  = 8'b00011101; // 5454 :  29 - 0x1d
      13'h154F: dout  = 8'b00101111; // 5455 :  47 - 0x2f
      13'h1550: dout  = 8'b11111111; // 5456 : 255 - 0xff -- Background 0x55
      13'h1551: dout  = 8'b11011110; // 5457 : 222 - 0xde
      13'h1552: dout  = 8'b10001110; // 5458 : 142 - 0x8e
      13'h1553: dout  = 8'b11000101; // 5459 : 197 - 0xc5
      13'h1554: dout  = 8'b10010010; // 5460 : 146 - 0x92
      13'h1555: dout  = 8'b01000111; // 5461 :  71 - 0x47
      13'h1556: dout  = 8'b11100010; // 5462 : 226 - 0xe2
      13'h1557: dout  = 8'b01010000; // 5463 :  80 - 0x50
      13'h1558: dout  = 8'b00000000; // 5464 :   0 - 0x0
      13'h1559: dout  = 8'b00100001; // 5465 :  33 - 0x21
      13'h155A: dout  = 8'b01110001; // 5466 : 113 - 0x71
      13'h155B: dout  = 8'b00111010; // 5467 :  58 - 0x3a
      13'h155C: dout  = 8'b01101101; // 5468 : 109 - 0x6d
      13'h155D: dout  = 8'b10111000; // 5469 : 184 - 0xb8
      13'h155E: dout  = 8'b00011101; // 5470 :  29 - 0x1d
      13'h155F: dout  = 8'b10101111; // 5471 : 175 - 0xaf
      13'h1560: dout  = 8'b11111110; // 5472 : 254 - 0xfe -- Background 0x56
      13'h1561: dout  = 8'b11011111; // 5473 : 223 - 0xdf
      13'h1562: dout  = 8'b10001111; // 5474 : 143 - 0x8f
      13'h1563: dout  = 8'b11000101; // 5475 : 197 - 0xc5
      13'h1564: dout  = 8'b10010011; // 5476 : 147 - 0x93
      13'h1565: dout  = 8'b01000111; // 5477 :  71 - 0x47
      13'h1566: dout  = 8'b11100011; // 5478 : 227 - 0xe3
      13'h1567: dout  = 8'b01010001; // 5479 :  81 - 0x51
      13'h1568: dout  = 8'b00000000; // 5480 :   0 - 0x0
      13'h1569: dout  = 8'b00100000; // 5481 :  32 - 0x20
      13'h156A: dout  = 8'b01110000; // 5482 : 112 - 0x70
      13'h156B: dout  = 8'b00111010; // 5483 :  58 - 0x3a
      13'h156C: dout  = 8'b01101100; // 5484 : 108 - 0x6c
      13'h156D: dout  = 8'b10111000; // 5485 : 184 - 0xb8
      13'h156E: dout  = 8'b00011100; // 5486 :  28 - 0x1c
      13'h156F: dout  = 8'b10101110; // 5487 : 174 - 0xae
      13'h1570: dout  = 8'b01111111; // 5488 : 127 - 0x7f -- Background 0x57
      13'h1571: dout  = 8'b10000000; // 5489 : 128 - 0x80
      13'h1572: dout  = 8'b10110011; // 5490 : 179 - 0xb3
      13'h1573: dout  = 8'b01001100; // 5491 :  76 - 0x4c
      13'h1574: dout  = 8'b00111111; // 5492 :  63 - 0x3f
      13'h1575: dout  = 8'b00000011; // 5493 :   3 - 0x3
      13'h1576: dout  = 8'b00000000; // 5494 :   0 - 0x0
      13'h1577: dout  = 8'b00000000; // 5495 :   0 - 0x0
      13'h1578: dout  = 8'b00000000; // 5496 :   0 - 0x0
      13'h1579: dout  = 8'b01111111; // 5497 : 127 - 0x7f
      13'h157A: dout  = 8'b01001100; // 5498 :  76 - 0x4c
      13'h157B: dout  = 8'b00110011; // 5499 :  51 - 0x33
      13'h157C: dout  = 8'b00000000; // 5500 :   0 - 0x0
      13'h157D: dout  = 8'b00000000; // 5501 :   0 - 0x0
      13'h157E: dout  = 8'b00000000; // 5502 :   0 - 0x0
      13'h157F: dout  = 8'b00000000; // 5503 :   0 - 0x0
      13'h1580: dout  = 8'b11111111; // 5504 : 255 - 0xff -- Background 0x58
      13'h1581: dout  = 8'b00000000; // 5505 :   0 - 0x0
      13'h1582: dout  = 8'b00110011; // 5506 :  51 - 0x33
      13'h1583: dout  = 8'b11001100; // 5507 : 204 - 0xcc
      13'h1584: dout  = 8'b00110011; // 5508 :  51 - 0x33
      13'h1585: dout  = 8'b11111111; // 5509 : 255 - 0xff
      13'h1586: dout  = 8'b00000000; // 5510 :   0 - 0x0
      13'h1587: dout  = 8'b00000000; // 5511 :   0 - 0x0
      13'h1588: dout  = 8'b00000000; // 5512 :   0 - 0x0
      13'h1589: dout  = 8'b11111111; // 5513 : 255 - 0xff
      13'h158A: dout  = 8'b11001100; // 5514 : 204 - 0xcc
      13'h158B: dout  = 8'b00110011; // 5515 :  51 - 0x33
      13'h158C: dout  = 8'b11001100; // 5516 : 204 - 0xcc
      13'h158D: dout  = 8'b00000000; // 5517 :   0 - 0x0
      13'h158E: dout  = 8'b00000000; // 5518 :   0 - 0x0
      13'h158F: dout  = 8'b00000000; // 5519 :   0 - 0x0
      13'h1590: dout  = 8'b11111110; // 5520 : 254 - 0xfe -- Background 0x59
      13'h1591: dout  = 8'b00000001; // 5521 :   1 - 0x1
      13'h1592: dout  = 8'b00110011; // 5522 :  51 - 0x33
      13'h1593: dout  = 8'b11001110; // 5523 : 206 - 0xce
      13'h1594: dout  = 8'b00111100; // 5524 :  60 - 0x3c
      13'h1595: dout  = 8'b11000000; // 5525 : 192 - 0xc0
      13'h1596: dout  = 8'b00000000; // 5526 :   0 - 0x0
      13'h1597: dout  = 8'b00000000; // 5527 :   0 - 0x0
      13'h1598: dout  = 8'b00000000; // 5528 :   0 - 0x0
      13'h1599: dout  = 8'b11111110; // 5529 : 254 - 0xfe
      13'h159A: dout  = 8'b11001100; // 5530 : 204 - 0xcc
      13'h159B: dout  = 8'b00110000; // 5531 :  48 - 0x30
      13'h159C: dout  = 8'b11000000; // 5532 : 192 - 0xc0
      13'h159D: dout  = 8'b00000000; // 5533 :   0 - 0x0
      13'h159E: dout  = 8'b00000000; // 5534 :   0 - 0x0
      13'h159F: dout  = 8'b00000000; // 5535 :   0 - 0x0
      13'h15A0: dout  = 8'b00000000; // 5536 :   0 - 0x0 -- Background 0x5a
      13'h15A1: dout  = 8'b00000000; // 5537 :   0 - 0x0
      13'h15A2: dout  = 8'b00000000; // 5538 :   0 - 0x0
      13'h15A3: dout  = 8'b00000000; // 5539 :   0 - 0x0
      13'h15A4: dout  = 8'b00000000; // 5540 :   0 - 0x0
      13'h15A5: dout  = 8'b00000000; // 5541 :   0 - 0x0
      13'h15A6: dout  = 8'b00000000; // 5542 :   0 - 0x0
      13'h15A7: dout  = 8'b00000000; // 5543 :   0 - 0x0
      13'h15A8: dout  = 8'b00000000; // 5544 :   0 - 0x0
      13'h15A9: dout  = 8'b00000000; // 5545 :   0 - 0x0
      13'h15AA: dout  = 8'b00000000; // 5546 :   0 - 0x0
      13'h15AB: dout  = 8'b00000000; // 5547 :   0 - 0x0
      13'h15AC: dout  = 8'b00000000; // 5548 :   0 - 0x0
      13'h15AD: dout  = 8'b00000000; // 5549 :   0 - 0x0
      13'h15AE: dout  = 8'b00000000; // 5550 :   0 - 0x0
      13'h15AF: dout  = 8'b00000000; // 5551 :   0 - 0x0
      13'h15B0: dout  = 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout  = 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout  = 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout  = 8'b00000001; // 5555 :   1 - 0x1
      13'h15B4: dout  = 8'b00000011; // 5556 :   3 - 0x3
      13'h15B5: dout  = 8'b00000011; // 5557 :   3 - 0x3
      13'h15B6: dout  = 8'b00000111; // 5558 :   7 - 0x7
      13'h15B7: dout  = 8'b00111111; // 5559 :  63 - 0x3f
      13'h15B8: dout  = 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout  = 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout  = 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout  = 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout  = 8'b00000001; // 5564 :   1 - 0x1
      13'h15BD: dout  = 8'b00000001; // 5565 :   1 - 0x1
      13'h15BE: dout  = 8'b00000011; // 5566 :   3 - 0x3
      13'h15BF: dout  = 8'b00000011; // 5567 :   3 - 0x3
      13'h15C0: dout  = 8'b00000000; // 5568 :   0 - 0x0 -- Background 0x5c
      13'h15C1: dout  = 8'b00000001; // 5569 :   1 - 0x1
      13'h15C2: dout  = 8'b01111111; // 5570 : 127 - 0x7f
      13'h15C3: dout  = 8'b11111111; // 5571 : 255 - 0xff
      13'h15C4: dout  = 8'b11111111; // 5572 : 255 - 0xff
      13'h15C5: dout  = 8'b11111111; // 5573 : 255 - 0xff
      13'h15C6: dout  = 8'b11111111; // 5574 : 255 - 0xff
      13'h15C7: dout  = 8'b11111111; // 5575 : 255 - 0xff
      13'h15C8: dout  = 8'b00000000; // 5576 :   0 - 0x0
      13'h15C9: dout  = 8'b00000000; // 5577 :   0 - 0x0
      13'h15CA: dout  = 8'b00000001; // 5578 :   1 - 0x1
      13'h15CB: dout  = 8'b01111110; // 5579 : 126 - 0x7e
      13'h15CC: dout  = 8'b11111111; // 5580 : 255 - 0xff
      13'h15CD: dout  = 8'b11111111; // 5581 : 255 - 0xff
      13'h15CE: dout  = 8'b11111111; // 5582 : 255 - 0xff
      13'h15CF: dout  = 8'b11111111; // 5583 : 255 - 0xff
      13'h15D0: dout  = 8'b11111111; // 5584 : 255 - 0xff -- Background 0x5d
      13'h15D1: dout  = 8'b11111111; // 5585 : 255 - 0xff
      13'h15D2: dout  = 8'b11111111; // 5586 : 255 - 0xff
      13'h15D3: dout  = 8'b11111111; // 5587 : 255 - 0xff
      13'h15D4: dout  = 8'b11111111; // 5588 : 255 - 0xff
      13'h15D5: dout  = 8'b11111111; // 5589 : 255 - 0xff
      13'h15D6: dout  = 8'b11111111; // 5590 : 255 - 0xff
      13'h15D7: dout  = 8'b11111111; // 5591 : 255 - 0xff
      13'h15D8: dout  = 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout  = 8'b11111111; // 5593 : 255 - 0xff
      13'h15DA: dout  = 8'b11111111; // 5594 : 255 - 0xff
      13'h15DB: dout  = 8'b11111111; // 5595 : 255 - 0xff
      13'h15DC: dout  = 8'b01111111; // 5596 : 127 - 0x7f
      13'h15DD: dout  = 8'b11111111; // 5597 : 255 - 0xff
      13'h15DE: dout  = 8'b11111111; // 5598 : 255 - 0xff
      13'h15DF: dout  = 8'b11111111; // 5599 : 255 - 0xff
      13'h15E0: dout  = 8'b00000000; // 5600 :   0 - 0x0 -- Background 0x5e
      13'h15E1: dout  = 8'b10000000; // 5601 : 128 - 0x80
      13'h15E2: dout  = 8'b11111110; // 5602 : 254 - 0xfe
      13'h15E3: dout  = 8'b11111111; // 5603 : 255 - 0xff
      13'h15E4: dout  = 8'b11111111; // 5604 : 255 - 0xff
      13'h15E5: dout  = 8'b11111111; // 5605 : 255 - 0xff
      13'h15E6: dout  = 8'b11111111; // 5606 : 255 - 0xff
      13'h15E7: dout  = 8'b11111111; // 5607 : 255 - 0xff
      13'h15E8: dout  = 8'b00000000; // 5608 :   0 - 0x0
      13'h15E9: dout  = 8'b00000000; // 5609 :   0 - 0x0
      13'h15EA: dout  = 8'b10000000; // 5610 : 128 - 0x80
      13'h15EB: dout  = 8'b01111110; // 5611 : 126 - 0x7e
      13'h15EC: dout  = 8'b10111111; // 5612 : 191 - 0xbf
      13'h15ED: dout  = 8'b11111111; // 5613 : 255 - 0xff
      13'h15EE: dout  = 8'b11111111; // 5614 : 255 - 0xff
      13'h15EF: dout  = 8'b11111111; // 5615 : 255 - 0xff
      13'h15F0: dout  = 8'b00000000; // 5616 :   0 - 0x0 -- Background 0x5f
      13'h15F1: dout  = 8'b00000000; // 5617 :   0 - 0x0
      13'h15F2: dout  = 8'b00000000; // 5618 :   0 - 0x0
      13'h15F3: dout  = 8'b10000000; // 5619 : 128 - 0x80
      13'h15F4: dout  = 8'b11000000; // 5620 : 192 - 0xc0
      13'h15F5: dout  = 8'b11000000; // 5621 : 192 - 0xc0
      13'h15F6: dout  = 8'b11100000; // 5622 : 224 - 0xe0
      13'h15F7: dout  = 8'b11111000; // 5623 : 248 - 0xf8
      13'h15F8: dout  = 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout  = 8'b00000000; // 5625 :   0 - 0x0
      13'h15FA: dout  = 8'b00000000; // 5626 :   0 - 0x0
      13'h15FB: dout  = 8'b00000000; // 5627 :   0 - 0x0
      13'h15FC: dout  = 8'b10000000; // 5628 : 128 - 0x80
      13'h15FD: dout  = 8'b10000000; // 5629 : 128 - 0x80
      13'h15FE: dout  = 8'b11000000; // 5630 : 192 - 0xc0
      13'h15FF: dout  = 8'b11000000; // 5631 : 192 - 0xc0
      13'h1600: dout  = 8'b11111111; // 5632 : 255 - 0xff -- Background 0x60
      13'h1601: dout  = 8'b11111111; // 5633 : 255 - 0xff
      13'h1602: dout  = 8'b11111111; // 5634 : 255 - 0xff
      13'h1603: dout  = 8'b11111111; // 5635 : 255 - 0xff
      13'h1604: dout  = 8'b11111111; // 5636 : 255 - 0xff
      13'h1605: dout  = 8'b11111111; // 5637 : 255 - 0xff
      13'h1606: dout  = 8'b11111111; // 5638 : 255 - 0xff
      13'h1607: dout  = 8'b11111111; // 5639 : 255 - 0xff
      13'h1608: dout  = 8'b01111111; // 5640 : 127 - 0x7f
      13'h1609: dout  = 8'b01111111; // 5641 : 127 - 0x7f
      13'h160A: dout  = 8'b01111101; // 5642 : 125 - 0x7d
      13'h160B: dout  = 8'b01111111; // 5643 : 127 - 0x7f
      13'h160C: dout  = 8'b00111111; // 5644 :  63 - 0x3f
      13'h160D: dout  = 8'b01111111; // 5645 : 127 - 0x7f
      13'h160E: dout  = 8'b01111111; // 5646 : 127 - 0x7f
      13'h160F: dout  = 8'b01110111; // 5647 : 119 - 0x77
      13'h1610: dout  = 8'b11111111; // 5648 : 255 - 0xff -- Background 0x61
      13'h1611: dout  = 8'b11111111; // 5649 : 255 - 0xff
      13'h1612: dout  = 8'b11111111; // 5650 : 255 - 0xff
      13'h1613: dout  = 8'b11111111; // 5651 : 255 - 0xff
      13'h1614: dout  = 8'b11111111; // 5652 : 255 - 0xff
      13'h1615: dout  = 8'b11111111; // 5653 : 255 - 0xff
      13'h1616: dout  = 8'b11111111; // 5654 : 255 - 0xff
      13'h1617: dout  = 8'b11111111; // 5655 : 255 - 0xff
      13'h1618: dout  = 8'b11111110; // 5656 : 254 - 0xfe
      13'h1619: dout  = 8'b11111110; // 5657 : 254 - 0xfe
      13'h161A: dout  = 8'b11111100; // 5658 : 252 - 0xfc
      13'h161B: dout  = 8'b11111110; // 5659 : 254 - 0xfe
      13'h161C: dout  = 8'b10111110; // 5660 : 190 - 0xbe
      13'h161D: dout  = 8'b11111110; // 5661 : 254 - 0xfe
      13'h161E: dout  = 8'b11111110; // 5662 : 254 - 0xfe
      13'h161F: dout  = 8'b11110110; // 5663 : 246 - 0xf6
      13'h1620: dout  = 8'b01111000; // 5664 : 120 - 0x78 -- Background 0x62
      13'h1621: dout  = 8'b01100000; // 5665 :  96 - 0x60
      13'h1622: dout  = 8'b01000000; // 5666 :  64 - 0x40
      13'h1623: dout  = 8'b01000000; // 5667 :  64 - 0x40
      13'h1624: dout  = 8'b01000000; // 5668 :  64 - 0x40
      13'h1625: dout  = 8'b01100000; // 5669 :  96 - 0x60
      13'h1626: dout  = 8'b00110000; // 5670 :  48 - 0x30
      13'h1627: dout  = 8'b00011111; // 5671 :  31 - 0x1f
      13'h1628: dout  = 8'b00000111; // 5672 :   7 - 0x7
      13'h1629: dout  = 8'b00011111; // 5673 :  31 - 0x1f
      13'h162A: dout  = 8'b00111111; // 5674 :  63 - 0x3f
      13'h162B: dout  = 8'b00111111; // 5675 :  63 - 0x3f
      13'h162C: dout  = 8'b00111111; // 5676 :  63 - 0x3f
      13'h162D: dout  = 8'b00011111; // 5677 :  31 - 0x1f
      13'h162E: dout  = 8'b00001111; // 5678 :  15 - 0xf
      13'h162F: dout  = 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout  = 8'b10000001; // 5680 : 129 - 0x81 -- Background 0x63
      13'h1631: dout  = 8'b10000011; // 5681 : 131 - 0x83
      13'h1632: dout  = 8'b11000001; // 5682 : 193 - 0xc1
      13'h1633: dout  = 8'b01000011; // 5683 :  67 - 0x43
      13'h1634: dout  = 8'b01000001; // 5684 :  65 - 0x41
      13'h1635: dout  = 8'b01100011; // 5685 :  99 - 0x63
      13'h1636: dout  = 8'b00100110; // 5686 :  38 - 0x26
      13'h1637: dout  = 8'b11111000; // 5687 : 248 - 0xf8
      13'h1638: dout  = 8'b01111110; // 5688 : 126 - 0x7e
      13'h1639: dout  = 8'b01111100; // 5689 : 124 - 0x7c
      13'h163A: dout  = 8'b00111110; // 5690 :  62 - 0x3e
      13'h163B: dout  = 8'b10111100; // 5691 : 188 - 0xbc
      13'h163C: dout  = 8'b10111110; // 5692 : 190 - 0xbe
      13'h163D: dout  = 8'b10011100; // 5693 : 156 - 0x9c
      13'h163E: dout  = 8'b11011000; // 5694 : 216 - 0xd8
      13'h163F: dout  = 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout  = 8'b10111001; // 5696 : 185 - 0xb9 -- Background 0x64
      13'h1641: dout  = 8'b10010100; // 5697 : 148 - 0x94
      13'h1642: dout  = 8'b10001110; // 5698 : 142 - 0x8e
      13'h1643: dout  = 8'b11000101; // 5699 : 197 - 0xc5
      13'h1644: dout  = 8'b10010010; // 5700 : 146 - 0x92
      13'h1645: dout  = 8'b11000111; // 5701 : 199 - 0xc7
      13'h1646: dout  = 8'b11100010; // 5702 : 226 - 0xe2
      13'h1647: dout  = 8'b11010000; // 5703 : 208 - 0xd0
      13'h1648: dout  = 8'b01000110; // 5704 :  70 - 0x46
      13'h1649: dout  = 8'b01101011; // 5705 : 107 - 0x6b
      13'h164A: dout  = 8'b01110001; // 5706 : 113 - 0x71
      13'h164B: dout  = 8'b00111010; // 5707 :  58 - 0x3a
      13'h164C: dout  = 8'b01101101; // 5708 : 109 - 0x6d
      13'h164D: dout  = 8'b00111000; // 5709 :  56 - 0x38
      13'h164E: dout  = 8'b00011101; // 5710 :  29 - 0x1d
      13'h164F: dout  = 8'b00101111; // 5711 :  47 - 0x2f
      13'h1650: dout  = 8'b10111001; // 5712 : 185 - 0xb9 -- Background 0x65
      13'h1651: dout  = 8'b00010100; // 5713 :  20 - 0x14
      13'h1652: dout  = 8'b10001110; // 5714 : 142 - 0x8e
      13'h1653: dout  = 8'b11000101; // 5715 : 197 - 0xc5
      13'h1654: dout  = 8'b10010010; // 5716 : 146 - 0x92
      13'h1655: dout  = 8'b01000111; // 5717 :  71 - 0x47
      13'h1656: dout  = 8'b11100010; // 5718 : 226 - 0xe2
      13'h1657: dout  = 8'b01010000; // 5719 :  80 - 0x50
      13'h1658: dout  = 8'b01000110; // 5720 :  70 - 0x46
      13'h1659: dout  = 8'b11101011; // 5721 : 235 - 0xeb
      13'h165A: dout  = 8'b01110001; // 5722 : 113 - 0x71
      13'h165B: dout  = 8'b00111010; // 5723 :  58 - 0x3a
      13'h165C: dout  = 8'b01101101; // 5724 : 109 - 0x6d
      13'h165D: dout  = 8'b10111000; // 5725 : 184 - 0xb8
      13'h165E: dout  = 8'b00011101; // 5726 :  29 - 0x1d
      13'h165F: dout  = 8'b10101111; // 5727 : 175 - 0xaf
      13'h1660: dout  = 8'b10111001; // 5728 : 185 - 0xb9 -- Background 0x66
      13'h1661: dout  = 8'b00010101; // 5729 :  21 - 0x15
      13'h1662: dout  = 8'b10001111; // 5730 : 143 - 0x8f
      13'h1663: dout  = 8'b11000101; // 5731 : 197 - 0xc5
      13'h1664: dout  = 8'b10010011; // 5732 : 147 - 0x93
      13'h1665: dout  = 8'b01000111; // 5733 :  71 - 0x47
      13'h1666: dout  = 8'b11100011; // 5734 : 227 - 0xe3
      13'h1667: dout  = 8'b01010001; // 5735 :  81 - 0x51
      13'h1668: dout  = 8'b01000110; // 5736 :  70 - 0x46
      13'h1669: dout  = 8'b11101010; // 5737 : 234 - 0xea
      13'h166A: dout  = 8'b01110000; // 5738 : 112 - 0x70
      13'h166B: dout  = 8'b00111010; // 5739 :  58 - 0x3a
      13'h166C: dout  = 8'b01101100; // 5740 : 108 - 0x6c
      13'h166D: dout  = 8'b10111000; // 5741 : 184 - 0xb8
      13'h166E: dout  = 8'b00011100; // 5742 :  28 - 0x1c
      13'h166F: dout  = 8'b10101110; // 5743 : 174 - 0xae
      13'h1670: dout  = 8'b01111111; // 5744 : 127 - 0x7f -- Background 0x67
      13'h1671: dout  = 8'b10000000; // 5745 : 128 - 0x80
      13'h1672: dout  = 8'b11001100; // 5746 : 204 - 0xcc
      13'h1673: dout  = 8'b01111111; // 5747 : 127 - 0x7f
      13'h1674: dout  = 8'b00111111; // 5748 :  63 - 0x3f
      13'h1675: dout  = 8'b00000011; // 5749 :   3 - 0x3
      13'h1676: dout  = 8'b00000000; // 5750 :   0 - 0x0
      13'h1677: dout  = 8'b00000000; // 5751 :   0 - 0x0
      13'h1678: dout  = 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout  = 8'b01111111; // 5753 : 127 - 0x7f
      13'h167A: dout  = 8'b01111111; // 5754 : 127 - 0x7f
      13'h167B: dout  = 8'b00110011; // 5755 :  51 - 0x33
      13'h167C: dout  = 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout  = 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout  = 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout  = 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout  = 8'b11111111; // 5760 : 255 - 0xff -- Background 0x68
      13'h1681: dout  = 8'b00000000; // 5761 :   0 - 0x0
      13'h1682: dout  = 8'b11001100; // 5762 : 204 - 0xcc
      13'h1683: dout  = 8'b00110011; // 5763 :  51 - 0x33
      13'h1684: dout  = 8'b11111111; // 5764 : 255 - 0xff
      13'h1685: dout  = 8'b11111111; // 5765 : 255 - 0xff
      13'h1686: dout  = 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout  = 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout  = 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout  = 8'b11111111; // 5769 : 255 - 0xff
      13'h168A: dout  = 8'b11111111; // 5770 : 255 - 0xff
      13'h168B: dout  = 8'b11111111; // 5771 : 255 - 0xff
      13'h168C: dout  = 8'b11001100; // 5772 : 204 - 0xcc
      13'h168D: dout  = 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout  = 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout  = 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout  = 8'b11111110; // 5776 : 254 - 0xfe -- Background 0x69
      13'h1691: dout  = 8'b00000001; // 5777 :   1 - 0x1
      13'h1692: dout  = 8'b11001101; // 5778 : 205 - 0xcd
      13'h1693: dout  = 8'b00111110; // 5779 :  62 - 0x3e
      13'h1694: dout  = 8'b11111100; // 5780 : 252 - 0xfc
      13'h1695: dout  = 8'b11000000; // 5781 : 192 - 0xc0
      13'h1696: dout  = 8'b00000000; // 5782 :   0 - 0x0
      13'h1697: dout  = 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout  = 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout  = 8'b11111110; // 5785 : 254 - 0xfe
      13'h169A: dout  = 8'b11111110; // 5786 : 254 - 0xfe
      13'h169B: dout  = 8'b11110000; // 5787 : 240 - 0xf0
      13'h169C: dout  = 8'b11000000; // 5788 : 192 - 0xc0
      13'h169D: dout  = 8'b00000000; // 5789 :   0 - 0x0
      13'h169E: dout  = 8'b00000000; // 5790 :   0 - 0x0
      13'h169F: dout  = 8'b00000000; // 5791 :   0 - 0x0
      13'h16A0: dout  = 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout  = 8'b00000000; // 5793 :   0 - 0x0
      13'h16A2: dout  = 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout  = 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout  = 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout  = 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout  = 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout  = 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout  = 8'b00000000; // 5800 :   0 - 0x0
      13'h16A9: dout  = 8'b00000000; // 5801 :   0 - 0x0
      13'h16AA: dout  = 8'b00000000; // 5802 :   0 - 0x0
      13'h16AB: dout  = 8'b00000000; // 5803 :   0 - 0x0
      13'h16AC: dout  = 8'b00000000; // 5804 :   0 - 0x0
      13'h16AD: dout  = 8'b00000000; // 5805 :   0 - 0x0
      13'h16AE: dout  = 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout  = 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout  = 8'b01111111; // 5808 : 127 - 0x7f -- Background 0x6b
      13'h16B1: dout  = 8'b11111111; // 5809 : 255 - 0xff
      13'h16B2: dout  = 8'b11111111; // 5810 : 255 - 0xff
      13'h16B3: dout  = 8'b11111111; // 5811 : 255 - 0xff
      13'h16B4: dout  = 8'b01111111; // 5812 : 127 - 0x7f
      13'h16B5: dout  = 8'b00110000; // 5813 :  48 - 0x30
      13'h16B6: dout  = 8'b00001111; // 5814 :  15 - 0xf
      13'h16B7: dout  = 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout  = 8'b00111101; // 5816 :  61 - 0x3d
      13'h16B9: dout  = 8'b01111111; // 5817 : 127 - 0x7f
      13'h16BA: dout  = 8'b01111111; // 5818 : 127 - 0x7f
      13'h16BB: dout  = 8'b01111111; // 5819 : 127 - 0x7f
      13'h16BC: dout  = 8'b00111111; // 5820 :  63 - 0x3f
      13'h16BD: dout  = 8'b00001111; // 5821 :  15 - 0xf
      13'h16BE: dout  = 8'b00000000; // 5822 :   0 - 0x0
      13'h16BF: dout  = 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout  = 8'b11111111; // 5824 : 255 - 0xff -- Background 0x6c
      13'h16C1: dout  = 8'b11111111; // 5825 : 255 - 0xff
      13'h16C2: dout  = 8'b11111111; // 5826 : 255 - 0xff
      13'h16C3: dout  = 8'b11111111; // 5827 : 255 - 0xff
      13'h16C4: dout  = 8'b11111111; // 5828 : 255 - 0xff
      13'h16C5: dout  = 8'b11111110; // 5829 : 254 - 0xfe
      13'h16C6: dout  = 8'b00000001; // 5830 :   1 - 0x1
      13'h16C7: dout  = 8'b11111110; // 5831 : 254 - 0xfe
      13'h16C8: dout  = 8'b11111111; // 5832 : 255 - 0xff
      13'h16C9: dout  = 8'b11111111; // 5833 : 255 - 0xff
      13'h16CA: dout  = 8'b11111111; // 5834 : 255 - 0xff
      13'h16CB: dout  = 8'b11111111; // 5835 : 255 - 0xff
      13'h16CC: dout  = 8'b11111111; // 5836 : 255 - 0xff
      13'h16CD: dout  = 8'b11111111; // 5837 : 255 - 0xff
      13'h16CE: dout  = 8'b11111110; // 5838 : 254 - 0xfe
      13'h16CF: dout  = 8'b00000000; // 5839 :   0 - 0x0
      13'h16D0: dout  = 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout  = 8'b00000000; // 5841 :   0 - 0x0
      13'h16D2: dout  = 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout  = 8'b00000000; // 5843 :   0 - 0x0
      13'h16D4: dout  = 8'b00000000; // 5844 :   0 - 0x0
      13'h16D5: dout  = 8'b00000000; // 5845 :   0 - 0x0
      13'h16D6: dout  = 8'b00000000; // 5846 :   0 - 0x0
      13'h16D7: dout  = 8'b00000000; // 5847 :   0 - 0x0
      13'h16D8: dout  = 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout  = 8'b00000000; // 5849 :   0 - 0x0
      13'h16DA: dout  = 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout  = 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout  = 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout  = 8'b00000000; // 5853 :   0 - 0x0
      13'h16DE: dout  = 8'b00000000; // 5854 :   0 - 0x0
      13'h16DF: dout  = 8'b00000000; // 5855 :   0 - 0x0
      13'h16E0: dout  = 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout  = 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout  = 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout  = 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout  = 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout  = 8'b00000000; // 5861 :   0 - 0x0
      13'h16E6: dout  = 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout  = 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout  = 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout  = 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout  = 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout  = 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout  = 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout  = 8'b00000000; // 5869 :   0 - 0x0
      13'h16EE: dout  = 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout  = 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout  = 8'b11111100; // 5872 : 252 - 0xfc -- Background 0x6f
      13'h16F1: dout  = 8'b11111110; // 5873 : 254 - 0xfe
      13'h16F2: dout  = 8'b11111111; // 5874 : 255 - 0xff
      13'h16F3: dout  = 8'b11111111; // 5875 : 255 - 0xff
      13'h16F4: dout  = 8'b11110010; // 5876 : 242 - 0xf2
      13'h16F5: dout  = 8'b00001100; // 5877 :  12 - 0xc
      13'h16F6: dout  = 8'b11110000; // 5878 : 240 - 0xf0
      13'h16F7: dout  = 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout  = 8'b10111000; // 5880 : 184 - 0xb8
      13'h16F9: dout  = 8'b11111100; // 5881 : 252 - 0xfc
      13'h16FA: dout  = 8'b11111110; // 5882 : 254 - 0xfe
      13'h16FB: dout  = 8'b11111110; // 5883 : 254 - 0xfe
      13'h16FC: dout  = 8'b11111100; // 5884 : 252 - 0xfc
      13'h16FD: dout  = 8'b11110000; // 5885 : 240 - 0xf0
      13'h16FE: dout  = 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout  = 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout  = 8'b01111111; // 5888 : 127 - 0x7f -- Background 0x70
      13'h1701: dout  = 8'b11000000; // 5889 : 192 - 0xc0
      13'h1702: dout  = 8'b10000000; // 5890 : 128 - 0x80
      13'h1703: dout  = 8'b10000000; // 5891 : 128 - 0x80
      13'h1704: dout  = 8'b11100011; // 5892 : 227 - 0xe3
      13'h1705: dout  = 8'b11111111; // 5893 : 255 - 0xff
      13'h1706: dout  = 8'b11111111; // 5894 : 255 - 0xff
      13'h1707: dout  = 8'b11111111; // 5895 : 255 - 0xff
      13'h1708: dout  = 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout  = 8'b00111111; // 5897 :  63 - 0x3f
      13'h170A: dout  = 8'b01111111; // 5898 : 127 - 0x7f
      13'h170B: dout  = 8'b01111111; // 5899 : 127 - 0x7f
      13'h170C: dout  = 8'b00011100; // 5900 :  28 - 0x1c
      13'h170D: dout  = 8'b00000000; // 5901 :   0 - 0x0
      13'h170E: dout  = 8'b00000000; // 5902 :   0 - 0x0
      13'h170F: dout  = 8'b00000000; // 5903 :   0 - 0x0
      13'h1710: dout  = 8'b11111111; // 5904 : 255 - 0xff -- Background 0x71
      13'h1711: dout  = 8'b00000000; // 5905 :   0 - 0x0
      13'h1712: dout  = 8'b00000000; // 5906 :   0 - 0x0
      13'h1713: dout  = 8'b00000000; // 5907 :   0 - 0x0
      13'h1714: dout  = 8'b00000000; // 5908 :   0 - 0x0
      13'h1715: dout  = 8'b11000011; // 5909 : 195 - 0xc3
      13'h1716: dout  = 8'b11111111; // 5910 : 255 - 0xff
      13'h1717: dout  = 8'b11111111; // 5911 : 255 - 0xff
      13'h1718: dout  = 8'b00000000; // 5912 :   0 - 0x0
      13'h1719: dout  = 8'b11111111; // 5913 : 255 - 0xff
      13'h171A: dout  = 8'b11111111; // 5914 : 255 - 0xff
      13'h171B: dout  = 8'b11111111; // 5915 : 255 - 0xff
      13'h171C: dout  = 8'b11111111; // 5916 : 255 - 0xff
      13'h171D: dout  = 8'b00111100; // 5917 :  60 - 0x3c
      13'h171E: dout  = 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout  = 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout  = 8'b11111110; // 5920 : 254 - 0xfe -- Background 0x72
      13'h1721: dout  = 8'b00000011; // 5921 :   3 - 0x3
      13'h1722: dout  = 8'b00000001; // 5922 :   1 - 0x1
      13'h1723: dout  = 8'b00000001; // 5923 :   1 - 0x1
      13'h1724: dout  = 8'b11000111; // 5924 : 199 - 0xc7
      13'h1725: dout  = 8'b11111111; // 5925 : 255 - 0xff
      13'h1726: dout  = 8'b11111111; // 5926 : 255 - 0xff
      13'h1727: dout  = 8'b11111111; // 5927 : 255 - 0xff
      13'h1728: dout  = 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout  = 8'b11111100; // 5929 : 252 - 0xfc
      13'h172A: dout  = 8'b11111110; // 5930 : 254 - 0xfe
      13'h172B: dout  = 8'b11111110; // 5931 : 254 - 0xfe
      13'h172C: dout  = 8'b00111000; // 5932 :  56 - 0x38
      13'h172D: dout  = 8'b00000000; // 5933 :   0 - 0x0
      13'h172E: dout  = 8'b00000000; // 5934 :   0 - 0x0
      13'h172F: dout  = 8'b00000000; // 5935 :   0 - 0x0
      13'h1730: dout  = 8'b11111111; // 5936 : 255 - 0xff -- Background 0x73
      13'h1731: dout  = 8'b11111111; // 5937 : 255 - 0xff
      13'h1732: dout  = 8'b11111111; // 5938 : 255 - 0xff
      13'h1733: dout  = 8'b11111111; // 5939 : 255 - 0xff
      13'h1734: dout  = 8'b11111111; // 5940 : 255 - 0xff
      13'h1735: dout  = 8'b11111111; // 5941 : 255 - 0xff
      13'h1736: dout  = 8'b11111111; // 5942 : 255 - 0xff
      13'h1737: dout  = 8'b11111111; // 5943 : 255 - 0xff
      13'h1738: dout  = 8'b11111111; // 5944 : 255 - 0xff
      13'h1739: dout  = 8'b11111111; // 5945 : 255 - 0xff
      13'h173A: dout  = 8'b11111101; // 5946 : 253 - 0xfd
      13'h173B: dout  = 8'b11111111; // 5947 : 255 - 0xff
      13'h173C: dout  = 8'b10111111; // 5948 : 191 - 0xbf
      13'h173D: dout  = 8'b11111111; // 5949 : 255 - 0xff
      13'h173E: dout  = 8'b11111111; // 5950 : 255 - 0xff
      13'h173F: dout  = 8'b11110111; // 5951 : 247 - 0xf7
      13'h1740: dout  = 8'b10111001; // 5952 : 185 - 0xb9 -- Background 0x74
      13'h1741: dout  = 8'b10010100; // 5953 : 148 - 0x94
      13'h1742: dout  = 8'b10001110; // 5954 : 142 - 0x8e
      13'h1743: dout  = 8'b11000101; // 5955 : 197 - 0xc5
      13'h1744: dout  = 8'b10010010; // 5956 : 146 - 0x92
      13'h1745: dout  = 8'b11000111; // 5957 : 199 - 0xc7
      13'h1746: dout  = 8'b11100010; // 5958 : 226 - 0xe2
      13'h1747: dout  = 8'b01111111; // 5959 : 127 - 0x7f
      13'h1748: dout  = 8'b01000110; // 5960 :  70 - 0x46
      13'h1749: dout  = 8'b01101011; // 5961 : 107 - 0x6b
      13'h174A: dout  = 8'b01110001; // 5962 : 113 - 0x71
      13'h174B: dout  = 8'b00111010; // 5963 :  58 - 0x3a
      13'h174C: dout  = 8'b01101101; // 5964 : 109 - 0x6d
      13'h174D: dout  = 8'b00111000; // 5965 :  56 - 0x38
      13'h174E: dout  = 8'b00011101; // 5966 :  29 - 0x1d
      13'h174F: dout  = 8'b00000000; // 5967 :   0 - 0x0
      13'h1750: dout  = 8'b10111001; // 5968 : 185 - 0xb9 -- Background 0x75
      13'h1751: dout  = 8'b00010100; // 5969 :  20 - 0x14
      13'h1752: dout  = 8'b10001110; // 5970 : 142 - 0x8e
      13'h1753: dout  = 8'b11000101; // 5971 : 197 - 0xc5
      13'h1754: dout  = 8'b10010010; // 5972 : 146 - 0x92
      13'h1755: dout  = 8'b01000111; // 5973 :  71 - 0x47
      13'h1756: dout  = 8'b11100010; // 5974 : 226 - 0xe2
      13'h1757: dout  = 8'b11111111; // 5975 : 255 - 0xff
      13'h1758: dout  = 8'b01000110; // 5976 :  70 - 0x46
      13'h1759: dout  = 8'b11101011; // 5977 : 235 - 0xeb
      13'h175A: dout  = 8'b01110001; // 5978 : 113 - 0x71
      13'h175B: dout  = 8'b00111010; // 5979 :  58 - 0x3a
      13'h175C: dout  = 8'b01101101; // 5980 : 109 - 0x6d
      13'h175D: dout  = 8'b10111000; // 5981 : 184 - 0xb8
      13'h175E: dout  = 8'b00011101; // 5982 :  29 - 0x1d
      13'h175F: dout  = 8'b00000000; // 5983 :   0 - 0x0
      13'h1760: dout  = 8'b10111001; // 5984 : 185 - 0xb9 -- Background 0x76
      13'h1761: dout  = 8'b00010101; // 5985 :  21 - 0x15
      13'h1762: dout  = 8'b10001111; // 5986 : 143 - 0x8f
      13'h1763: dout  = 8'b11000101; // 5987 : 197 - 0xc5
      13'h1764: dout  = 8'b10010011; // 5988 : 147 - 0x93
      13'h1765: dout  = 8'b01000111; // 5989 :  71 - 0x47
      13'h1766: dout  = 8'b11100011; // 5990 : 227 - 0xe3
      13'h1767: dout  = 8'b11111110; // 5991 : 254 - 0xfe
      13'h1768: dout  = 8'b01000110; // 5992 :  70 - 0x46
      13'h1769: dout  = 8'b11101010; // 5993 : 234 - 0xea
      13'h176A: dout  = 8'b01110000; // 5994 : 112 - 0x70
      13'h176B: dout  = 8'b00111010; // 5995 :  58 - 0x3a
      13'h176C: dout  = 8'b01101100; // 5996 : 108 - 0x6c
      13'h176D: dout  = 8'b10111000; // 5997 : 184 - 0xb8
      13'h176E: dout  = 8'b00011100; // 5998 :  28 - 0x1c
      13'h176F: dout  = 8'b00000000; // 5999 :   0 - 0x0
      13'h1770: dout  = 8'b11111111; // 6000 : 255 - 0xff -- Background 0x77
      13'h1771: dout  = 8'b11111111; // 6001 : 255 - 0xff
      13'h1772: dout  = 8'b11111111; // 6002 : 255 - 0xff
      13'h1773: dout  = 8'b11111111; // 6003 : 255 - 0xff
      13'h1774: dout  = 8'b11111111; // 6004 : 255 - 0xff
      13'h1775: dout  = 8'b11111111; // 6005 : 255 - 0xff
      13'h1776: dout  = 8'b11111111; // 6006 : 255 - 0xff
      13'h1777: dout  = 8'b11111111; // 6007 : 255 - 0xff
      13'h1778: dout  = 8'b10000001; // 6008 : 129 - 0x81
      13'h1779: dout  = 8'b11111111; // 6009 : 255 - 0xff
      13'h177A: dout  = 8'b11111101; // 6010 : 253 - 0xfd
      13'h177B: dout  = 8'b11111111; // 6011 : 255 - 0xff
      13'h177C: dout  = 8'b10111111; // 6012 : 191 - 0xbf
      13'h177D: dout  = 8'b11111111; // 6013 : 255 - 0xff
      13'h177E: dout  = 8'b11111111; // 6014 : 255 - 0xff
      13'h177F: dout  = 8'b11110111; // 6015 : 247 - 0xf7
      13'h1780: dout  = 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout  = 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout  = 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout  = 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout  = 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout  = 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout  = 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout  = 8'b00000000; // 6023 :   0 - 0x0
      13'h1788: dout  = 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout  = 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout  = 8'b00000000; // 6026 :   0 - 0x0
      13'h178B: dout  = 8'b00000000; // 6027 :   0 - 0x0
      13'h178C: dout  = 8'b00000000; // 6028 :   0 - 0x0
      13'h178D: dout  = 8'b00000000; // 6029 :   0 - 0x0
      13'h178E: dout  = 8'b00000000; // 6030 :   0 - 0x0
      13'h178F: dout  = 8'b00000000; // 6031 :   0 - 0x0
      13'h1790: dout  = 8'b00000000; // 6032 :   0 - 0x0 -- Background 0x79
      13'h1791: dout  = 8'b00000000; // 6033 :   0 - 0x0
      13'h1792: dout  = 8'b00000000; // 6034 :   0 - 0x0
      13'h1793: dout  = 8'b00000000; // 6035 :   0 - 0x0
      13'h1794: dout  = 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout  = 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout  = 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout  = 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout  = 8'b00000000; // 6040 :   0 - 0x0
      13'h1799: dout  = 8'b00000000; // 6041 :   0 - 0x0
      13'h179A: dout  = 8'b00000000; // 6042 :   0 - 0x0
      13'h179B: dout  = 8'b00000000; // 6043 :   0 - 0x0
      13'h179C: dout  = 8'b00000000; // 6044 :   0 - 0x0
      13'h179D: dout  = 8'b00000000; // 6045 :   0 - 0x0
      13'h179E: dout  = 8'b00000000; // 6046 :   0 - 0x0
      13'h179F: dout  = 8'b00000000; // 6047 :   0 - 0x0
      13'h17A0: dout  = 8'b00000000; // 6048 :   0 - 0x0 -- Background 0x7a
      13'h17A1: dout  = 8'b00000000; // 6049 :   0 - 0x0
      13'h17A2: dout  = 8'b00000000; // 6050 :   0 - 0x0
      13'h17A3: dout  = 8'b00000000; // 6051 :   0 - 0x0
      13'h17A4: dout  = 8'b00000000; // 6052 :   0 - 0x0
      13'h17A5: dout  = 8'b00000000; // 6053 :   0 - 0x0
      13'h17A6: dout  = 8'b00000000; // 6054 :   0 - 0x0
      13'h17A7: dout  = 8'b00000000; // 6055 :   0 - 0x0
      13'h17A8: dout  = 8'b00000000; // 6056 :   0 - 0x0
      13'h17A9: dout  = 8'b00000000; // 6057 :   0 - 0x0
      13'h17AA: dout  = 8'b00000000; // 6058 :   0 - 0x0
      13'h17AB: dout  = 8'b00000000; // 6059 :   0 - 0x0
      13'h17AC: dout  = 8'b00000000; // 6060 :   0 - 0x0
      13'h17AD: dout  = 8'b00000000; // 6061 :   0 - 0x0
      13'h17AE: dout  = 8'b00000000; // 6062 :   0 - 0x0
      13'h17AF: dout  = 8'b00000000; // 6063 :   0 - 0x0
      13'h17B0: dout  = 8'b00000000; // 6064 :   0 - 0x0 -- Background 0x7b
      13'h17B1: dout  = 8'b00000000; // 6065 :   0 - 0x0
      13'h17B2: dout  = 8'b00000000; // 6066 :   0 - 0x0
      13'h17B3: dout  = 8'b00000000; // 6067 :   0 - 0x0
      13'h17B4: dout  = 8'b00000000; // 6068 :   0 - 0x0
      13'h17B5: dout  = 8'b00000000; // 6069 :   0 - 0x0
      13'h17B6: dout  = 8'b00000000; // 6070 :   0 - 0x0
      13'h17B7: dout  = 8'b00000000; // 6071 :   0 - 0x0
      13'h17B8: dout  = 8'b00000000; // 6072 :   0 - 0x0
      13'h17B9: dout  = 8'b00000000; // 6073 :   0 - 0x0
      13'h17BA: dout  = 8'b00000000; // 6074 :   0 - 0x0
      13'h17BB: dout  = 8'b00000000; // 6075 :   0 - 0x0
      13'h17BC: dout  = 8'b00000000; // 6076 :   0 - 0x0
      13'h17BD: dout  = 8'b00000000; // 6077 :   0 - 0x0
      13'h17BE: dout  = 8'b00000000; // 6078 :   0 - 0x0
      13'h17BF: dout  = 8'b00000000; // 6079 :   0 - 0x0
      13'h17C0: dout  = 8'b00100010; // 6080 :  34 - 0x22 -- Background 0x7c
      13'h17C1: dout  = 8'b01010101; // 6081 :  85 - 0x55
      13'h17C2: dout  = 8'b10101010; // 6082 : 170 - 0xaa
      13'h17C3: dout  = 8'b00000101; // 6083 :   5 - 0x5
      13'h17C4: dout  = 8'b00000100; // 6084 :   4 - 0x4
      13'h17C5: dout  = 8'b00001010; // 6085 :  10 - 0xa
      13'h17C6: dout  = 8'b01010000; // 6086 :  80 - 0x50
      13'h17C7: dout  = 8'b00000010; // 6087 :   2 - 0x2
      13'h17C8: dout  = 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout  = 8'b00100010; // 6089 :  34 - 0x22
      13'h17CA: dout  = 8'b01110111; // 6090 : 119 - 0x77
      13'h17CB: dout  = 8'b11111111; // 6091 : 255 - 0xff
      13'h17CC: dout  = 8'b11111011; // 6092 : 251 - 0xfb
      13'h17CD: dout  = 8'b11110101; // 6093 : 245 - 0xf5
      13'h17CE: dout  = 8'b11101111; // 6094 : 239 - 0xef
      13'h17CF: dout  = 8'b11111111; // 6095 : 255 - 0xff
      13'h17D0: dout  = 8'b01110011; // 6096 : 115 - 0x73 -- Background 0x7d
      13'h17D1: dout  = 8'b11111111; // 6097 : 255 - 0xff
      13'h17D2: dout  = 8'b11111111; // 6098 : 255 - 0xff
      13'h17D3: dout  = 8'b10111101; // 6099 : 189 - 0xbd
      13'h17D4: dout  = 8'b01101110; // 6100 : 110 - 0x6e
      13'h17D5: dout  = 8'b00001010; // 6101 :  10 - 0xa
      13'h17D6: dout  = 8'b01010000; // 6102 :  80 - 0x50
      13'h17D7: dout  = 8'b00000010; // 6103 :   2 - 0x2
      13'h17D8: dout  = 8'b00000000; // 6104 :   0 - 0x0
      13'h17D9: dout  = 8'b01110011; // 6105 : 115 - 0x73
      13'h17DA: dout  = 8'b11111111; // 6106 : 255 - 0xff
      13'h17DB: dout  = 8'b11111111; // 6107 : 255 - 0xff
      13'h17DC: dout  = 8'b11111011; // 6108 : 251 - 0xfb
      13'h17DD: dout  = 8'b11111101; // 6109 : 253 - 0xfd
      13'h17DE: dout  = 8'b11101111; // 6110 : 239 - 0xef
      13'h17DF: dout  = 8'b11111111; // 6111 : 255 - 0xff
      13'h17E0: dout  = 8'b00100000; // 6112 :  32 - 0x20 -- Background 0x7e
      13'h17E1: dout  = 8'b01010000; // 6113 :  80 - 0x50
      13'h17E2: dout  = 8'b10000100; // 6114 : 132 - 0x84
      13'h17E3: dout  = 8'b00000000; // 6115 :   0 - 0x0
      13'h17E4: dout  = 8'b00100100; // 6116 :  36 - 0x24
      13'h17E5: dout  = 8'b01011010; // 6117 :  90 - 0x5a
      13'h17E6: dout  = 8'b00010000; // 6118 :  16 - 0x10
      13'h17E7: dout  = 8'b00000000; // 6119 :   0 - 0x0
      13'h17E8: dout  = 8'b11011111; // 6120 : 223 - 0xdf
      13'h17E9: dout  = 8'b10101111; // 6121 : 175 - 0xaf
      13'h17EA: dout  = 8'b01111111; // 6122 : 127 - 0x7f
      13'h17EB: dout  = 8'b11111111; // 6123 : 255 - 0xff
      13'h17EC: dout  = 8'b11111011; // 6124 : 251 - 0xfb
      13'h17ED: dout  = 8'b11110101; // 6125 : 245 - 0xf5
      13'h17EE: dout  = 8'b11101111; // 6126 : 239 - 0xef
      13'h17EF: dout  = 8'b11111111; // 6127 : 255 - 0xff
      13'h17F0: dout  = 8'b11111111; // 6128 : 255 - 0xff -- Background 0x7f
      13'h17F1: dout  = 8'b01010000; // 6129 :  80 - 0x50
      13'h17F2: dout  = 8'b10000100; // 6130 : 132 - 0x84
      13'h17F3: dout  = 8'b00000000; // 6131 :   0 - 0x0
      13'h17F4: dout  = 8'b00100100; // 6132 :  36 - 0x24
      13'h17F5: dout  = 8'b01011010; // 6133 :  90 - 0x5a
      13'h17F6: dout  = 8'b00010000; // 6134 :  16 - 0x10
      13'h17F7: dout  = 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout  = 8'b00000000; // 6136 :   0 - 0x0
      13'h17F9: dout  = 8'b10101111; // 6137 : 175 - 0xaf
      13'h17FA: dout  = 8'b01111111; // 6138 : 127 - 0x7f
      13'h17FB: dout  = 8'b11111111; // 6139 : 255 - 0xff
      13'h17FC: dout  = 8'b11111011; // 6140 : 251 - 0xfb
      13'h17FD: dout  = 8'b11110101; // 6141 : 245 - 0xf5
      13'h17FE: dout  = 8'b11101111; // 6142 : 239 - 0xef
      13'h17FF: dout  = 8'b11111111; // 6143 : 255 - 0xff
      13'h1800: dout  = 8'b11111111; // 6144 : 255 - 0xff -- Background 0x80
      13'h1801: dout  = 8'b10000000; // 6145 : 128 - 0x80
      13'h1802: dout  = 8'b11001111; // 6146 : 207 - 0xcf
      13'h1803: dout  = 8'b01001000; // 6147 :  72 - 0x48
      13'h1804: dout  = 8'b11001111; // 6148 : 207 - 0xcf
      13'h1805: dout  = 8'b10000000; // 6149 : 128 - 0x80
      13'h1806: dout  = 8'b11001111; // 6150 : 207 - 0xcf
      13'h1807: dout  = 8'b01001000; // 6151 :  72 - 0x48
      13'h1808: dout  = 8'b00000000; // 6152 :   0 - 0x0
      13'h1809: dout  = 8'b01111111; // 6153 : 127 - 0x7f
      13'h180A: dout  = 8'b00110000; // 6154 :  48 - 0x30
      13'h180B: dout  = 8'b00110000; // 6155 :  48 - 0x30
      13'h180C: dout  = 8'b00110000; // 6156 :  48 - 0x30
      13'h180D: dout  = 8'b01111111; // 6157 : 127 - 0x7f
      13'h180E: dout  = 8'b00110000; // 6158 :  48 - 0x30
      13'h180F: dout  = 8'b00110000; // 6159 :  48 - 0x30
      13'h1810: dout  = 8'b11111111; // 6160 : 255 - 0xff -- Background 0x81
      13'h1811: dout  = 8'b10000000; // 6161 : 128 - 0x80
      13'h1812: dout  = 8'b11111111; // 6162 : 255 - 0xff
      13'h1813: dout  = 8'b10000000; // 6163 : 128 - 0x80
      13'h1814: dout  = 8'b10000000; // 6164 : 128 - 0x80
      13'h1815: dout  = 8'b11011111; // 6165 : 223 - 0xdf
      13'h1816: dout  = 8'b10110000; // 6166 : 176 - 0xb0
      13'h1817: dout  = 8'b11000000; // 6167 : 192 - 0xc0
      13'h1818: dout  = 8'b00000000; // 6168 :   0 - 0x0
      13'h1819: dout  = 8'b01111111; // 6169 : 127 - 0x7f
      13'h181A: dout  = 8'b00000000; // 6170 :   0 - 0x0
      13'h181B: dout  = 8'b01111111; // 6171 : 127 - 0x7f
      13'h181C: dout  = 8'b01111111; // 6172 : 127 - 0x7f
      13'h181D: dout  = 8'b00100000; // 6173 :  32 - 0x20
      13'h181E: dout  = 8'b01000000; // 6174 :  64 - 0x40
      13'h181F: dout  = 8'b00000000; // 6175 :   0 - 0x0
      13'h1820: dout  = 8'b11111111; // 6176 : 255 - 0xff -- Background 0x82
      13'h1821: dout  = 8'b00000001; // 6177 :   1 - 0x1
      13'h1822: dout  = 8'b11110011; // 6178 : 243 - 0xf3
      13'h1823: dout  = 8'b00010010; // 6179 :  18 - 0x12
      13'h1824: dout  = 8'b11110011; // 6180 : 243 - 0xf3
      13'h1825: dout  = 8'b00000001; // 6181 :   1 - 0x1
      13'h1826: dout  = 8'b11110011; // 6182 : 243 - 0xf3
      13'h1827: dout  = 8'b00010010; // 6183 :  18 - 0x12
      13'h1828: dout  = 8'b00000000; // 6184 :   0 - 0x0
      13'h1829: dout  = 8'b11111110; // 6185 : 254 - 0xfe
      13'h182A: dout  = 8'b00001100; // 6186 :  12 - 0xc
      13'h182B: dout  = 8'b00001100; // 6187 :  12 - 0xc
      13'h182C: dout  = 8'b00001100; // 6188 :  12 - 0xc
      13'h182D: dout  = 8'b11111110; // 6189 : 254 - 0xfe
      13'h182E: dout  = 8'b00001100; // 6190 :  12 - 0xc
      13'h182F: dout  = 8'b00001100; // 6191 :  12 - 0xc
      13'h1830: dout  = 8'b11111111; // 6192 : 255 - 0xff -- Background 0x83
      13'h1831: dout  = 8'b00000000; // 6193 :   0 - 0x0
      13'h1832: dout  = 8'b11111111; // 6194 : 255 - 0xff
      13'h1833: dout  = 8'b00000000; // 6195 :   0 - 0x0
      13'h1834: dout  = 8'b00000000; // 6196 :   0 - 0x0
      13'h1835: dout  = 8'b11111111; // 6197 : 255 - 0xff
      13'h1836: dout  = 8'b00000000; // 6198 :   0 - 0x0
      13'h1837: dout  = 8'b00000000; // 6199 :   0 - 0x0
      13'h1838: dout  = 8'b00000000; // 6200 :   0 - 0x0
      13'h1839: dout  = 8'b11111111; // 6201 : 255 - 0xff
      13'h183A: dout  = 8'b00000000; // 6202 :   0 - 0x0
      13'h183B: dout  = 8'b11111111; // 6203 : 255 - 0xff
      13'h183C: dout  = 8'b11111111; // 6204 : 255 - 0xff
      13'h183D: dout  = 8'b00000000; // 6205 :   0 - 0x0
      13'h183E: dout  = 8'b00000000; // 6206 :   0 - 0x0
      13'h183F: dout  = 8'b00000000; // 6207 :   0 - 0x0
      13'h1840: dout  = 8'b11111111; // 6208 : 255 - 0xff -- Background 0x84
      13'h1841: dout  = 8'b10000010; // 6209 : 130 - 0x82
      13'h1842: dout  = 8'b00010000; // 6210 :  16 - 0x10
      13'h1843: dout  = 8'b00000000; // 6211 :   0 - 0x0
      13'h1844: dout  = 8'b00000000; // 6212 :   0 - 0x0
      13'h1845: dout  = 8'b00010000; // 6213 :  16 - 0x10
      13'h1846: dout  = 8'b01000100; // 6214 :  68 - 0x44
      13'h1847: dout  = 8'b11111111; // 6215 : 255 - 0xff
      13'h1848: dout  = 8'b00000000; // 6216 :   0 - 0x0
      13'h1849: dout  = 8'b11111111; // 6217 : 255 - 0xff
      13'h184A: dout  = 8'b11111111; // 6218 : 255 - 0xff
      13'h184B: dout  = 8'b11111111; // 6219 : 255 - 0xff
      13'h184C: dout  = 8'b11111111; // 6220 : 255 - 0xff
      13'h184D: dout  = 8'b11101111; // 6221 : 239 - 0xef
      13'h184E: dout  = 8'b10111011; // 6222 : 187 - 0xbb
      13'h184F: dout  = 8'b00000000; // 6223 :   0 - 0x0
      13'h1850: dout  = 8'b11111111; // 6224 : 255 - 0xff -- Background 0x85
      13'h1851: dout  = 8'b00000001; // 6225 :   1 - 0x1
      13'h1852: dout  = 8'b11111111; // 6226 : 255 - 0xff
      13'h1853: dout  = 8'b00000001; // 6227 :   1 - 0x1
      13'h1854: dout  = 8'b00000001; // 6228 :   1 - 0x1
      13'h1855: dout  = 8'b11110011; // 6229 : 243 - 0xf3
      13'h1856: dout  = 8'b00001101; // 6230 :  13 - 0xd
      13'h1857: dout  = 8'b00000011; // 6231 :   3 - 0x3
      13'h1858: dout  = 8'b00000000; // 6232 :   0 - 0x0
      13'h1859: dout  = 8'b11111110; // 6233 : 254 - 0xfe
      13'h185A: dout  = 8'b00000000; // 6234 :   0 - 0x0
      13'h185B: dout  = 8'b11111110; // 6235 : 254 - 0xfe
      13'h185C: dout  = 8'b11111110; // 6236 : 254 - 0xfe
      13'h185D: dout  = 8'b00001100; // 6237 :  12 - 0xc
      13'h185E: dout  = 8'b00000010; // 6238 :   2 - 0x2
      13'h185F: dout  = 8'b00000000; // 6239 :   0 - 0x0
      13'h1860: dout  = 8'b00000000; // 6240 :   0 - 0x0 -- Background 0x86
      13'h1861: dout  = 8'b00000000; // 6241 :   0 - 0x0
      13'h1862: dout  = 8'b00000000; // 6242 :   0 - 0x0
      13'h1863: dout  = 8'b00000000; // 6243 :   0 - 0x0
      13'h1864: dout  = 8'b00000000; // 6244 :   0 - 0x0
      13'h1865: dout  = 8'b00000000; // 6245 :   0 - 0x0
      13'h1866: dout  = 8'b00000000; // 6246 :   0 - 0x0
      13'h1867: dout  = 8'b00000000; // 6247 :   0 - 0x0
      13'h1868: dout  = 8'b00000000; // 6248 :   0 - 0x0
      13'h1869: dout  = 8'b00000000; // 6249 :   0 - 0x0
      13'h186A: dout  = 8'b00000000; // 6250 :   0 - 0x0
      13'h186B: dout  = 8'b00000000; // 6251 :   0 - 0x0
      13'h186C: dout  = 8'b00000000; // 6252 :   0 - 0x0
      13'h186D: dout  = 8'b00000000; // 6253 :   0 - 0x0
      13'h186E: dout  = 8'b00000000; // 6254 :   0 - 0x0
      13'h186F: dout  = 8'b00000000; // 6255 :   0 - 0x0
      13'h1870: dout  = 8'b00000000; // 6256 :   0 - 0x0 -- Background 0x87
      13'h1871: dout  = 8'b00000000; // 6257 :   0 - 0x0
      13'h1872: dout  = 8'b00000000; // 6258 :   0 - 0x0
      13'h1873: dout  = 8'b00000000; // 6259 :   0 - 0x0
      13'h1874: dout  = 8'b00000000; // 6260 :   0 - 0x0
      13'h1875: dout  = 8'b00000000; // 6261 :   0 - 0x0
      13'h1876: dout  = 8'b00000000; // 6262 :   0 - 0x0
      13'h1877: dout  = 8'b00000000; // 6263 :   0 - 0x0
      13'h1878: dout  = 8'b00000000; // 6264 :   0 - 0x0
      13'h1879: dout  = 8'b00000000; // 6265 :   0 - 0x0
      13'h187A: dout  = 8'b00000000; // 6266 :   0 - 0x0
      13'h187B: dout  = 8'b00000000; // 6267 :   0 - 0x0
      13'h187C: dout  = 8'b00000000; // 6268 :   0 - 0x0
      13'h187D: dout  = 8'b00000000; // 6269 :   0 - 0x0
      13'h187E: dout  = 8'b00000000; // 6270 :   0 - 0x0
      13'h187F: dout  = 8'b00000000; // 6271 :   0 - 0x0
      13'h1880: dout  = 8'b00000111; // 6272 :   7 - 0x7 -- Background 0x88
      13'h1881: dout  = 8'b00011110; // 6273 :  30 - 0x1e
      13'h1882: dout  = 8'b00101111; // 6274 :  47 - 0x2f
      13'h1883: dout  = 8'b01010011; // 6275 :  83 - 0x53
      13'h1884: dout  = 8'b01101110; // 6276 : 110 - 0x6e
      13'h1885: dout  = 8'b11011011; // 6277 : 219 - 0xdb
      13'h1886: dout  = 8'b11111010; // 6278 : 250 - 0xfa
      13'h1887: dout  = 8'b11010101; // 6279 : 213 - 0xd5
      13'h1888: dout  = 8'b00000000; // 6280 :   0 - 0x0
      13'h1889: dout  = 8'b00000111; // 6281 :   7 - 0x7
      13'h188A: dout  = 8'b00011111; // 6282 :  31 - 0x1f
      13'h188B: dout  = 8'b00111100; // 6283 :  60 - 0x3c
      13'h188C: dout  = 8'b00110001; // 6284 :  49 - 0x31
      13'h188D: dout  = 8'b01110100; // 6285 : 116 - 0x74
      13'h188E: dout  = 8'b01100101; // 6286 : 101 - 0x65
      13'h188F: dout  = 8'b01101010; // 6287 : 106 - 0x6a
      13'h1890: dout  = 8'b10111011; // 6288 : 187 - 0xbb -- Background 0x89
      13'h1891: dout  = 8'b11110010; // 6289 : 242 - 0xf2
      13'h1892: dout  = 8'b11011101; // 6290 : 221 - 0xdd
      13'h1893: dout  = 8'b01001111; // 6291 :  79 - 0x4f
      13'h1894: dout  = 8'b01111011; // 6292 : 123 - 0x7b
      13'h1895: dout  = 8'b00110010; // 6293 :  50 - 0x32
      13'h1896: dout  = 8'b00011111; // 6294 :  31 - 0x1f
      13'h1897: dout  = 8'b00000111; // 6295 :   7 - 0x7
      13'h1898: dout  = 8'b01100100; // 6296 : 100 - 0x64
      13'h1899: dout  = 8'b01101101; // 6297 : 109 - 0x6d
      13'h189A: dout  = 8'b01110010; // 6298 : 114 - 0x72
      13'h189B: dout  = 8'b00110000; // 6299 :  48 - 0x30
      13'h189C: dout  = 8'b00111100; // 6300 :  60 - 0x3c
      13'h189D: dout  = 8'b00011111; // 6301 :  31 - 0x1f
      13'h189E: dout  = 8'b00000111; // 6302 :   7 - 0x7
      13'h189F: dout  = 8'b00000000; // 6303 :   0 - 0x0
      13'h18A0: dout  = 8'b11100000; // 6304 : 224 - 0xe0 -- Background 0x8a
      13'h18A1: dout  = 8'b11011000; // 6305 : 216 - 0xd8
      13'h18A2: dout  = 8'b01010100; // 6306 :  84 - 0x54
      13'h18A3: dout  = 8'b11101010; // 6307 : 234 - 0xea
      13'h18A4: dout  = 8'b10111010; // 6308 : 186 - 0xba
      13'h18A5: dout  = 8'b10010011; // 6309 : 147 - 0x93
      13'h18A6: dout  = 8'b11011111; // 6310 : 223 - 0xdf
      13'h18A7: dout  = 8'b10111101; // 6311 : 189 - 0xbd
      13'h18A8: dout  = 8'b00000000; // 6312 :   0 - 0x0
      13'h18A9: dout  = 8'b11100000; // 6313 : 224 - 0xe0
      13'h18AA: dout  = 8'b11111000; // 6314 : 248 - 0xf8
      13'h18AB: dout  = 8'b00111100; // 6315 :  60 - 0x3c
      13'h18AC: dout  = 8'b01001100; // 6316 :  76 - 0x4c
      13'h18AD: dout  = 8'b01101110; // 6317 : 110 - 0x6e
      13'h18AE: dout  = 8'b00100110; // 6318 :  38 - 0x26
      13'h18AF: dout  = 8'b01000110; // 6319 :  70 - 0x46
      13'h18B0: dout  = 8'b01101011; // 6320 : 107 - 0x6b -- Background 0x8b
      13'h18B1: dout  = 8'b10011111; // 6321 : 159 - 0x9f
      13'h18B2: dout  = 8'b01011101; // 6322 :  93 - 0x5d
      13'h18B3: dout  = 8'b10110110; // 6323 : 182 - 0xb6
      13'h18B4: dout  = 8'b11101010; // 6324 : 234 - 0xea
      13'h18B5: dout  = 8'b11001100; // 6325 : 204 - 0xcc
      13'h18B6: dout  = 8'b01111000; // 6326 : 120 - 0x78
      13'h18B7: dout  = 8'b11100000; // 6327 : 224 - 0xe0
      13'h18B8: dout  = 8'b10010110; // 6328 : 150 - 0x96
      13'h18B9: dout  = 8'b01100110; // 6329 : 102 - 0x66
      13'h18BA: dout  = 8'b10101110; // 6330 : 174 - 0xae
      13'h18BB: dout  = 8'b01001100; // 6331 :  76 - 0x4c
      13'h18BC: dout  = 8'b00111100; // 6332 :  60 - 0x3c
      13'h18BD: dout  = 8'b11111000; // 6333 : 248 - 0xf8
      13'h18BE: dout  = 8'b11100000; // 6334 : 224 - 0xe0
      13'h18BF: dout  = 8'b00000000; // 6335 :   0 - 0x0
      13'h18C0: dout  = 8'b00000111; // 6336 :   7 - 0x7 -- Background 0x8c
      13'h18C1: dout  = 8'b00011000; // 6337 :  24 - 0x18
      13'h18C2: dout  = 8'b00100011; // 6338 :  35 - 0x23
      13'h18C3: dout  = 8'b01001100; // 6339 :  76 - 0x4c
      13'h18C4: dout  = 8'b01110000; // 6340 : 112 - 0x70
      13'h18C5: dout  = 8'b10100001; // 6341 : 161 - 0xa1
      13'h18C6: dout  = 8'b10100110; // 6342 : 166 - 0xa6
      13'h18C7: dout  = 8'b10101000; // 6343 : 168 - 0xa8
      13'h18C8: dout  = 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout  = 8'b00000111; // 6345 :   7 - 0x7
      13'h18CA: dout  = 8'b00011111; // 6346 :  31 - 0x1f
      13'h18CB: dout  = 8'b00111111; // 6347 :  63 - 0x3f
      13'h18CC: dout  = 8'b00111111; // 6348 :  63 - 0x3f
      13'h18CD: dout  = 8'b01111111; // 6349 : 127 - 0x7f
      13'h18CE: dout  = 8'b01111111; // 6350 : 127 - 0x7f
      13'h18CF: dout  = 8'b01111111; // 6351 : 127 - 0x7f
      13'h18D0: dout  = 8'b10100101; // 6352 : 165 - 0xa5 -- Background 0x8d
      13'h18D1: dout  = 8'b10100010; // 6353 : 162 - 0xa2
      13'h18D2: dout  = 8'b10010000; // 6354 : 144 - 0x90
      13'h18D3: dout  = 8'b01001000; // 6355 :  72 - 0x48
      13'h18D4: dout  = 8'b01000111; // 6356 :  71 - 0x47
      13'h18D5: dout  = 8'b00100000; // 6357 :  32 - 0x20
      13'h18D6: dout  = 8'b00011001; // 6358 :  25 - 0x19
      13'h18D7: dout  = 8'b00000111; // 6359 :   7 - 0x7
      13'h18D8: dout  = 8'b01111111; // 6360 : 127 - 0x7f
      13'h18D9: dout  = 8'b01111111; // 6361 : 127 - 0x7f
      13'h18DA: dout  = 8'b01111111; // 6362 : 127 - 0x7f
      13'h18DB: dout  = 8'b00111111; // 6363 :  63 - 0x3f
      13'h18DC: dout  = 8'b00111111; // 6364 :  63 - 0x3f
      13'h18DD: dout  = 8'b00011111; // 6365 :  31 - 0x1f
      13'h18DE: dout  = 8'b00000111; // 6366 :   7 - 0x7
      13'h18DF: dout  = 8'b00000000; // 6367 :   0 - 0x0
      13'h18E0: dout  = 8'b11100000; // 6368 : 224 - 0xe0 -- Background 0x8e
      13'h18E1: dout  = 8'b00011000; // 6369 :  24 - 0x18
      13'h18E2: dout  = 8'b00000100; // 6370 :   4 - 0x4
      13'h18E3: dout  = 8'b11000010; // 6371 : 194 - 0xc2
      13'h18E4: dout  = 8'b00110010; // 6372 :  50 - 0x32
      13'h18E5: dout  = 8'b00001001; // 6373 :   9 - 0x9
      13'h18E6: dout  = 8'b11000101; // 6374 : 197 - 0xc5
      13'h18E7: dout  = 8'b00100101; // 6375 :  37 - 0x25
      13'h18E8: dout  = 8'b00000000; // 6376 :   0 - 0x0
      13'h18E9: dout  = 8'b11100000; // 6377 : 224 - 0xe0
      13'h18EA: dout  = 8'b11111000; // 6378 : 248 - 0xf8
      13'h18EB: dout  = 8'b11111100; // 6379 : 252 - 0xfc
      13'h18EC: dout  = 8'b11111100; // 6380 : 252 - 0xfc
      13'h18ED: dout  = 8'b11111110; // 6381 : 254 - 0xfe
      13'h18EE: dout  = 8'b11111110; // 6382 : 254 - 0xfe
      13'h18EF: dout  = 8'b11111110; // 6383 : 254 - 0xfe
      13'h18F0: dout  = 8'b10100101; // 6384 : 165 - 0xa5 -- Background 0x8f
      13'h18F1: dout  = 8'b01100101; // 6385 : 101 - 0x65
      13'h18F2: dout  = 8'b01000101; // 6386 :  69 - 0x45
      13'h18F3: dout  = 8'b10001010; // 6387 : 138 - 0x8a
      13'h18F4: dout  = 8'b10010010; // 6388 : 146 - 0x92
      13'h18F5: dout  = 8'b00100100; // 6389 :  36 - 0x24
      13'h18F6: dout  = 8'b11011000; // 6390 : 216 - 0xd8
      13'h18F7: dout  = 8'b11100000; // 6391 : 224 - 0xe0
      13'h18F8: dout  = 8'b11111110; // 6392 : 254 - 0xfe
      13'h18F9: dout  = 8'b11111110; // 6393 : 254 - 0xfe
      13'h18FA: dout  = 8'b11111110; // 6394 : 254 - 0xfe
      13'h18FB: dout  = 8'b11111100; // 6395 : 252 - 0xfc
      13'h18FC: dout  = 8'b11111100; // 6396 : 252 - 0xfc
      13'h18FD: dout  = 8'b11111000; // 6397 : 248 - 0xf8
      13'h18FE: dout  = 8'b11100000; // 6398 : 224 - 0xe0
      13'h18FF: dout  = 8'b00000000; // 6399 :   0 - 0x0
      13'h1900: dout  = 8'b00000000; // 6400 :   0 - 0x0 -- Background 0x90
      13'h1901: dout  = 8'b00000000; // 6401 :   0 - 0x0
      13'h1902: dout  = 8'b00100000; // 6402 :  32 - 0x20
      13'h1903: dout  = 8'b00110000; // 6403 :  48 - 0x30
      13'h1904: dout  = 8'b00101100; // 6404 :  44 - 0x2c
      13'h1905: dout  = 8'b00100010; // 6405 :  34 - 0x22
      13'h1906: dout  = 8'b00010001; // 6406 :  17 - 0x11
      13'h1907: dout  = 8'b00001000; // 6407 :   8 - 0x8
      13'h1908: dout  = 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout  = 8'b00000000; // 6409 :   0 - 0x0
      13'h190A: dout  = 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout  = 8'b00000000; // 6411 :   0 - 0x0
      13'h190C: dout  = 8'b00010000; // 6412 :  16 - 0x10
      13'h190D: dout  = 8'b00011100; // 6413 :  28 - 0x1c
      13'h190E: dout  = 8'b00001110; // 6414 :  14 - 0xe
      13'h190F: dout  = 8'b00000111; // 6415 :   7 - 0x7
      13'h1910: dout  = 8'b00000100; // 6416 :   4 - 0x4 -- Background 0x91
      13'h1911: dout  = 8'b11110010; // 6417 : 242 - 0xf2
      13'h1912: dout  = 8'b11001111; // 6418 : 207 - 0xcf
      13'h1913: dout  = 8'b00110000; // 6419 :  48 - 0x30
      13'h1914: dout  = 8'b00001100; // 6420 :  12 - 0xc
      13'h1915: dout  = 8'b11111111; // 6421 : 255 - 0xff
      13'h1916: dout  = 8'b10000000; // 6422 : 128 - 0x80
      13'h1917: dout  = 8'b11111111; // 6423 : 255 - 0xff
      13'h1918: dout  = 8'b00000011; // 6424 :   3 - 0x3
      13'h1919: dout  = 8'b00000001; // 6425 :   1 - 0x1
      13'h191A: dout  = 8'b00110000; // 6426 :  48 - 0x30
      13'h191B: dout  = 8'b00001111; // 6427 :  15 - 0xf
      13'h191C: dout  = 8'b00000011; // 6428 :   3 - 0x3
      13'h191D: dout  = 8'b00000000; // 6429 :   0 - 0x0
      13'h191E: dout  = 8'b01111111; // 6430 : 127 - 0x7f
      13'h191F: dout  = 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout  = 8'b01000010; // 6432 :  66 - 0x42 -- Background 0x92
      13'h1921: dout  = 8'b10100101; // 6433 : 165 - 0xa5
      13'h1922: dout  = 8'b10100101; // 6434 : 165 - 0xa5
      13'h1923: dout  = 8'b10011001; // 6435 : 153 - 0x99
      13'h1924: dout  = 8'b10011001; // 6436 : 153 - 0x99
      13'h1925: dout  = 8'b10011001; // 6437 : 153 - 0x99
      13'h1926: dout  = 8'b00000001; // 6438 :   1 - 0x1
      13'h1927: dout  = 8'b00000000; // 6439 :   0 - 0x0
      13'h1928: dout  = 8'b00000000; // 6440 :   0 - 0x0
      13'h1929: dout  = 8'b01000010; // 6441 :  66 - 0x42
      13'h192A: dout  = 8'b01000010; // 6442 :  66 - 0x42
      13'h192B: dout  = 8'b01100110; // 6443 : 102 - 0x66
      13'h192C: dout  = 8'b01100110; // 6444 : 102 - 0x66
      13'h192D: dout  = 8'b01100110; // 6445 : 102 - 0x66
      13'h192E: dout  = 8'b11111110; // 6446 : 254 - 0xfe
      13'h192F: dout  = 8'b11111111; // 6447 : 255 - 0xff
      13'h1930: dout  = 8'b11111111; // 6448 : 255 - 0xff -- Background 0x93
      13'h1931: dout  = 8'b11111111; // 6449 : 255 - 0xff
      13'h1932: dout  = 8'b11111111; // 6450 : 255 - 0xff
      13'h1933: dout  = 8'b10000001; // 6451 : 129 - 0x81
      13'h1934: dout  = 8'b11111111; // 6452 : 255 - 0xff
      13'h1935: dout  = 8'b11111111; // 6453 : 255 - 0xff
      13'h1936: dout  = 8'b11111111; // 6454 : 255 - 0xff
      13'h1937: dout  = 8'b10000001; // 6455 : 129 - 0x81
      13'h1938: dout  = 8'b01111110; // 6456 : 126 - 0x7e
      13'h1939: dout  = 8'b01111110; // 6457 : 126 - 0x7e
      13'h193A: dout  = 8'b01111110; // 6458 : 126 - 0x7e
      13'h193B: dout  = 8'b01111110; // 6459 : 126 - 0x7e
      13'h193C: dout  = 8'b01111110; // 6460 : 126 - 0x7e
      13'h193D: dout  = 8'b01111110; // 6461 : 126 - 0x7e
      13'h193E: dout  = 8'b01111110; // 6462 : 126 - 0x7e
      13'h193F: dout  = 8'b01111110; // 6463 : 126 - 0x7e
      13'h1940: dout  = 8'b00000000; // 6464 :   0 - 0x0 -- Background 0x94
      13'h1941: dout  = 8'b00000000; // 6465 :   0 - 0x0
      13'h1942: dout  = 8'b00000100; // 6466 :   4 - 0x4
      13'h1943: dout  = 8'b00001100; // 6467 :  12 - 0xc
      13'h1944: dout  = 8'b00110100; // 6468 :  52 - 0x34
      13'h1945: dout  = 8'b01000100; // 6469 :  68 - 0x44
      13'h1946: dout  = 8'b10001000; // 6470 : 136 - 0x88
      13'h1947: dout  = 8'b00010000; // 6471 :  16 - 0x10
      13'h1948: dout  = 8'b00000000; // 6472 :   0 - 0x0
      13'h1949: dout  = 8'b00000000; // 6473 :   0 - 0x0
      13'h194A: dout  = 8'b00000000; // 6474 :   0 - 0x0
      13'h194B: dout  = 8'b00000000; // 6475 :   0 - 0x0
      13'h194C: dout  = 8'b00001000; // 6476 :   8 - 0x8
      13'h194D: dout  = 8'b00111000; // 6477 :  56 - 0x38
      13'h194E: dout  = 8'b01110000; // 6478 : 112 - 0x70
      13'h194F: dout  = 8'b11100000; // 6479 : 224 - 0xe0
      13'h1950: dout  = 8'b00100000; // 6480 :  32 - 0x20 -- Background 0x95
      13'h1951: dout  = 8'b01001111; // 6481 :  79 - 0x4f
      13'h1952: dout  = 8'b11110011; // 6482 : 243 - 0xf3
      13'h1953: dout  = 8'b00001100; // 6483 :  12 - 0xc
      13'h1954: dout  = 8'b00110000; // 6484 :  48 - 0x30
      13'h1955: dout  = 8'b11111111; // 6485 : 255 - 0xff
      13'h1956: dout  = 8'b00000001; // 6486 :   1 - 0x1
      13'h1957: dout  = 8'b11111111; // 6487 : 255 - 0xff
      13'h1958: dout  = 8'b11000000; // 6488 : 192 - 0xc0
      13'h1959: dout  = 8'b10000000; // 6489 : 128 - 0x80
      13'h195A: dout  = 8'b00001100; // 6490 :  12 - 0xc
      13'h195B: dout  = 8'b11110000; // 6491 : 240 - 0xf0
      13'h195C: dout  = 8'b11000000; // 6492 : 192 - 0xc0
      13'h195D: dout  = 8'b00000000; // 6493 :   0 - 0x0
      13'h195E: dout  = 8'b11111110; // 6494 : 254 - 0xfe
      13'h195F: dout  = 8'b00000000; // 6495 :   0 - 0x0
      13'h1960: dout  = 8'b01111111; // 6496 : 127 - 0x7f -- Background 0x96
      13'h1961: dout  = 8'b11111111; // 6497 : 255 - 0xff
      13'h1962: dout  = 8'b11111111; // 6498 : 255 - 0xff
      13'h1963: dout  = 8'b11111111; // 6499 : 255 - 0xff
      13'h1964: dout  = 8'b11111011; // 6500 : 251 - 0xfb
      13'h1965: dout  = 8'b11111111; // 6501 : 255 - 0xff
      13'h1966: dout  = 8'b11111111; // 6502 : 255 - 0xff
      13'h1967: dout  = 8'b11111111; // 6503 : 255 - 0xff
      13'h1968: dout  = 8'b00000000; // 6504 :   0 - 0x0
      13'h1969: dout  = 8'b00111111; // 6505 :  63 - 0x3f
      13'h196A: dout  = 8'b01111111; // 6506 : 127 - 0x7f
      13'h196B: dout  = 8'b01111111; // 6507 : 127 - 0x7f
      13'h196C: dout  = 8'b01111111; // 6508 : 127 - 0x7f
      13'h196D: dout  = 8'b01111111; // 6509 : 127 - 0x7f
      13'h196E: dout  = 8'b01111111; // 6510 : 127 - 0x7f
      13'h196F: dout  = 8'b01111111; // 6511 : 127 - 0x7f
      13'h1970: dout  = 8'b11111111; // 6512 : 255 - 0xff -- Background 0x97
      13'h1971: dout  = 8'b11111111; // 6513 : 255 - 0xff
      13'h1972: dout  = 8'b11111111; // 6514 : 255 - 0xff
      13'h1973: dout  = 8'b11111111; // 6515 : 255 - 0xff
      13'h1974: dout  = 8'b11111111; // 6516 : 255 - 0xff
      13'h1975: dout  = 8'b11111111; // 6517 : 255 - 0xff
      13'h1976: dout  = 8'b11111110; // 6518 : 254 - 0xfe
      13'h1977: dout  = 8'b11111111; // 6519 : 255 - 0xff
      13'h1978: dout  = 8'b01111111; // 6520 : 127 - 0x7f
      13'h1979: dout  = 8'b01111111; // 6521 : 127 - 0x7f
      13'h197A: dout  = 8'b00111111; // 6522 :  63 - 0x3f
      13'h197B: dout  = 8'b01111111; // 6523 : 127 - 0x7f
      13'h197C: dout  = 8'b01111111; // 6524 : 127 - 0x7f
      13'h197D: dout  = 8'b01111111; // 6525 : 127 - 0x7f
      13'h197E: dout  = 8'b01111111; // 6526 : 127 - 0x7f
      13'h197F: dout  = 8'b01111111; // 6527 : 127 - 0x7f
      13'h1980: dout  = 8'b11111111; // 6528 : 255 - 0xff -- Background 0x98
      13'h1981: dout  = 8'b10111111; // 6529 : 191 - 0xbf
      13'h1982: dout  = 8'b11111111; // 6530 : 255 - 0xff
      13'h1983: dout  = 8'b11111111; // 6531 : 255 - 0xff
      13'h1984: dout  = 8'b11111011; // 6532 : 251 - 0xfb
      13'h1985: dout  = 8'b11111111; // 6533 : 255 - 0xff
      13'h1986: dout  = 8'b11111111; // 6534 : 255 - 0xff
      13'h1987: dout  = 8'b11111111; // 6535 : 255 - 0xff
      13'h1988: dout  = 8'b00000000; // 6536 :   0 - 0x0
      13'h1989: dout  = 8'b11011111; // 6537 : 223 - 0xdf
      13'h198A: dout  = 8'b11111111; // 6538 : 255 - 0xff
      13'h198B: dout  = 8'b11111111; // 6539 : 255 - 0xff
      13'h198C: dout  = 8'b11111111; // 6540 : 255 - 0xff
      13'h198D: dout  = 8'b11111111; // 6541 : 255 - 0xff
      13'h198E: dout  = 8'b11111111; // 6542 : 255 - 0xff
      13'h198F: dout  = 8'b11111111; // 6543 : 255 - 0xff
      13'h1990: dout  = 8'b11111111; // 6544 : 255 - 0xff -- Background 0x99
      13'h1991: dout  = 8'b11111111; // 6545 : 255 - 0xff
      13'h1992: dout  = 8'b11111111; // 6546 : 255 - 0xff
      13'h1993: dout  = 8'b11111111; // 6547 : 255 - 0xff
      13'h1994: dout  = 8'b11111111; // 6548 : 255 - 0xff
      13'h1995: dout  = 8'b11111111; // 6549 : 255 - 0xff
      13'h1996: dout  = 8'b11111110; // 6550 : 254 - 0xfe
      13'h1997: dout  = 8'b11111111; // 6551 : 255 - 0xff
      13'h1998: dout  = 8'b11111111; // 6552 : 255 - 0xff
      13'h1999: dout  = 8'b11111111; // 6553 : 255 - 0xff
      13'h199A: dout  = 8'b10111111; // 6554 : 191 - 0xbf
      13'h199B: dout  = 8'b11111111; // 6555 : 255 - 0xff
      13'h199C: dout  = 8'b11111111; // 6556 : 255 - 0xff
      13'h199D: dout  = 8'b11111111; // 6557 : 255 - 0xff
      13'h199E: dout  = 8'b11111111; // 6558 : 255 - 0xff
      13'h199F: dout  = 8'b11111111; // 6559 : 255 - 0xff
      13'h19A0: dout  = 8'b11111110; // 6560 : 254 - 0xfe -- Background 0x9a
      13'h19A1: dout  = 8'b11111111; // 6561 : 255 - 0xff
      13'h19A2: dout  = 8'b11111111; // 6562 : 255 - 0xff
      13'h19A3: dout  = 8'b11111111; // 6563 : 255 - 0xff
      13'h19A4: dout  = 8'b11111011; // 6564 : 251 - 0xfb
      13'h19A5: dout  = 8'b11111111; // 6565 : 255 - 0xff
      13'h19A6: dout  = 8'b11111111; // 6566 : 255 - 0xff
      13'h19A7: dout  = 8'b11111111; // 6567 : 255 - 0xff
      13'h19A8: dout  = 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout  = 8'b10111100; // 6569 : 188 - 0xbc
      13'h19AA: dout  = 8'b11111110; // 6570 : 254 - 0xfe
      13'h19AB: dout  = 8'b11111110; // 6571 : 254 - 0xfe
      13'h19AC: dout  = 8'b11111110; // 6572 : 254 - 0xfe
      13'h19AD: dout  = 8'b11111110; // 6573 : 254 - 0xfe
      13'h19AE: dout  = 8'b11111110; // 6574 : 254 - 0xfe
      13'h19AF: dout  = 8'b11111110; // 6575 : 254 - 0xfe
      13'h19B0: dout  = 8'b11111111; // 6576 : 255 - 0xff -- Background 0x9b
      13'h19B1: dout  = 8'b11111111; // 6577 : 255 - 0xff
      13'h19B2: dout  = 8'b11111111; // 6578 : 255 - 0xff
      13'h19B3: dout  = 8'b11111111; // 6579 : 255 - 0xff
      13'h19B4: dout  = 8'b11111111; // 6580 : 255 - 0xff
      13'h19B5: dout  = 8'b11111111; // 6581 : 255 - 0xff
      13'h19B6: dout  = 8'b11111111; // 6582 : 255 - 0xff
      13'h19B7: dout  = 8'b11111111; // 6583 : 255 - 0xff
      13'h19B8: dout  = 8'b11111110; // 6584 : 254 - 0xfe
      13'h19B9: dout  = 8'b11111110; // 6585 : 254 - 0xfe
      13'h19BA: dout  = 8'b10111110; // 6586 : 190 - 0xbe
      13'h19BB: dout  = 8'b11111110; // 6587 : 254 - 0xfe
      13'h19BC: dout  = 8'b11111110; // 6588 : 254 - 0xfe
      13'h19BD: dout  = 8'b11111110; // 6589 : 254 - 0xfe
      13'h19BE: dout  = 8'b11111110; // 6590 : 254 - 0xfe
      13'h19BF: dout  = 8'b11111110; // 6591 : 254 - 0xfe
      13'h19C0: dout  = 8'b11111111; // 6592 : 255 - 0xff -- Background 0x9c
      13'h19C1: dout  = 8'b11111111; // 6593 : 255 - 0xff
      13'h19C2: dout  = 8'b10100000; // 6594 : 160 - 0xa0
      13'h19C3: dout  = 8'b10010000; // 6595 : 144 - 0x90
      13'h19C4: dout  = 8'b10001000; // 6596 : 136 - 0x88
      13'h19C5: dout  = 8'b10000100; // 6597 : 132 - 0x84
      13'h19C6: dout  = 8'b01101010; // 6598 : 106 - 0x6a
      13'h19C7: dout  = 8'b00111111; // 6599 :  63 - 0x3f
      13'h19C8: dout  = 8'b00000000; // 6600 :   0 - 0x0
      13'h19C9: dout  = 8'b00111111; // 6601 :  63 - 0x3f
      13'h19CA: dout  = 8'b01011111; // 6602 :  95 - 0x5f
      13'h19CB: dout  = 8'b01101111; // 6603 : 111 - 0x6f
      13'h19CC: dout  = 8'b01110111; // 6604 : 119 - 0x77
      13'h19CD: dout  = 8'b01111011; // 6605 : 123 - 0x7b
      13'h19CE: dout  = 8'b00010101; // 6606 :  21 - 0x15
      13'h19CF: dout  = 8'b00000000; // 6607 :   0 - 0x0
      13'h19D0: dout  = 8'b11111111; // 6608 : 255 - 0xff -- Background 0x9d
      13'h19D1: dout  = 8'b11111111; // 6609 : 255 - 0xff
      13'h19D2: dout  = 8'b00100001; // 6610 :  33 - 0x21
      13'h19D3: dout  = 8'b00010001; // 6611 :  17 - 0x11
      13'h19D4: dout  = 8'b00001001; // 6612 :   9 - 0x9
      13'h19D5: dout  = 8'b00000101; // 6613 :   5 - 0x5
      13'h19D6: dout  = 8'b10101010; // 6614 : 170 - 0xaa
      13'h19D7: dout  = 8'b11111100; // 6615 : 252 - 0xfc
      13'h19D8: dout  = 8'b00000000; // 6616 :   0 - 0x0
      13'h19D9: dout  = 8'b10111110; // 6617 : 190 - 0xbe
      13'h19DA: dout  = 8'b11011110; // 6618 : 222 - 0xde
      13'h19DB: dout  = 8'b11101110; // 6619 : 238 - 0xee
      13'h19DC: dout  = 8'b11110110; // 6620 : 246 - 0xf6
      13'h19DD: dout  = 8'b11111010; // 6621 : 250 - 0xfa
      13'h19DE: dout  = 8'b01010100; // 6622 :  84 - 0x54
      13'h19DF: dout  = 8'b00000000; // 6623 :   0 - 0x0
      13'h19E0: dout  = 8'b11111111; // 6624 : 255 - 0xff -- Background 0x9e
      13'h19E1: dout  = 8'b11111111; // 6625 : 255 - 0xff
      13'h19E2: dout  = 8'b00100000; // 6626 :  32 - 0x20
      13'h19E3: dout  = 8'b00010000; // 6627 :  16 - 0x10
      13'h19E4: dout  = 8'b00001000; // 6628 :   8 - 0x8
      13'h19E5: dout  = 8'b00000100; // 6629 :   4 - 0x4
      13'h19E6: dout  = 8'b10101010; // 6630 : 170 - 0xaa
      13'h19E7: dout  = 8'b11111111; // 6631 : 255 - 0xff
      13'h19E8: dout  = 8'b00000000; // 6632 :   0 - 0x0
      13'h19E9: dout  = 8'b10111111; // 6633 : 191 - 0xbf
      13'h19EA: dout  = 8'b11011111; // 6634 : 223 - 0xdf
      13'h19EB: dout  = 8'b11101111; // 6635 : 239 - 0xef
      13'h19EC: dout  = 8'b11110111; // 6636 : 247 - 0xf7
      13'h19ED: dout  = 8'b11111011; // 6637 : 251 - 0xfb
      13'h19EE: dout  = 8'b01010101; // 6638 :  85 - 0x55
      13'h19EF: dout  = 8'b00000000; // 6639 :   0 - 0x0
      13'h19F0: dout  = 8'b00000000; // 6640 :   0 - 0x0 -- Background 0x9f
      13'h19F1: dout  = 8'b00000000; // 6641 :   0 - 0x0
      13'h19F2: dout  = 8'b00000000; // 6642 :   0 - 0x0
      13'h19F3: dout  = 8'b00000000; // 6643 :   0 - 0x0
      13'h19F4: dout  = 8'b00000000; // 6644 :   0 - 0x0
      13'h19F5: dout  = 8'b00000000; // 6645 :   0 - 0x0
      13'h19F6: dout  = 8'b00000000; // 6646 :   0 - 0x0
      13'h19F7: dout  = 8'b00000000; // 6647 :   0 - 0x0
      13'h19F8: dout  = 8'b00000000; // 6648 :   0 - 0x0
      13'h19F9: dout  = 8'b00000000; // 6649 :   0 - 0x0
      13'h19FA: dout  = 8'b00000000; // 6650 :   0 - 0x0
      13'h19FB: dout  = 8'b00000000; // 6651 :   0 - 0x0
      13'h19FC: dout  = 8'b00000000; // 6652 :   0 - 0x0
      13'h19FD: dout  = 8'b00000000; // 6653 :   0 - 0x0
      13'h19FE: dout  = 8'b00000000; // 6654 :   0 - 0x0
      13'h19FF: dout  = 8'b00000000; // 6655 :   0 - 0x0
      13'h1A00: dout  = 8'b11111111; // 6656 : 255 - 0xff -- Background 0xa0
      13'h1A01: dout  = 8'b11010101; // 6657 : 213 - 0xd5
      13'h1A02: dout  = 8'b11111111; // 6658 : 255 - 0xff
      13'h1A03: dout  = 8'b00000010; // 6659 :   2 - 0x2
      13'h1A04: dout  = 8'b00000010; // 6660 :   2 - 0x2
      13'h1A05: dout  = 8'b00000010; // 6661 :   2 - 0x2
      13'h1A06: dout  = 8'b00000010; // 6662 :   2 - 0x2
      13'h1A07: dout  = 8'b00000010; // 6663 :   2 - 0x2
      13'h1A08: dout  = 8'b00000000; // 6664 :   0 - 0x0
      13'h1A09: dout  = 8'b01111111; // 6665 : 127 - 0x7f
      13'h1A0A: dout  = 8'b00000000; // 6666 :   0 - 0x0
      13'h1A0B: dout  = 8'b00000001; // 6667 :   1 - 0x1
      13'h1A0C: dout  = 8'b00000001; // 6668 :   1 - 0x1
      13'h1A0D: dout  = 8'b00000001; // 6669 :   1 - 0x1
      13'h1A0E: dout  = 8'b00000001; // 6670 :   1 - 0x1
      13'h1A0F: dout  = 8'b00000001; // 6671 :   1 - 0x1
      13'h1A10: dout  = 8'b00000010; // 6672 :   2 - 0x2 -- Background 0xa1
      13'h1A11: dout  = 8'b00000010; // 6673 :   2 - 0x2
      13'h1A12: dout  = 8'b00000010; // 6674 :   2 - 0x2
      13'h1A13: dout  = 8'b00000010; // 6675 :   2 - 0x2
      13'h1A14: dout  = 8'b00000010; // 6676 :   2 - 0x2
      13'h1A15: dout  = 8'b00000010; // 6677 :   2 - 0x2
      13'h1A16: dout  = 8'b00000010; // 6678 :   2 - 0x2
      13'h1A17: dout  = 8'b00000010; // 6679 :   2 - 0x2
      13'h1A18: dout  = 8'b00000001; // 6680 :   1 - 0x1
      13'h1A19: dout  = 8'b00000001; // 6681 :   1 - 0x1
      13'h1A1A: dout  = 8'b00000001; // 6682 :   1 - 0x1
      13'h1A1B: dout  = 8'b00000001; // 6683 :   1 - 0x1
      13'h1A1C: dout  = 8'b00000001; // 6684 :   1 - 0x1
      13'h1A1D: dout  = 8'b00000001; // 6685 :   1 - 0x1
      13'h1A1E: dout  = 8'b00000001; // 6686 :   1 - 0x1
      13'h1A1F: dout  = 8'b00000001; // 6687 :   1 - 0x1
      13'h1A20: dout  = 8'b11111111; // 6688 : 255 - 0xff -- Background 0xa2
      13'h1A21: dout  = 8'b01010101; // 6689 :  85 - 0x55
      13'h1A22: dout  = 8'b11111111; // 6690 : 255 - 0xff
      13'h1A23: dout  = 8'b01000000; // 6691 :  64 - 0x40
      13'h1A24: dout  = 8'b01000000; // 6692 :  64 - 0x40
      13'h1A25: dout  = 8'b01000000; // 6693 :  64 - 0x40
      13'h1A26: dout  = 8'b01000000; // 6694 :  64 - 0x40
      13'h1A27: dout  = 8'b01000000; // 6695 :  64 - 0x40
      13'h1A28: dout  = 8'b00000000; // 6696 :   0 - 0x0
      13'h1A29: dout  = 8'b11111110; // 6697 : 254 - 0xfe
      13'h1A2A: dout  = 8'b00000000; // 6698 :   0 - 0x0
      13'h1A2B: dout  = 8'b10000000; // 6699 : 128 - 0x80
      13'h1A2C: dout  = 8'b10000000; // 6700 : 128 - 0x80
      13'h1A2D: dout  = 8'b10000000; // 6701 : 128 - 0x80
      13'h1A2E: dout  = 8'b10000000; // 6702 : 128 - 0x80
      13'h1A2F: dout  = 8'b10000000; // 6703 : 128 - 0x80
      13'h1A30: dout  = 8'b01000000; // 6704 :  64 - 0x40 -- Background 0xa3
      13'h1A31: dout  = 8'b01000000; // 6705 :  64 - 0x40
      13'h1A32: dout  = 8'b01000000; // 6706 :  64 - 0x40
      13'h1A33: dout  = 8'b01000000; // 6707 :  64 - 0x40
      13'h1A34: dout  = 8'b01000000; // 6708 :  64 - 0x40
      13'h1A35: dout  = 8'b01000000; // 6709 :  64 - 0x40
      13'h1A36: dout  = 8'b01000000; // 6710 :  64 - 0x40
      13'h1A37: dout  = 8'b01000000; // 6711 :  64 - 0x40
      13'h1A38: dout  = 8'b10000000; // 6712 : 128 - 0x80
      13'h1A39: dout  = 8'b10000000; // 6713 : 128 - 0x80
      13'h1A3A: dout  = 8'b10000000; // 6714 : 128 - 0x80
      13'h1A3B: dout  = 8'b10000000; // 6715 : 128 - 0x80
      13'h1A3C: dout  = 8'b10000000; // 6716 : 128 - 0x80
      13'h1A3D: dout  = 8'b10000000; // 6717 : 128 - 0x80
      13'h1A3E: dout  = 8'b10000000; // 6718 : 128 - 0x80
      13'h1A3F: dout  = 8'b10000000; // 6719 : 128 - 0x80
      13'h1A40: dout  = 8'b00110001; // 6720 :  49 - 0x31 -- Background 0xa4
      13'h1A41: dout  = 8'b01001000; // 6721 :  72 - 0x48
      13'h1A42: dout  = 8'b01000101; // 6722 :  69 - 0x45
      13'h1A43: dout  = 8'b10000101; // 6723 : 133 - 0x85
      13'h1A44: dout  = 8'b10000011; // 6724 : 131 - 0x83
      13'h1A45: dout  = 8'b10000010; // 6725 : 130 - 0x82
      13'h1A46: dout  = 8'b01100010; // 6726 :  98 - 0x62
      13'h1A47: dout  = 8'b00010010; // 6727 :  18 - 0x12
      13'h1A48: dout  = 8'b00000000; // 6728 :   0 - 0x0
      13'h1A49: dout  = 8'b00110000; // 6729 :  48 - 0x30
      13'h1A4A: dout  = 8'b00111000; // 6730 :  56 - 0x38
      13'h1A4B: dout  = 8'b01111000; // 6731 : 120 - 0x78
      13'h1A4C: dout  = 8'b01111100; // 6732 : 124 - 0x7c
      13'h1A4D: dout  = 8'b01111101; // 6733 : 125 - 0x7d
      13'h1A4E: dout  = 8'b00011101; // 6734 :  29 - 0x1d
      13'h1A4F: dout  = 8'b00001101; // 6735 :  13 - 0xd
      13'h1A50: dout  = 8'b00110010; // 6736 :  50 - 0x32 -- Background 0xa5
      13'h1A51: dout  = 8'b00100010; // 6737 :  34 - 0x22
      13'h1A52: dout  = 8'b01000010; // 6738 :  66 - 0x42
      13'h1A53: dout  = 8'b01000000; // 6739 :  64 - 0x40
      13'h1A54: dout  = 8'b01000000; // 6740 :  64 - 0x40
      13'h1A55: dout  = 8'b00100000; // 6741 :  32 - 0x20
      13'h1A56: dout  = 8'b00011110; // 6742 :  30 - 0x1e
      13'h1A57: dout  = 8'b00000111; // 6743 :   7 - 0x7
      13'h1A58: dout  = 8'b00001101; // 6744 :  13 - 0xd
      13'h1A59: dout  = 8'b00011101; // 6745 :  29 - 0x1d
      13'h1A5A: dout  = 8'b00111101; // 6746 :  61 - 0x3d
      13'h1A5B: dout  = 8'b00111111; // 6747 :  63 - 0x3f
      13'h1A5C: dout  = 8'b00111111; // 6748 :  63 - 0x3f
      13'h1A5D: dout  = 8'b00011111; // 6749 :  31 - 0x1f
      13'h1A5E: dout  = 8'b00000001; // 6750 :   1 - 0x1
      13'h1A5F: dout  = 8'b00000000; // 6751 :   0 - 0x0
      13'h1A60: dout  = 8'b10000000; // 6752 : 128 - 0x80 -- Background 0xa6
      13'h1A61: dout  = 8'b11100000; // 6753 : 224 - 0xe0
      13'h1A62: dout  = 8'b00111000; // 6754 :  56 - 0x38
      13'h1A63: dout  = 8'b00100100; // 6755 :  36 - 0x24
      13'h1A64: dout  = 8'b00000100; // 6756 :   4 - 0x4
      13'h1A65: dout  = 8'b00001000; // 6757 :   8 - 0x8
      13'h1A66: dout  = 8'b00110000; // 6758 :  48 - 0x30
      13'h1A67: dout  = 8'b00100000; // 6759 :  32 - 0x20
      13'h1A68: dout  = 8'b00000000; // 6760 :   0 - 0x0
      13'h1A69: dout  = 8'b00000000; // 6761 :   0 - 0x0
      13'h1A6A: dout  = 8'b11100000; // 6762 : 224 - 0xe0
      13'h1A6B: dout  = 8'b11111000; // 6763 : 248 - 0xf8
      13'h1A6C: dout  = 8'b11111000; // 6764 : 248 - 0xf8
      13'h1A6D: dout  = 8'b11110000; // 6765 : 240 - 0xf0
      13'h1A6E: dout  = 8'b11000000; // 6766 : 192 - 0xc0
      13'h1A6F: dout  = 8'b11000000; // 6767 : 192 - 0xc0
      13'h1A70: dout  = 8'b00110000; // 6768 :  48 - 0x30 -- Background 0xa7
      13'h1A71: dout  = 8'b00001000; // 6769 :   8 - 0x8
      13'h1A72: dout  = 8'b00001000; // 6770 :   8 - 0x8
      13'h1A73: dout  = 8'b00110000; // 6771 :  48 - 0x30
      13'h1A74: dout  = 8'b00100000; // 6772 :  32 - 0x20
      13'h1A75: dout  = 8'b00100000; // 6773 :  32 - 0x20
      13'h1A76: dout  = 8'b00110000; // 6774 :  48 - 0x30
      13'h1A77: dout  = 8'b11110000; // 6775 : 240 - 0xf0
      13'h1A78: dout  = 8'b11000000; // 6776 : 192 - 0xc0
      13'h1A79: dout  = 8'b11110000; // 6777 : 240 - 0xf0
      13'h1A7A: dout  = 8'b11110000; // 6778 : 240 - 0xf0
      13'h1A7B: dout  = 8'b11000000; // 6779 : 192 - 0xc0
      13'h1A7C: dout  = 8'b11000000; // 6780 : 192 - 0xc0
      13'h1A7D: dout  = 8'b11000000; // 6781 : 192 - 0xc0
      13'h1A7E: dout  = 8'b11000000; // 6782 : 192 - 0xc0
      13'h1A7F: dout  = 8'b00000000; // 6783 :   0 - 0x0
      13'h1A80: dout  = 8'b11111111; // 6784 : 255 - 0xff -- Background 0xa8
      13'h1A81: dout  = 8'b11010010; // 6785 : 210 - 0xd2
      13'h1A82: dout  = 8'b11110100; // 6786 : 244 - 0xf4
      13'h1A83: dout  = 8'b11011000; // 6787 : 216 - 0xd8
      13'h1A84: dout  = 8'b11111000; // 6788 : 248 - 0xf8
      13'h1A85: dout  = 8'b11010100; // 6789 : 212 - 0xd4
      13'h1A86: dout  = 8'b11110010; // 6790 : 242 - 0xf2
      13'h1A87: dout  = 8'b11010001; // 6791 : 209 - 0xd1
      13'h1A88: dout  = 8'b00000000; // 6792 :   0 - 0x0
      13'h1A89: dout  = 8'b01100000; // 6793 :  96 - 0x60
      13'h1A8A: dout  = 8'b01100000; // 6794 :  96 - 0x60
      13'h1A8B: dout  = 8'b01100000; // 6795 :  96 - 0x60
      13'h1A8C: dout  = 8'b01100000; // 6796 :  96 - 0x60
      13'h1A8D: dout  = 8'b01100000; // 6797 :  96 - 0x60
      13'h1A8E: dout  = 8'b01100000; // 6798 :  96 - 0x60
      13'h1A8F: dout  = 8'b01100000; // 6799 :  96 - 0x60
      13'h1A90: dout  = 8'b11110001; // 6800 : 241 - 0xf1 -- Background 0xa9
      13'h1A91: dout  = 8'b11010010; // 6801 : 210 - 0xd2
      13'h1A92: dout  = 8'b11110100; // 6802 : 244 - 0xf4
      13'h1A93: dout  = 8'b11011000; // 6803 : 216 - 0xd8
      13'h1A94: dout  = 8'b11111000; // 6804 : 248 - 0xf8
      13'h1A95: dout  = 8'b11010100; // 6805 : 212 - 0xd4
      13'h1A96: dout  = 8'b11110010; // 6806 : 242 - 0xf2
      13'h1A97: dout  = 8'b11111111; // 6807 : 255 - 0xff
      13'h1A98: dout  = 8'b01100000; // 6808 :  96 - 0x60
      13'h1A99: dout  = 8'b01100000; // 6809 :  96 - 0x60
      13'h1A9A: dout  = 8'b01100000; // 6810 :  96 - 0x60
      13'h1A9B: dout  = 8'b01100000; // 6811 :  96 - 0x60
      13'h1A9C: dout  = 8'b01100000; // 6812 :  96 - 0x60
      13'h1A9D: dout  = 8'b01100000; // 6813 :  96 - 0x60
      13'h1A9E: dout  = 8'b01100000; // 6814 :  96 - 0x60
      13'h1A9F: dout  = 8'b00000000; // 6815 :   0 - 0x0
      13'h1AA0: dout  = 8'b11111111; // 6816 : 255 - 0xff -- Background 0xaa
      13'h1AA1: dout  = 8'b01000010; // 6817 :  66 - 0x42
      13'h1AA2: dout  = 8'b00100100; // 6818 :  36 - 0x24
      13'h1AA3: dout  = 8'b00011000; // 6819 :  24 - 0x18
      13'h1AA4: dout  = 8'b00011000; // 6820 :  24 - 0x18
      13'h1AA5: dout  = 8'b00100100; // 6821 :  36 - 0x24
      13'h1AA6: dout  = 8'b01000010; // 6822 :  66 - 0x42
      13'h1AA7: dout  = 8'b10000001; // 6823 : 129 - 0x81
      13'h1AA8: dout  = 8'b00000000; // 6824 :   0 - 0x0
      13'h1AA9: dout  = 8'b00000000; // 6825 :   0 - 0x0
      13'h1AAA: dout  = 8'b00000000; // 6826 :   0 - 0x0
      13'h1AAB: dout  = 8'b00000000; // 6827 :   0 - 0x0
      13'h1AAC: dout  = 8'b00000000; // 6828 :   0 - 0x0
      13'h1AAD: dout  = 8'b00000000; // 6829 :   0 - 0x0
      13'h1AAE: dout  = 8'b00000000; // 6830 :   0 - 0x0
      13'h1AAF: dout  = 8'b00000000; // 6831 :   0 - 0x0
      13'h1AB0: dout  = 8'b10000001; // 6832 : 129 - 0x81 -- Background 0xab
      13'h1AB1: dout  = 8'b01000010; // 6833 :  66 - 0x42
      13'h1AB2: dout  = 8'b00100100; // 6834 :  36 - 0x24
      13'h1AB3: dout  = 8'b00011000; // 6835 :  24 - 0x18
      13'h1AB4: dout  = 8'b00011000; // 6836 :  24 - 0x18
      13'h1AB5: dout  = 8'b00100100; // 6837 :  36 - 0x24
      13'h1AB6: dout  = 8'b01000010; // 6838 :  66 - 0x42
      13'h1AB7: dout  = 8'b11111111; // 6839 : 255 - 0xff
      13'h1AB8: dout  = 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout  = 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout  = 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout  = 8'b00000000; // 6843 :   0 - 0x0
      13'h1ABC: dout  = 8'b00000000; // 6844 :   0 - 0x0
      13'h1ABD: dout  = 8'b00000000; // 6845 :   0 - 0x0
      13'h1ABE: dout  = 8'b00000000; // 6846 :   0 - 0x0
      13'h1ABF: dout  = 8'b00000000; // 6847 :   0 - 0x0
      13'h1AC0: dout  = 8'b11111111; // 6848 : 255 - 0xff -- Background 0xac
      13'h1AC1: dout  = 8'b01001101; // 6849 :  77 - 0x4d
      13'h1AC2: dout  = 8'b00101111; // 6850 :  47 - 0x2f
      13'h1AC3: dout  = 8'b00011101; // 6851 :  29 - 0x1d
      13'h1AC4: dout  = 8'b00011111; // 6852 :  31 - 0x1f
      13'h1AC5: dout  = 8'b00101101; // 6853 :  45 - 0x2d
      13'h1AC6: dout  = 8'b01001111; // 6854 :  79 - 0x4f
      13'h1AC7: dout  = 8'b10001101; // 6855 : 141 - 0x8d
      13'h1AC8: dout  = 8'b00000000; // 6856 :   0 - 0x0
      13'h1AC9: dout  = 8'b00000110; // 6857 :   6 - 0x6
      13'h1ACA: dout  = 8'b00000110; // 6858 :   6 - 0x6
      13'h1ACB: dout  = 8'b00000110; // 6859 :   6 - 0x6
      13'h1ACC: dout  = 8'b00000110; // 6860 :   6 - 0x6
      13'h1ACD: dout  = 8'b00000110; // 6861 :   6 - 0x6
      13'h1ACE: dout  = 8'b00000110; // 6862 :   6 - 0x6
      13'h1ACF: dout  = 8'b00000110; // 6863 :   6 - 0x6
      13'h1AD0: dout  = 8'b10001111; // 6864 : 143 - 0x8f -- Background 0xad
      13'h1AD1: dout  = 8'b01001101; // 6865 :  77 - 0x4d
      13'h1AD2: dout  = 8'b00101111; // 6866 :  47 - 0x2f
      13'h1AD3: dout  = 8'b00011101; // 6867 :  29 - 0x1d
      13'h1AD4: dout  = 8'b00011111; // 6868 :  31 - 0x1f
      13'h1AD5: dout  = 8'b00101101; // 6869 :  45 - 0x2d
      13'h1AD6: dout  = 8'b01001111; // 6870 :  79 - 0x4f
      13'h1AD7: dout  = 8'b11111111; // 6871 : 255 - 0xff
      13'h1AD8: dout  = 8'b00000110; // 6872 :   6 - 0x6
      13'h1AD9: dout  = 8'b00000110; // 6873 :   6 - 0x6
      13'h1ADA: dout  = 8'b00000110; // 6874 :   6 - 0x6
      13'h1ADB: dout  = 8'b00000110; // 6875 :   6 - 0x6
      13'h1ADC: dout  = 8'b00000110; // 6876 :   6 - 0x6
      13'h1ADD: dout  = 8'b00000110; // 6877 :   6 - 0x6
      13'h1ADE: dout  = 8'b00000110; // 6878 :   6 - 0x6
      13'h1ADF: dout  = 8'b00000000; // 6879 :   0 - 0x0
      13'h1AE0: dout  = 8'b00000001; // 6880 :   1 - 0x1 -- Background 0xae
      13'h1AE1: dout  = 8'b00000011; // 6881 :   3 - 0x3
      13'h1AE2: dout  = 8'b00000110; // 6882 :   6 - 0x6
      13'h1AE3: dout  = 8'b00000111; // 6883 :   7 - 0x7
      13'h1AE4: dout  = 8'b00000111; // 6884 :   7 - 0x7
      13'h1AE5: dout  = 8'b00000111; // 6885 :   7 - 0x7
      13'h1AE6: dout  = 8'b00000110; // 6886 :   6 - 0x6
      13'h1AE7: dout  = 8'b00000111; // 6887 :   7 - 0x7
      13'h1AE8: dout  = 8'b00000000; // 6888 :   0 - 0x0
      13'h1AE9: dout  = 8'b00000001; // 6889 :   1 - 0x1
      13'h1AEA: dout  = 8'b00000011; // 6890 :   3 - 0x3
      13'h1AEB: dout  = 8'b00000010; // 6891 :   2 - 0x2
      13'h1AEC: dout  = 8'b00000010; // 6892 :   2 - 0x2
      13'h1AED: dout  = 8'b00000000; // 6893 :   0 - 0x0
      13'h1AEE: dout  = 8'b00000011; // 6894 :   3 - 0x3
      13'h1AEF: dout  = 8'b00000010; // 6895 :   2 - 0x2
      13'h1AF0: dout  = 8'b00000110; // 6896 :   6 - 0x6 -- Background 0xaf
      13'h1AF1: dout  = 8'b00000110; // 6897 :   6 - 0x6
      13'h1AF2: dout  = 8'b00001110; // 6898 :  14 - 0xe
      13'h1AF3: dout  = 8'b00001111; // 6899 :  15 - 0xf
      13'h1AF4: dout  = 8'b00001110; // 6900 :  14 - 0xe
      13'h1AF5: dout  = 8'b00011010; // 6901 :  26 - 0x1a
      13'h1AF6: dout  = 8'b00011011; // 6902 :  27 - 0x1b
      13'h1AF7: dout  = 8'b00001111; // 6903 :  15 - 0xf
      13'h1AF8: dout  = 8'b00000001; // 6904 :   1 - 0x1
      13'h1AF9: dout  = 8'b00000011; // 6905 :   3 - 0x3
      13'h1AFA: dout  = 8'b00000101; // 6906 :   5 - 0x5
      13'h1AFB: dout  = 8'b00000100; // 6907 :   4 - 0x4
      13'h1AFC: dout  = 8'b00000101; // 6908 :   5 - 0x5
      13'h1AFD: dout  = 8'b00001101; // 6909 :  13 - 0xd
      13'h1AFE: dout  = 8'b00001100; // 6910 :  12 - 0xc
      13'h1AFF: dout  = 8'b00000001; // 6911 :   1 - 0x1
      13'h1B00: dout  = 8'b00000000; // 6912 :   0 - 0x0 -- Background 0xb0
      13'h1B01: dout  = 8'b11000000; // 6913 : 192 - 0xc0
      13'h1B02: dout  = 8'b11110000; // 6914 : 240 - 0xf0
      13'h1B03: dout  = 8'b10001000; // 6915 : 136 - 0x88
      13'h1B04: dout  = 8'b00010100; // 6916 :  20 - 0x14
      13'h1B05: dout  = 8'b01101000; // 6917 : 104 - 0x68
      13'h1B06: dout  = 8'b10101000; // 6918 : 168 - 0xa8
      13'h1B07: dout  = 8'b00101100; // 6919 :  44 - 0x2c
      13'h1B08: dout  = 8'b00000000; // 6920 :   0 - 0x0
      13'h1B09: dout  = 8'b00000000; // 6921 :   0 - 0x0
      13'h1B0A: dout  = 8'b01000000; // 6922 :  64 - 0x40
      13'h1B0B: dout  = 8'b11110000; // 6923 : 240 - 0xf0
      13'h1B0C: dout  = 8'b11101000; // 6924 : 232 - 0xe8
      13'h1B0D: dout  = 8'b10010000; // 6925 : 144 - 0x90
      13'h1B0E: dout  = 8'b01010000; // 6926 :  80 - 0x50
      13'h1B0F: dout  = 8'b11010000; // 6927 : 208 - 0xd0
      13'h1B10: dout  = 8'b00000100; // 6928 :   4 - 0x4 -- Background 0xb1
      13'h1B11: dout  = 8'b00111000; // 6929 :  56 - 0x38
      13'h1B12: dout  = 8'b00010000; // 6930 :  16 - 0x10
      13'h1B13: dout  = 8'b10100000; // 6931 : 160 - 0xa0
      13'h1B14: dout  = 8'b01100000; // 6932 :  96 - 0x60
      13'h1B15: dout  = 8'b00100000; // 6933 :  32 - 0x20
      13'h1B16: dout  = 8'b00010000; // 6934 :  16 - 0x10
      13'h1B17: dout  = 8'b10001000; // 6935 : 136 - 0x88
      13'h1B18: dout  = 8'b11111000; // 6936 : 248 - 0xf8
      13'h1B19: dout  = 8'b11000000; // 6937 : 192 - 0xc0
      13'h1B1A: dout  = 8'b11100000; // 6938 : 224 - 0xe0
      13'h1B1B: dout  = 8'b01000000; // 6939 :  64 - 0x40
      13'h1B1C: dout  = 8'b10000000; // 6940 : 128 - 0x80
      13'h1B1D: dout  = 8'b11000000; // 6941 : 192 - 0xc0
      13'h1B1E: dout  = 8'b11100000; // 6942 : 224 - 0xe0
      13'h1B1F: dout  = 8'b01110000; // 6943 : 112 - 0x70
      13'h1B20: dout  = 8'b00001111; // 6944 :  15 - 0xf -- Background 0xb2
      13'h1B21: dout  = 8'b00011011; // 6945 :  27 - 0x1b
      13'h1B22: dout  = 8'b00011011; // 6946 :  27 - 0x1b
      13'h1B23: dout  = 8'b00001110; // 6947 :  14 - 0xe
      13'h1B24: dout  = 8'b00000110; // 6948 :   6 - 0x6
      13'h1B25: dout  = 8'b00001100; // 6949 :  12 - 0xc
      13'h1B26: dout  = 8'b00001100; // 6950 :  12 - 0xc
      13'h1B27: dout  = 8'b00111111; // 6951 :  63 - 0x3f
      13'h1B28: dout  = 8'b00000001; // 6952 :   1 - 0x1
      13'h1B29: dout  = 8'b00001101; // 6953 :  13 - 0xd
      13'h1B2A: dout  = 8'b00001101; // 6954 :  13 - 0xd
      13'h1B2B: dout  = 8'b00000011; // 6955 :   3 - 0x3
      13'h1B2C: dout  = 8'b00000011; // 6956 :   3 - 0x3
      13'h1B2D: dout  = 8'b00000111; // 6957 :   7 - 0x7
      13'h1B2E: dout  = 8'b00000111; // 6958 :   7 - 0x7
      13'h1B2F: dout  = 8'b00000000; // 6959 :   0 - 0x0
      13'h1B30: dout  = 8'b01111111; // 6960 : 127 - 0x7f -- Background 0xb3
      13'h1B31: dout  = 8'b01100000; // 6961 :  96 - 0x60
      13'h1B32: dout  = 8'b01100000; // 6962 :  96 - 0x60
      13'h1B33: dout  = 8'b01100000; // 6963 :  96 - 0x60
      13'h1B34: dout  = 8'b01100000; // 6964 :  96 - 0x60
      13'h1B35: dout  = 8'b01100000; // 6965 :  96 - 0x60
      13'h1B36: dout  = 8'b01101010; // 6966 : 106 - 0x6a
      13'h1B37: dout  = 8'b01111111; // 6967 : 127 - 0x7f
      13'h1B38: dout  = 8'b00111111; // 6968 :  63 - 0x3f
      13'h1B39: dout  = 8'b00111111; // 6969 :  63 - 0x3f
      13'h1B3A: dout  = 8'b00111111; // 6970 :  63 - 0x3f
      13'h1B3B: dout  = 8'b00111111; // 6971 :  63 - 0x3f
      13'h1B3C: dout  = 8'b00111111; // 6972 :  63 - 0x3f
      13'h1B3D: dout  = 8'b00111111; // 6973 :  63 - 0x3f
      13'h1B3E: dout  = 8'b00110101; // 6974 :  53 - 0x35
      13'h1B3F: dout  = 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout  = 8'b01001000; // 6976 :  72 - 0x48 -- Background 0xb4
      13'h1B41: dout  = 8'b00110000; // 6977 :  48 - 0x30
      13'h1B42: dout  = 8'b00010000; // 6978 :  16 - 0x10
      13'h1B43: dout  = 8'b00010000; // 6979 :  16 - 0x10
      13'h1B44: dout  = 8'b00001000; // 6980 :   8 - 0x8
      13'h1B45: dout  = 8'b00001000; // 6981 :   8 - 0x8
      13'h1B46: dout  = 8'b00001000; // 6982 :   8 - 0x8
      13'h1B47: dout  = 8'b11111100; // 6983 : 252 - 0xfc
      13'h1B48: dout  = 8'b10110000; // 6984 : 176 - 0xb0
      13'h1B49: dout  = 8'b11000000; // 6985 : 192 - 0xc0
      13'h1B4A: dout  = 8'b11100000; // 6986 : 224 - 0xe0
      13'h1B4B: dout  = 8'b11100000; // 6987 : 224 - 0xe0
      13'h1B4C: dout  = 8'b11110000; // 6988 : 240 - 0xf0
      13'h1B4D: dout  = 8'b11110000; // 6989 : 240 - 0xf0
      13'h1B4E: dout  = 8'b11110000; // 6990 : 240 - 0xf0
      13'h1B4F: dout  = 8'b00000000; // 6991 :   0 - 0x0
      13'h1B50: dout  = 8'b11111110; // 6992 : 254 - 0xfe -- Background 0xb5
      13'h1B51: dout  = 8'b00000110; // 6993 :   6 - 0x6
      13'h1B52: dout  = 8'b00000010; // 6994 :   2 - 0x2
      13'h1B53: dout  = 8'b00000110; // 6995 :   6 - 0x6
      13'h1B54: dout  = 8'b00000010; // 6996 :   2 - 0x2
      13'h1B55: dout  = 8'b00000110; // 6997 :   6 - 0x6
      13'h1B56: dout  = 8'b10101010; // 6998 : 170 - 0xaa
      13'h1B57: dout  = 8'b11111110; // 6999 : 254 - 0xfe
      13'h1B58: dout  = 8'b11111100; // 7000 : 252 - 0xfc
      13'h1B59: dout  = 8'b11111000; // 7001 : 248 - 0xf8
      13'h1B5A: dout  = 8'b11111100; // 7002 : 252 - 0xfc
      13'h1B5B: dout  = 8'b11111000; // 7003 : 248 - 0xf8
      13'h1B5C: dout  = 8'b11111100; // 7004 : 252 - 0xfc
      13'h1B5D: dout  = 8'b11111000; // 7005 : 248 - 0xf8
      13'h1B5E: dout  = 8'b01010100; // 7006 :  84 - 0x54
      13'h1B5F: dout  = 8'b00000000; // 7007 :   0 - 0x0
      13'h1B60: dout  = 8'b11111111; // 7008 : 255 - 0xff -- Background 0xb6
      13'h1B61: dout  = 8'b10000000; // 7009 : 128 - 0x80
      13'h1B62: dout  = 8'b10000000; // 7010 : 128 - 0x80
      13'h1B63: dout  = 8'b10000000; // 7011 : 128 - 0x80
      13'h1B64: dout  = 8'b10000000; // 7012 : 128 - 0x80
      13'h1B65: dout  = 8'b10000000; // 7013 : 128 - 0x80
      13'h1B66: dout  = 8'b10010101; // 7014 : 149 - 0x95
      13'h1B67: dout  = 8'b11111111; // 7015 : 255 - 0xff
      13'h1B68: dout  = 8'b00000000; // 7016 :   0 - 0x0
      13'h1B69: dout  = 8'b01111111; // 7017 : 127 - 0x7f
      13'h1B6A: dout  = 8'b01111111; // 7018 : 127 - 0x7f
      13'h1B6B: dout  = 8'b01111111; // 7019 : 127 - 0x7f
      13'h1B6C: dout  = 8'b01111111; // 7020 : 127 - 0x7f
      13'h1B6D: dout  = 8'b01111111; // 7021 : 127 - 0x7f
      13'h1B6E: dout  = 8'b01101010; // 7022 : 106 - 0x6a
      13'h1B6F: dout  = 8'b00000000; // 7023 :   0 - 0x0
      13'h1B70: dout  = 8'b11111111; // 7024 : 255 - 0xff -- Background 0xb7
      13'h1B71: dout  = 8'b10000100; // 7025 : 132 - 0x84
      13'h1B72: dout  = 8'b10001100; // 7026 : 140 - 0x8c
      13'h1B73: dout  = 8'b10000100; // 7027 : 132 - 0x84
      13'h1B74: dout  = 8'b10001100; // 7028 : 140 - 0x8c
      13'h1B75: dout  = 8'b10000100; // 7029 : 132 - 0x84
      13'h1B76: dout  = 8'b10101100; // 7030 : 172 - 0xac
      13'h1B77: dout  = 8'b11111111; // 7031 : 255 - 0xff
      13'h1B78: dout  = 8'b00000000; // 7032 :   0 - 0x0
      13'h1B79: dout  = 8'b01111011; // 7033 : 123 - 0x7b
      13'h1B7A: dout  = 8'b01110011; // 7034 : 115 - 0x73
      13'h1B7B: dout  = 8'b01111011; // 7035 : 123 - 0x7b
      13'h1B7C: dout  = 8'b01110011; // 7036 : 115 - 0x73
      13'h1B7D: dout  = 8'b01111011; // 7037 : 123 - 0x7b
      13'h1B7E: dout  = 8'b01010011; // 7038 :  83 - 0x53
      13'h1B7F: dout  = 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout  = 8'b11111111; // 7040 : 255 - 0xff -- Background 0xb8
      13'h1B81: dout  = 8'b00100001; // 7041 :  33 - 0x21
      13'h1B82: dout  = 8'b01100001; // 7042 :  97 - 0x61
      13'h1B83: dout  = 8'b00100011; // 7043 :  35 - 0x23
      13'h1B84: dout  = 8'b01100001; // 7044 :  97 - 0x61
      13'h1B85: dout  = 8'b00100011; // 7045 :  35 - 0x23
      13'h1B86: dout  = 8'b01100101; // 7046 : 101 - 0x65
      13'h1B87: dout  = 8'b11111111; // 7047 : 255 - 0xff
      13'h1B88: dout  = 8'b00000000; // 7048 :   0 - 0x0
      13'h1B89: dout  = 8'b11011110; // 7049 : 222 - 0xde
      13'h1B8A: dout  = 8'b10011110; // 7050 : 158 - 0x9e
      13'h1B8B: dout  = 8'b11011100; // 7051 : 220 - 0xdc
      13'h1B8C: dout  = 8'b10011110; // 7052 : 158 - 0x9e
      13'h1B8D: dout  = 8'b11011100; // 7053 : 220 - 0xdc
      13'h1B8E: dout  = 8'b10011010; // 7054 : 154 - 0x9a
      13'h1B8F: dout  = 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout  = 8'b11111111; // 7056 : 255 - 0xff -- Background 0xb9
      13'h1B91: dout  = 8'b00000001; // 7057 :   1 - 0x1
      13'h1B92: dout  = 8'b00000011; // 7058 :   3 - 0x3
      13'h1B93: dout  = 8'b00000001; // 7059 :   1 - 0x1
      13'h1B94: dout  = 8'b00000011; // 7060 :   3 - 0x3
      13'h1B95: dout  = 8'b00000001; // 7061 :   1 - 0x1
      13'h1B96: dout  = 8'b10101011; // 7062 : 171 - 0xab
      13'h1B97: dout  = 8'b11111111; // 7063 : 255 - 0xff
      13'h1B98: dout  = 8'b00000000; // 7064 :   0 - 0x0
      13'h1B99: dout  = 8'b11111110; // 7065 : 254 - 0xfe
      13'h1B9A: dout  = 8'b11111100; // 7066 : 252 - 0xfc
      13'h1B9B: dout  = 8'b11111110; // 7067 : 254 - 0xfe
      13'h1B9C: dout  = 8'b11111100; // 7068 : 252 - 0xfc
      13'h1B9D: dout  = 8'b11111110; // 7069 : 254 - 0xfe
      13'h1B9E: dout  = 8'b01010100; // 7070 :  84 - 0x54
      13'h1B9F: dout  = 8'b00000000; // 7071 :   0 - 0x0
      13'h1BA0: dout  = 8'b11111111; // 7072 : 255 - 0xff -- Background 0xba
      13'h1BA1: dout  = 8'b11010101; // 7073 : 213 - 0xd5
      13'h1BA2: dout  = 8'b10101010; // 7074 : 170 - 0xaa
      13'h1BA3: dout  = 8'b11111111; // 7075 : 255 - 0xff
      13'h1BA4: dout  = 8'b10000000; // 7076 : 128 - 0x80
      13'h1BA5: dout  = 8'b10000000; // 7077 : 128 - 0x80
      13'h1BA6: dout  = 8'b10010101; // 7078 : 149 - 0x95
      13'h1BA7: dout  = 8'b11111111; // 7079 : 255 - 0xff
      13'h1BA8: dout  = 8'b00000000; // 7080 :   0 - 0x0
      13'h1BA9: dout  = 8'b01111111; // 7081 : 127 - 0x7f
      13'h1BAA: dout  = 8'b01111111; // 7082 : 127 - 0x7f
      13'h1BAB: dout  = 8'b00000000; // 7083 :   0 - 0x0
      13'h1BAC: dout  = 8'b01111111; // 7084 : 127 - 0x7f
      13'h1BAD: dout  = 8'b01111111; // 7085 : 127 - 0x7f
      13'h1BAE: dout  = 8'b01101010; // 7086 : 106 - 0x6a
      13'h1BAF: dout  = 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout  = 8'b00000000; // 7088 :   0 - 0x0 -- Background 0xbb
      13'h1BB1: dout  = 8'b00000000; // 7089 :   0 - 0x0
      13'h1BB2: dout  = 8'b00000000; // 7090 :   0 - 0x0
      13'h1BB3: dout  = 8'b00000000; // 7091 :   0 - 0x0
      13'h1BB4: dout  = 8'b00000000; // 7092 :   0 - 0x0
      13'h1BB5: dout  = 8'b00000000; // 7093 :   0 - 0x0
      13'h1BB6: dout  = 8'b00000000; // 7094 :   0 - 0x0
      13'h1BB7: dout  = 8'b00000000; // 7095 :   0 - 0x0
      13'h1BB8: dout  = 8'b00000000; // 7096 :   0 - 0x0
      13'h1BB9: dout  = 8'b00000000; // 7097 :   0 - 0x0
      13'h1BBA: dout  = 8'b00000000; // 7098 :   0 - 0x0
      13'h1BBB: dout  = 8'b00000000; // 7099 :   0 - 0x0
      13'h1BBC: dout  = 8'b00000000; // 7100 :   0 - 0x0
      13'h1BBD: dout  = 8'b00000000; // 7101 :   0 - 0x0
      13'h1BBE: dout  = 8'b00000000; // 7102 :   0 - 0x0
      13'h1BBF: dout  = 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout  = 8'b11111111; // 7104 : 255 - 0xff -- Background 0xbc
      13'h1BC1: dout  = 8'b01010101; // 7105 :  85 - 0x55
      13'h1BC2: dout  = 8'b10101011; // 7106 : 171 - 0xab
      13'h1BC3: dout  = 8'b11111111; // 7107 : 255 - 0xff
      13'h1BC4: dout  = 8'b01100001; // 7108 :  97 - 0x61
      13'h1BC5: dout  = 8'b00100011; // 7109 :  35 - 0x23
      13'h1BC6: dout  = 8'b01100101; // 7110 : 101 - 0x65
      13'h1BC7: dout  = 8'b11111111; // 7111 : 255 - 0xff
      13'h1BC8: dout  = 8'b00000000; // 7112 :   0 - 0x0
      13'h1BC9: dout  = 8'b11111110; // 7113 : 254 - 0xfe
      13'h1BCA: dout  = 8'b11111110; // 7114 : 254 - 0xfe
      13'h1BCB: dout  = 8'b00000000; // 7115 :   0 - 0x0
      13'h1BCC: dout  = 8'b10011110; // 7116 : 158 - 0x9e
      13'h1BCD: dout  = 8'b11011100; // 7117 : 220 - 0xdc
      13'h1BCE: dout  = 8'b10011010; // 7118 : 154 - 0x9a
      13'h1BCF: dout  = 8'b00000000; // 7119 :   0 - 0x0
      13'h1BD0: dout  = 8'b00000000; // 7120 :   0 - 0x0 -- Background 0xbd
      13'h1BD1: dout  = 8'b00000000; // 7121 :   0 - 0x0
      13'h1BD2: dout  = 8'b00000000; // 7122 :   0 - 0x0
      13'h1BD3: dout  = 8'b00000000; // 7123 :   0 - 0x0
      13'h1BD4: dout  = 8'b00000000; // 7124 :   0 - 0x0
      13'h1BD5: dout  = 8'b00000000; // 7125 :   0 - 0x0
      13'h1BD6: dout  = 8'b00000000; // 7126 :   0 - 0x0
      13'h1BD7: dout  = 8'b00000000; // 7127 :   0 - 0x0
      13'h1BD8: dout  = 8'b00000000; // 7128 :   0 - 0x0
      13'h1BD9: dout  = 8'b00000000; // 7129 :   0 - 0x0
      13'h1BDA: dout  = 8'b00000000; // 7130 :   0 - 0x0
      13'h1BDB: dout  = 8'b00000000; // 7131 :   0 - 0x0
      13'h1BDC: dout  = 8'b00000000; // 7132 :   0 - 0x0
      13'h1BDD: dout  = 8'b00000000; // 7133 :   0 - 0x0
      13'h1BDE: dout  = 8'b00000000; // 7134 :   0 - 0x0
      13'h1BDF: dout  = 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout  = 8'b00000000; // 7136 :   0 - 0x0 -- Background 0xbe
      13'h1BE1: dout  = 8'b00000000; // 7137 :   0 - 0x0
      13'h1BE2: dout  = 8'b00000000; // 7138 :   0 - 0x0
      13'h1BE3: dout  = 8'b00000000; // 7139 :   0 - 0x0
      13'h1BE4: dout  = 8'b00000000; // 7140 :   0 - 0x0
      13'h1BE5: dout  = 8'b00000000; // 7141 :   0 - 0x0
      13'h1BE6: dout  = 8'b00000000; // 7142 :   0 - 0x0
      13'h1BE7: dout  = 8'b00000000; // 7143 :   0 - 0x0
      13'h1BE8: dout  = 8'b00000000; // 7144 :   0 - 0x0
      13'h1BE9: dout  = 8'b00000000; // 7145 :   0 - 0x0
      13'h1BEA: dout  = 8'b00000000; // 7146 :   0 - 0x0
      13'h1BEB: dout  = 8'b00000000; // 7147 :   0 - 0x0
      13'h1BEC: dout  = 8'b00000000; // 7148 :   0 - 0x0
      13'h1BED: dout  = 8'b00000000; // 7149 :   0 - 0x0
      13'h1BEE: dout  = 8'b00000000; // 7150 :   0 - 0x0
      13'h1BEF: dout  = 8'b00000000; // 7151 :   0 - 0x0
      13'h1BF0: dout  = 8'b00000000; // 7152 :   0 - 0x0 -- Background 0xbf
      13'h1BF1: dout  = 8'b00000000; // 7153 :   0 - 0x0
      13'h1BF2: dout  = 8'b00000000; // 7154 :   0 - 0x0
      13'h1BF3: dout  = 8'b00000000; // 7155 :   0 - 0x0
      13'h1BF4: dout  = 8'b00000000; // 7156 :   0 - 0x0
      13'h1BF5: dout  = 8'b00000000; // 7157 :   0 - 0x0
      13'h1BF6: dout  = 8'b00000000; // 7158 :   0 - 0x0
      13'h1BF7: dout  = 8'b00000000; // 7159 :   0 - 0x0
      13'h1BF8: dout  = 8'b00000000; // 7160 :   0 - 0x0
      13'h1BF9: dout  = 8'b00000000; // 7161 :   0 - 0x0
      13'h1BFA: dout  = 8'b00000000; // 7162 :   0 - 0x0
      13'h1BFB: dout  = 8'b00000000; // 7163 :   0 - 0x0
      13'h1BFC: dout  = 8'b00000000; // 7164 :   0 - 0x0
      13'h1BFD: dout  = 8'b00000000; // 7165 :   0 - 0x0
      13'h1BFE: dout  = 8'b00000000; // 7166 :   0 - 0x0
      13'h1BFF: dout  = 8'b00000000; // 7167 :   0 - 0x0
      13'h1C00: dout  = 8'b00000000; // 7168 :   0 - 0x0 -- Background 0xc0
      13'h1C01: dout  = 8'b00000000; // 7169 :   0 - 0x0
      13'h1C02: dout  = 8'b00000000; // 7170 :   0 - 0x0
      13'h1C03: dout  = 8'b00000000; // 7171 :   0 - 0x0
      13'h1C04: dout  = 8'b00000000; // 7172 :   0 - 0x0
      13'h1C05: dout  = 8'b00000000; // 7173 :   0 - 0x0
      13'h1C06: dout  = 8'b00000000; // 7174 :   0 - 0x0
      13'h1C07: dout  = 8'b00000000; // 7175 :   0 - 0x0
      13'h1C08: dout  = 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout  = 8'b00000000; // 7177 :   0 - 0x0
      13'h1C0A: dout  = 8'b00000000; // 7178 :   0 - 0x0
      13'h1C0B: dout  = 8'b00000000; // 7179 :   0 - 0x0
      13'h1C0C: dout  = 8'b00000000; // 7180 :   0 - 0x0
      13'h1C0D: dout  = 8'b00000000; // 7181 :   0 - 0x0
      13'h1C0E: dout  = 8'b00000000; // 7182 :   0 - 0x0
      13'h1C0F: dout  = 8'b00000000; // 7183 :   0 - 0x0
      13'h1C10: dout  = 8'b00000000; // 7184 :   0 - 0x0 -- Background 0xc1
      13'h1C11: dout  = 8'b00000000; // 7185 :   0 - 0x0
      13'h1C12: dout  = 8'b00000000; // 7186 :   0 - 0x0
      13'h1C13: dout  = 8'b00000000; // 7187 :   0 - 0x0
      13'h1C14: dout  = 8'b00000000; // 7188 :   0 - 0x0
      13'h1C15: dout  = 8'b00000000; // 7189 :   0 - 0x0
      13'h1C16: dout  = 8'b00000000; // 7190 :   0 - 0x0
      13'h1C17: dout  = 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout  = 8'b00000000; // 7192 :   0 - 0x0
      13'h1C19: dout  = 8'b00000000; // 7193 :   0 - 0x0
      13'h1C1A: dout  = 8'b00000000; // 7194 :   0 - 0x0
      13'h1C1B: dout  = 8'b00000000; // 7195 :   0 - 0x0
      13'h1C1C: dout  = 8'b00000000; // 7196 :   0 - 0x0
      13'h1C1D: dout  = 8'b00000000; // 7197 :   0 - 0x0
      13'h1C1E: dout  = 8'b00000000; // 7198 :   0 - 0x0
      13'h1C1F: dout  = 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout  = 8'b00000000; // 7200 :   0 - 0x0 -- Background 0xc2
      13'h1C21: dout  = 8'b00000000; // 7201 :   0 - 0x0
      13'h1C22: dout  = 8'b00000000; // 7202 :   0 - 0x0
      13'h1C23: dout  = 8'b00000000; // 7203 :   0 - 0x0
      13'h1C24: dout  = 8'b00000000; // 7204 :   0 - 0x0
      13'h1C25: dout  = 8'b00000000; // 7205 :   0 - 0x0
      13'h1C26: dout  = 8'b00000000; // 7206 :   0 - 0x0
      13'h1C27: dout  = 8'b00000000; // 7207 :   0 - 0x0
      13'h1C28: dout  = 8'b00000000; // 7208 :   0 - 0x0
      13'h1C29: dout  = 8'b00000000; // 7209 :   0 - 0x0
      13'h1C2A: dout  = 8'b00000000; // 7210 :   0 - 0x0
      13'h1C2B: dout  = 8'b00000000; // 7211 :   0 - 0x0
      13'h1C2C: dout  = 8'b00000000; // 7212 :   0 - 0x0
      13'h1C2D: dout  = 8'b00000000; // 7213 :   0 - 0x0
      13'h1C2E: dout  = 8'b00000000; // 7214 :   0 - 0x0
      13'h1C2F: dout  = 8'b00000000; // 7215 :   0 - 0x0
      13'h1C30: dout  = 8'b00000000; // 7216 :   0 - 0x0 -- Background 0xc3
      13'h1C31: dout  = 8'b00000000; // 7217 :   0 - 0x0
      13'h1C32: dout  = 8'b00000000; // 7218 :   0 - 0x0
      13'h1C33: dout  = 8'b00000000; // 7219 :   0 - 0x0
      13'h1C34: dout  = 8'b00000000; // 7220 :   0 - 0x0
      13'h1C35: dout  = 8'b00000000; // 7221 :   0 - 0x0
      13'h1C36: dout  = 8'b00000000; // 7222 :   0 - 0x0
      13'h1C37: dout  = 8'b00000000; // 7223 :   0 - 0x0
      13'h1C38: dout  = 8'b00000000; // 7224 :   0 - 0x0
      13'h1C39: dout  = 8'b00000000; // 7225 :   0 - 0x0
      13'h1C3A: dout  = 8'b00000000; // 7226 :   0 - 0x0
      13'h1C3B: dout  = 8'b00000000; // 7227 :   0 - 0x0
      13'h1C3C: dout  = 8'b00000000; // 7228 :   0 - 0x0
      13'h1C3D: dout  = 8'b00000000; // 7229 :   0 - 0x0
      13'h1C3E: dout  = 8'b00000000; // 7230 :   0 - 0x0
      13'h1C3F: dout  = 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout  = 8'b00000000; // 7232 :   0 - 0x0 -- Background 0xc4
      13'h1C41: dout  = 8'b00000000; // 7233 :   0 - 0x0
      13'h1C42: dout  = 8'b00000000; // 7234 :   0 - 0x0
      13'h1C43: dout  = 8'b00000000; // 7235 :   0 - 0x0
      13'h1C44: dout  = 8'b00000000; // 7236 :   0 - 0x0
      13'h1C45: dout  = 8'b00000000; // 7237 :   0 - 0x0
      13'h1C46: dout  = 8'b00000000; // 7238 :   0 - 0x0
      13'h1C47: dout  = 8'b00000000; // 7239 :   0 - 0x0
      13'h1C48: dout  = 8'b00000000; // 7240 :   0 - 0x0
      13'h1C49: dout  = 8'b00000000; // 7241 :   0 - 0x0
      13'h1C4A: dout  = 8'b00000000; // 7242 :   0 - 0x0
      13'h1C4B: dout  = 8'b00000000; // 7243 :   0 - 0x0
      13'h1C4C: dout  = 8'b00000000; // 7244 :   0 - 0x0
      13'h1C4D: dout  = 8'b00000000; // 7245 :   0 - 0x0
      13'h1C4E: dout  = 8'b00000000; // 7246 :   0 - 0x0
      13'h1C4F: dout  = 8'b00000000; // 7247 :   0 - 0x0
      13'h1C50: dout  = 8'b00000000; // 7248 :   0 - 0x0 -- Background 0xc5
      13'h1C51: dout  = 8'b00000000; // 7249 :   0 - 0x0
      13'h1C52: dout  = 8'b00000001; // 7250 :   1 - 0x1
      13'h1C53: dout  = 8'b00000110; // 7251 :   6 - 0x6
      13'h1C54: dout  = 8'b00001010; // 7252 :  10 - 0xa
      13'h1C55: dout  = 8'b00010100; // 7253 :  20 - 0x14
      13'h1C56: dout  = 8'b00010000; // 7254 :  16 - 0x10
      13'h1C57: dout  = 8'b00101000; // 7255 :  40 - 0x28
      13'h1C58: dout  = 8'b00000000; // 7256 :   0 - 0x0
      13'h1C59: dout  = 8'b00000000; // 7257 :   0 - 0x0
      13'h1C5A: dout  = 8'b00000000; // 7258 :   0 - 0x0
      13'h1C5B: dout  = 8'b00000001; // 7259 :   1 - 0x1
      13'h1C5C: dout  = 8'b00000111; // 7260 :   7 - 0x7
      13'h1C5D: dout  = 8'b00001111; // 7261 :  15 - 0xf
      13'h1C5E: dout  = 8'b00001111; // 7262 :  15 - 0xf
      13'h1C5F: dout  = 8'b00011111; // 7263 :  31 - 0x1f
      13'h1C60: dout  = 8'b00011111; // 7264 :  31 - 0x1f -- Background 0xc6
      13'h1C61: dout  = 8'b01100000; // 7265 :  96 - 0x60
      13'h1C62: dout  = 8'b10100000; // 7266 : 160 - 0xa0
      13'h1C63: dout  = 8'b01000000; // 7267 :  64 - 0x40
      13'h1C64: dout  = 8'b00000000; // 7268 :   0 - 0x0
      13'h1C65: dout  = 8'b00000000; // 7269 :   0 - 0x0
      13'h1C66: dout  = 8'b00000000; // 7270 :   0 - 0x0
      13'h1C67: dout  = 8'b00000000; // 7271 :   0 - 0x0
      13'h1C68: dout  = 8'b00000000; // 7272 :   0 - 0x0
      13'h1C69: dout  = 8'b00011111; // 7273 :  31 - 0x1f
      13'h1C6A: dout  = 8'b01111111; // 7274 : 127 - 0x7f
      13'h1C6B: dout  = 8'b11111111; // 7275 : 255 - 0xff
      13'h1C6C: dout  = 8'b11111111; // 7276 : 255 - 0xff
      13'h1C6D: dout  = 8'b11111111; // 7277 : 255 - 0xff
      13'h1C6E: dout  = 8'b11111111; // 7278 : 255 - 0xff
      13'h1C6F: dout  = 8'b11111111; // 7279 : 255 - 0xff
      13'h1C70: dout  = 8'b00110000; // 7280 :  48 - 0x30 -- Background 0xc7
      13'h1C71: dout  = 8'b01000000; // 7281 :  64 - 0x40
      13'h1C72: dout  = 8'b01100000; // 7282 :  96 - 0x60
      13'h1C73: dout  = 8'b11000000; // 7283 : 192 - 0xc0
      13'h1C74: dout  = 8'b10000000; // 7284 : 128 - 0x80
      13'h1C75: dout  = 8'b10100000; // 7285 : 160 - 0xa0
      13'h1C76: dout  = 8'b11000000; // 7286 : 192 - 0xc0
      13'h1C77: dout  = 8'b10000000; // 7287 : 128 - 0x80
      13'h1C78: dout  = 8'b00011111; // 7288 :  31 - 0x1f
      13'h1C79: dout  = 8'b00111111; // 7289 :  63 - 0x3f
      13'h1C7A: dout  = 8'b00111111; // 7290 :  63 - 0x3f
      13'h1C7B: dout  = 8'b01111111; // 7291 : 127 - 0x7f
      13'h1C7C: dout  = 8'b01111111; // 7292 : 127 - 0x7f
      13'h1C7D: dout  = 8'b01111111; // 7293 : 127 - 0x7f
      13'h1C7E: dout  = 8'b01111111; // 7294 : 127 - 0x7f
      13'h1C7F: dout  = 8'b01111111; // 7295 : 127 - 0x7f
      13'h1C80: dout  = 8'b11111111; // 7296 : 255 - 0xff -- Background 0xc8
      13'h1C81: dout  = 8'b00000000; // 7297 :   0 - 0x0
      13'h1C82: dout  = 8'b00000000; // 7298 :   0 - 0x0
      13'h1C83: dout  = 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout  = 8'b00000000; // 7300 :   0 - 0x0
      13'h1C85: dout  = 8'b00000000; // 7301 :   0 - 0x0
      13'h1C86: dout  = 8'b00000000; // 7302 :   0 - 0x0
      13'h1C87: dout  = 8'b00000000; // 7303 :   0 - 0x0
      13'h1C88: dout  = 8'b00000000; // 7304 :   0 - 0x0
      13'h1C89: dout  = 8'b11111111; // 7305 : 255 - 0xff
      13'h1C8A: dout  = 8'b11111111; // 7306 : 255 - 0xff
      13'h1C8B: dout  = 8'b11111111; // 7307 : 255 - 0xff
      13'h1C8C: dout  = 8'b11111111; // 7308 : 255 - 0xff
      13'h1C8D: dout  = 8'b11111111; // 7309 : 255 - 0xff
      13'h1C8E: dout  = 8'b11111111; // 7310 : 255 - 0xff
      13'h1C8F: dout  = 8'b11111111; // 7311 : 255 - 0xff
      13'h1C90: dout  = 8'b00010100; // 7312 :  20 - 0x14 -- Background 0xc9
      13'h1C91: dout  = 8'b00101010; // 7313 :  42 - 0x2a
      13'h1C92: dout  = 8'b00010110; // 7314 :  22 - 0x16
      13'h1C93: dout  = 8'b00101011; // 7315 :  43 - 0x2b
      13'h1C94: dout  = 8'b00010101; // 7316 :  21 - 0x15
      13'h1C95: dout  = 8'b00101011; // 7317 :  43 - 0x2b
      13'h1C96: dout  = 8'b00010101; // 7318 :  21 - 0x15
      13'h1C97: dout  = 8'b00101011; // 7319 :  43 - 0x2b
      13'h1C98: dout  = 8'b11101000; // 7320 : 232 - 0xe8
      13'h1C99: dout  = 8'b11010100; // 7321 : 212 - 0xd4
      13'h1C9A: dout  = 8'b11101000; // 7322 : 232 - 0xe8
      13'h1C9B: dout  = 8'b11010100; // 7323 : 212 - 0xd4
      13'h1C9C: dout  = 8'b11101010; // 7324 : 234 - 0xea
      13'h1C9D: dout  = 8'b11010100; // 7325 : 212 - 0xd4
      13'h1C9E: dout  = 8'b11101010; // 7326 : 234 - 0xea
      13'h1C9F: dout  = 8'b11010100; // 7327 : 212 - 0xd4
      13'h1CA0: dout  = 8'b00000000; // 7328 :   0 - 0x0 -- Background 0xca
      13'h1CA1: dout  = 8'b00000100; // 7329 :   4 - 0x4
      13'h1CA2: dout  = 8'b00000100; // 7330 :   4 - 0x4
      13'h1CA3: dout  = 8'b00000101; // 7331 :   5 - 0x5
      13'h1CA4: dout  = 8'b00010101; // 7332 :  21 - 0x15
      13'h1CA5: dout  = 8'b00010101; // 7333 :  21 - 0x15
      13'h1CA6: dout  = 8'b01010101; // 7334 :  85 - 0x55
      13'h1CA7: dout  = 8'b01010101; // 7335 :  85 - 0x55
      13'h1CA8: dout  = 8'b00000000; // 7336 :   0 - 0x0
      13'h1CA9: dout  = 8'b00000000; // 7337 :   0 - 0x0
      13'h1CAA: dout  = 8'b00000000; // 7338 :   0 - 0x0
      13'h1CAB: dout  = 8'b00000000; // 7339 :   0 - 0x0
      13'h1CAC: dout  = 8'b00000000; // 7340 :   0 - 0x0
      13'h1CAD: dout  = 8'b00000000; // 7341 :   0 - 0x0
      13'h1CAE: dout  = 8'b00000000; // 7342 :   0 - 0x0
      13'h1CAF: dout  = 8'b00000000; // 7343 :   0 - 0x0
      13'h1CB0: dout  = 8'b00000000; // 7344 :   0 - 0x0 -- Background 0xcb
      13'h1CB1: dout  = 8'b00000000; // 7345 :   0 - 0x0
      13'h1CB2: dout  = 8'b00010000; // 7346 :  16 - 0x10
      13'h1CB3: dout  = 8'b00010000; // 7347 :  16 - 0x10
      13'h1CB4: dout  = 8'b01010001; // 7348 :  81 - 0x51
      13'h1CB5: dout  = 8'b01010101; // 7349 :  85 - 0x55
      13'h1CB6: dout  = 8'b01010101; // 7350 :  85 - 0x55
      13'h1CB7: dout  = 8'b01010101; // 7351 :  85 - 0x55
      13'h1CB8: dout  = 8'b00000000; // 7352 :   0 - 0x0
      13'h1CB9: dout  = 8'b00000000; // 7353 :   0 - 0x0
      13'h1CBA: dout  = 8'b00000000; // 7354 :   0 - 0x0
      13'h1CBB: dout  = 8'b00000000; // 7355 :   0 - 0x0
      13'h1CBC: dout  = 8'b00000000; // 7356 :   0 - 0x0
      13'h1CBD: dout  = 8'b00000000; // 7357 :   0 - 0x0
      13'h1CBE: dout  = 8'b00000000; // 7358 :   0 - 0x0
      13'h1CBF: dout  = 8'b00000000; // 7359 :   0 - 0x0
      13'h1CC0: dout  = 8'b00000000; // 7360 :   0 - 0x0 -- Background 0xcc
      13'h1CC1: dout  = 8'b00000000; // 7361 :   0 - 0x0
      13'h1CC2: dout  = 8'b00000000; // 7362 :   0 - 0x0
      13'h1CC3: dout  = 8'b00000101; // 7363 :   5 - 0x5
      13'h1CC4: dout  = 8'b00001111; // 7364 :  15 - 0xf
      13'h1CC5: dout  = 8'b00000111; // 7365 :   7 - 0x7
      13'h1CC6: dout  = 8'b00000011; // 7366 :   3 - 0x3
      13'h1CC7: dout  = 8'b00000001; // 7367 :   1 - 0x1
      13'h1CC8: dout  = 8'b00000000; // 7368 :   0 - 0x0
      13'h1CC9: dout  = 8'b00000000; // 7369 :   0 - 0x0
      13'h1CCA: dout  = 8'b00000000; // 7370 :   0 - 0x0
      13'h1CCB: dout  = 8'b00000000; // 7371 :   0 - 0x0
      13'h1CCC: dout  = 8'b00000101; // 7372 :   5 - 0x5
      13'h1CCD: dout  = 8'b00000010; // 7373 :   2 - 0x2
      13'h1CCE: dout  = 8'b00000001; // 7374 :   1 - 0x1
      13'h1CCF: dout  = 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout  = 8'b00000000; // 7376 :   0 - 0x0 -- Background 0xcd
      13'h1CD1: dout  = 8'b00000000; // 7377 :   0 - 0x0
      13'h1CD2: dout  = 8'b10000000; // 7378 : 128 - 0x80
      13'h1CD3: dout  = 8'b11010000; // 7379 : 208 - 0xd0
      13'h1CD4: dout  = 8'b11111000; // 7380 : 248 - 0xf8
      13'h1CD5: dout  = 8'b11110000; // 7381 : 240 - 0xf0
      13'h1CD6: dout  = 8'b11100000; // 7382 : 224 - 0xe0
      13'h1CD7: dout  = 8'b11000000; // 7383 : 192 - 0xc0
      13'h1CD8: dout  = 8'b00000000; // 7384 :   0 - 0x0
      13'h1CD9: dout  = 8'b00000000; // 7385 :   0 - 0x0
      13'h1CDA: dout  = 8'b00000000; // 7386 :   0 - 0x0
      13'h1CDB: dout  = 8'b10000000; // 7387 : 128 - 0x80
      13'h1CDC: dout  = 8'b01010000; // 7388 :  80 - 0x50
      13'h1CDD: dout  = 8'b10100000; // 7389 : 160 - 0xa0
      13'h1CDE: dout  = 8'b01000000; // 7390 :  64 - 0x40
      13'h1CDF: dout  = 8'b10000000; // 7391 : 128 - 0x80
      13'h1CE0: dout  = 8'b00000000; // 7392 :   0 - 0x0 -- Background 0xce
      13'h1CE1: dout  = 8'b00000000; // 7393 :   0 - 0x0
      13'h1CE2: dout  = 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout  = 8'b01111000; // 7395 : 120 - 0x78
      13'h1CE4: dout  = 8'b11001111; // 7396 : 207 - 0xcf
      13'h1CE5: dout  = 8'b10000000; // 7397 : 128 - 0x80
      13'h1CE6: dout  = 8'b11001111; // 7398 : 207 - 0xcf
      13'h1CE7: dout  = 8'b01001000; // 7399 :  72 - 0x48
      13'h1CE8: dout  = 8'b00000000; // 7400 :   0 - 0x0
      13'h1CE9: dout  = 8'b00000000; // 7401 :   0 - 0x0
      13'h1CEA: dout  = 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout  = 8'b00000000; // 7403 :   0 - 0x0
      13'h1CEC: dout  = 8'b00110000; // 7404 :  48 - 0x30
      13'h1CED: dout  = 8'b01111111; // 7405 : 127 - 0x7f
      13'h1CEE: dout  = 8'b00110000; // 7406 :  48 - 0x30
      13'h1CEF: dout  = 8'b00110000; // 7407 :  48 - 0x30
      13'h1CF0: dout  = 8'b00000000; // 7408 :   0 - 0x0 -- Background 0xcf
      13'h1CF1: dout  = 8'b00000000; // 7409 :   0 - 0x0
      13'h1CF2: dout  = 8'b00000000; // 7410 :   0 - 0x0
      13'h1CF3: dout  = 8'b00011110; // 7411 :  30 - 0x1e
      13'h1CF4: dout  = 8'b11110011; // 7412 : 243 - 0xf3
      13'h1CF5: dout  = 8'b00000001; // 7413 :   1 - 0x1
      13'h1CF6: dout  = 8'b11110011; // 7414 : 243 - 0xf3
      13'h1CF7: dout  = 8'b00010010; // 7415 :  18 - 0x12
      13'h1CF8: dout  = 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout  = 8'b00000000; // 7417 :   0 - 0x0
      13'h1CFA: dout  = 8'b00000000; // 7418 :   0 - 0x0
      13'h1CFB: dout  = 8'b00000000; // 7419 :   0 - 0x0
      13'h1CFC: dout  = 8'b00001100; // 7420 :  12 - 0xc
      13'h1CFD: dout  = 8'b11111110; // 7421 : 254 - 0xfe
      13'h1CFE: dout  = 8'b00001100; // 7422 :  12 - 0xc
      13'h1CFF: dout  = 8'b00001100; // 7423 :  12 - 0xc
      13'h1D00: dout  = 8'b00000000; // 7424 :   0 - 0x0 -- Background 0xd0
      13'h1D01: dout  = 8'b00000000; // 7425 :   0 - 0x0
      13'h1D02: dout  = 8'b00000000; // 7426 :   0 - 0x0
      13'h1D03: dout  = 8'b00000000; // 7427 :   0 - 0x0
      13'h1D04: dout  = 8'b00000000; // 7428 :   0 - 0x0
      13'h1D05: dout  = 8'b00000000; // 7429 :   0 - 0x0
      13'h1D06: dout  = 8'b00000000; // 7430 :   0 - 0x0
      13'h1D07: dout  = 8'b00000000; // 7431 :   0 - 0x0
      13'h1D08: dout  = 8'b00000000; // 7432 :   0 - 0x0
      13'h1D09: dout  = 8'b00000000; // 7433 :   0 - 0x0
      13'h1D0A: dout  = 8'b00000000; // 7434 :   0 - 0x0
      13'h1D0B: dout  = 8'b00000000; // 7435 :   0 - 0x0
      13'h1D0C: dout  = 8'b00000000; // 7436 :   0 - 0x0
      13'h1D0D: dout  = 8'b00000000; // 7437 :   0 - 0x0
      13'h1D0E: dout  = 8'b00000000; // 7438 :   0 - 0x0
      13'h1D0F: dout  = 8'b00000000; // 7439 :   0 - 0x0
      13'h1D10: dout  = 8'b00000000; // 7440 :   0 - 0x0 -- Background 0xd1
      13'h1D11: dout  = 8'b00000000; // 7441 :   0 - 0x0
      13'h1D12: dout  = 8'b00000000; // 7442 :   0 - 0x0
      13'h1D13: dout  = 8'b00000000; // 7443 :   0 - 0x0
      13'h1D14: dout  = 8'b00000000; // 7444 :   0 - 0x0
      13'h1D15: dout  = 8'b00000000; // 7445 :   0 - 0x0
      13'h1D16: dout  = 8'b00000000; // 7446 :   0 - 0x0
      13'h1D17: dout  = 8'b00000000; // 7447 :   0 - 0x0
      13'h1D18: dout  = 8'b00000000; // 7448 :   0 - 0x0
      13'h1D19: dout  = 8'b00000000; // 7449 :   0 - 0x0
      13'h1D1A: dout  = 8'b00000000; // 7450 :   0 - 0x0
      13'h1D1B: dout  = 8'b00000000; // 7451 :   0 - 0x0
      13'h1D1C: dout  = 8'b00000000; // 7452 :   0 - 0x0
      13'h1D1D: dout  = 8'b00000000; // 7453 :   0 - 0x0
      13'h1D1E: dout  = 8'b00000000; // 7454 :   0 - 0x0
      13'h1D1F: dout  = 8'b00000000; // 7455 :   0 - 0x0
      13'h1D20: dout  = 8'b00001000; // 7456 :   8 - 0x8 -- Background 0xd2
      13'h1D21: dout  = 8'b00001100; // 7457 :  12 - 0xc
      13'h1D22: dout  = 8'b00001000; // 7458 :   8 - 0x8
      13'h1D23: dout  = 8'b00001000; // 7459 :   8 - 0x8
      13'h1D24: dout  = 8'b00001010; // 7460 :  10 - 0xa
      13'h1D25: dout  = 8'b00001000; // 7461 :   8 - 0x8
      13'h1D26: dout  = 8'b00001000; // 7462 :   8 - 0x8
      13'h1D27: dout  = 8'b00001100; // 7463 :  12 - 0xc
      13'h1D28: dout  = 8'b00000111; // 7464 :   7 - 0x7
      13'h1D29: dout  = 8'b00000111; // 7465 :   7 - 0x7
      13'h1D2A: dout  = 8'b00000111; // 7466 :   7 - 0x7
      13'h1D2B: dout  = 8'b00000111; // 7467 :   7 - 0x7
      13'h1D2C: dout  = 8'b00000111; // 7468 :   7 - 0x7
      13'h1D2D: dout  = 8'b00000111; // 7469 :   7 - 0x7
      13'h1D2E: dout  = 8'b00000111; // 7470 :   7 - 0x7
      13'h1D2F: dout  = 8'b00000111; // 7471 :   7 - 0x7
      13'h1D30: dout  = 8'b00010000; // 7472 :  16 - 0x10 -- Background 0xd3
      13'h1D31: dout  = 8'b00010000; // 7473 :  16 - 0x10
      13'h1D32: dout  = 8'b00110000; // 7474 :  48 - 0x30
      13'h1D33: dout  = 8'b00010000; // 7475 :  16 - 0x10
      13'h1D34: dout  = 8'b01010000; // 7476 :  80 - 0x50
      13'h1D35: dout  = 8'b00010000; // 7477 :  16 - 0x10
      13'h1D36: dout  = 8'b00110000; // 7478 :  48 - 0x30
      13'h1D37: dout  = 8'b00010000; // 7479 :  16 - 0x10
      13'h1D38: dout  = 8'b11100000; // 7480 : 224 - 0xe0
      13'h1D39: dout  = 8'b11100000; // 7481 : 224 - 0xe0
      13'h1D3A: dout  = 8'b11000000; // 7482 : 192 - 0xc0
      13'h1D3B: dout  = 8'b11100000; // 7483 : 224 - 0xe0
      13'h1D3C: dout  = 8'b10100000; // 7484 : 160 - 0xa0
      13'h1D3D: dout  = 8'b11100000; // 7485 : 224 - 0xe0
      13'h1D3E: dout  = 8'b11000000; // 7486 : 192 - 0xc0
      13'h1D3F: dout  = 8'b11100000; // 7487 : 224 - 0xe0
      13'h1D40: dout  = 8'b00000000; // 7488 :   0 - 0x0 -- Background 0xd4
      13'h1D41: dout  = 8'b00000000; // 7489 :   0 - 0x0
      13'h1D42: dout  = 8'b00000000; // 7490 :   0 - 0x0
      13'h1D43: dout  = 8'b00000000; // 7491 :   0 - 0x0
      13'h1D44: dout  = 8'b00000000; // 7492 :   0 - 0x0
      13'h1D45: dout  = 8'b00000000; // 7493 :   0 - 0x0
      13'h1D46: dout  = 8'b00000000; // 7494 :   0 - 0x0
      13'h1D47: dout  = 8'b00000000; // 7495 :   0 - 0x0
      13'h1D48: dout  = 8'b00000000; // 7496 :   0 - 0x0
      13'h1D49: dout  = 8'b00000000; // 7497 :   0 - 0x0
      13'h1D4A: dout  = 8'b00000000; // 7498 :   0 - 0x0
      13'h1D4B: dout  = 8'b00000000; // 7499 :   0 - 0x0
      13'h1D4C: dout  = 8'b00000000; // 7500 :   0 - 0x0
      13'h1D4D: dout  = 8'b00000000; // 7501 :   0 - 0x0
      13'h1D4E: dout  = 8'b00000000; // 7502 :   0 - 0x0
      13'h1D4F: dout  = 8'b00000000; // 7503 :   0 - 0x0
      13'h1D50: dout  = 8'b11111000; // 7504 : 248 - 0xf8 -- Background 0xd5
      13'h1D51: dout  = 8'b00000110; // 7505 :   6 - 0x6
      13'h1D52: dout  = 8'b00000001; // 7506 :   1 - 0x1
      13'h1D53: dout  = 8'b00000000; // 7507 :   0 - 0x0
      13'h1D54: dout  = 8'b00000000; // 7508 :   0 - 0x0
      13'h1D55: dout  = 8'b00000000; // 7509 :   0 - 0x0
      13'h1D56: dout  = 8'b00000000; // 7510 :   0 - 0x0
      13'h1D57: dout  = 8'b00000000; // 7511 :   0 - 0x0
      13'h1D58: dout  = 8'b00000000; // 7512 :   0 - 0x0
      13'h1D59: dout  = 8'b11111000; // 7513 : 248 - 0xf8
      13'h1D5A: dout  = 8'b11111110; // 7514 : 254 - 0xfe
      13'h1D5B: dout  = 8'b11111111; // 7515 : 255 - 0xff
      13'h1D5C: dout  = 8'b11111111; // 7516 : 255 - 0xff
      13'h1D5D: dout  = 8'b11111111; // 7517 : 255 - 0xff
      13'h1D5E: dout  = 8'b11111111; // 7518 : 255 - 0xff
      13'h1D5F: dout  = 8'b11111111; // 7519 : 255 - 0xff
      13'h1D60: dout  = 8'b00000000; // 7520 :   0 - 0x0 -- Background 0xd6
      13'h1D61: dout  = 8'b00000000; // 7521 :   0 - 0x0
      13'h1D62: dout  = 8'b10000000; // 7522 : 128 - 0x80
      13'h1D63: dout  = 8'b01100000; // 7523 :  96 - 0x60
      13'h1D64: dout  = 8'b01010000; // 7524 :  80 - 0x50
      13'h1D65: dout  = 8'b10101000; // 7525 : 168 - 0xa8
      13'h1D66: dout  = 8'b01011000; // 7526 :  88 - 0x58
      13'h1D67: dout  = 8'b00101100; // 7527 :  44 - 0x2c
      13'h1D68: dout  = 8'b00000000; // 7528 :   0 - 0x0
      13'h1D69: dout  = 8'b00000000; // 7529 :   0 - 0x0
      13'h1D6A: dout  = 8'b00000000; // 7530 :   0 - 0x0
      13'h1D6B: dout  = 8'b10000000; // 7531 : 128 - 0x80
      13'h1D6C: dout  = 8'b10100000; // 7532 : 160 - 0xa0
      13'h1D6D: dout  = 8'b01010000; // 7533 :  80 - 0x50
      13'h1D6E: dout  = 8'b10100000; // 7534 : 160 - 0xa0
      13'h1D6F: dout  = 8'b11010000; // 7535 : 208 - 0xd0
      13'h1D70: dout  = 8'b10100000; // 7536 : 160 - 0xa0 -- Background 0xd7
      13'h1D71: dout  = 8'b11000000; // 7537 : 192 - 0xc0
      13'h1D72: dout  = 8'b10000000; // 7538 : 128 - 0x80
      13'h1D73: dout  = 8'b01010000; // 7539 :  80 - 0x50
      13'h1D74: dout  = 8'b01100000; // 7540 :  96 - 0x60
      13'h1D75: dout  = 8'b00111000; // 7541 :  56 - 0x38
      13'h1D76: dout  = 8'b00001000; // 7542 :   8 - 0x8
      13'h1D77: dout  = 8'b00000111; // 7543 :   7 - 0x7
      13'h1D78: dout  = 8'b01111111; // 7544 : 127 - 0x7f
      13'h1D79: dout  = 8'b01111111; // 7545 : 127 - 0x7f
      13'h1D7A: dout  = 8'b01111111; // 7546 : 127 - 0x7f
      13'h1D7B: dout  = 8'b00111111; // 7547 :  63 - 0x3f
      13'h1D7C: dout  = 8'b00111111; // 7548 :  63 - 0x3f
      13'h1D7D: dout  = 8'b00001111; // 7549 :  15 - 0xf
      13'h1D7E: dout  = 8'b00000111; // 7550 :   7 - 0x7
      13'h1D7F: dout  = 8'b00000000; // 7551 :   0 - 0x0
      13'h1D80: dout  = 8'b00000000; // 7552 :   0 - 0x0 -- Background 0xd8
      13'h1D81: dout  = 8'b00000000; // 7553 :   0 - 0x0
      13'h1D82: dout  = 8'b00000000; // 7554 :   0 - 0x0
      13'h1D83: dout  = 8'b00000000; // 7555 :   0 - 0x0
      13'h1D84: dout  = 8'b00000000; // 7556 :   0 - 0x0
      13'h1D85: dout  = 8'b00000000; // 7557 :   0 - 0x0
      13'h1D86: dout  = 8'b00000000; // 7558 :   0 - 0x0
      13'h1D87: dout  = 8'b11111111; // 7559 : 255 - 0xff
      13'h1D88: dout  = 8'b11111111; // 7560 : 255 - 0xff
      13'h1D89: dout  = 8'b11111111; // 7561 : 255 - 0xff
      13'h1D8A: dout  = 8'b11111111; // 7562 : 255 - 0xff
      13'h1D8B: dout  = 8'b11111111; // 7563 : 255 - 0xff
      13'h1D8C: dout  = 8'b11111111; // 7564 : 255 - 0xff
      13'h1D8D: dout  = 8'b11111111; // 7565 : 255 - 0xff
      13'h1D8E: dout  = 8'b11111111; // 7566 : 255 - 0xff
      13'h1D8F: dout  = 8'b00000000; // 7567 :   0 - 0x0
      13'h1D90: dout  = 8'b00010101; // 7568 :  21 - 0x15 -- Background 0xd9
      13'h1D91: dout  = 8'b00101011; // 7569 :  43 - 0x2b
      13'h1D92: dout  = 8'b00010101; // 7570 :  21 - 0x15
      13'h1D93: dout  = 8'b00101010; // 7571 :  42 - 0x2a
      13'h1D94: dout  = 8'b01010110; // 7572 :  86 - 0x56
      13'h1D95: dout  = 8'b10101100; // 7573 : 172 - 0xac
      13'h1D96: dout  = 8'b01010000; // 7574 :  80 - 0x50
      13'h1D97: dout  = 8'b11100000; // 7575 : 224 - 0xe0
      13'h1D98: dout  = 8'b11101010; // 7576 : 234 - 0xea
      13'h1D99: dout  = 8'b11010100; // 7577 : 212 - 0xd4
      13'h1D9A: dout  = 8'b11101010; // 7578 : 234 - 0xea
      13'h1D9B: dout  = 8'b11010100; // 7579 : 212 - 0xd4
      13'h1D9C: dout  = 8'b10101000; // 7580 : 168 - 0xa8
      13'h1D9D: dout  = 8'b01010000; // 7581 :  80 - 0x50
      13'h1D9E: dout  = 8'b10100000; // 7582 : 160 - 0xa0
      13'h1D9F: dout  = 8'b00000000; // 7583 :   0 - 0x0
      13'h1DA0: dout  = 8'b00000001; // 7584 :   1 - 0x1 -- Background 0xda
      13'h1DA1: dout  = 8'b00001101; // 7585 :  13 - 0xd
      13'h1DA2: dout  = 8'b00010011; // 7586 :  19 - 0x13
      13'h1DA3: dout  = 8'b00001101; // 7587 :  13 - 0xd
      13'h1DA4: dout  = 8'b00000001; // 7588 :   1 - 0x1
      13'h1DA5: dout  = 8'b00000001; // 7589 :   1 - 0x1
      13'h1DA6: dout  = 8'b00000001; // 7590 :   1 - 0x1
      13'h1DA7: dout  = 8'b00000001; // 7591 :   1 - 0x1
      13'h1DA8: dout  = 8'b00000000; // 7592 :   0 - 0x0
      13'h1DA9: dout  = 8'b00000000; // 7593 :   0 - 0x0
      13'h1DAA: dout  = 8'b00001100; // 7594 :  12 - 0xc
      13'h1DAB: dout  = 8'b00000000; // 7595 :   0 - 0x0
      13'h1DAC: dout  = 8'b00000000; // 7596 :   0 - 0x0
      13'h1DAD: dout  = 8'b00000000; // 7597 :   0 - 0x0
      13'h1DAE: dout  = 8'b00000000; // 7598 :   0 - 0x0
      13'h1DAF: dout  = 8'b00000000; // 7599 :   0 - 0x0
      13'h1DB0: dout  = 8'b11000000; // 7600 : 192 - 0xc0 -- Background 0xdb
      13'h1DB1: dout  = 8'b01000000; // 7601 :  64 - 0x40
      13'h1DB2: dout  = 8'b01000000; // 7602 :  64 - 0x40
      13'h1DB3: dout  = 8'b01011000; // 7603 :  88 - 0x58
      13'h1DB4: dout  = 8'b01100100; // 7604 : 100 - 0x64
      13'h1DB5: dout  = 8'b01011000; // 7605 :  88 - 0x58
      13'h1DB6: dout  = 8'b01000000; // 7606 :  64 - 0x40
      13'h1DB7: dout  = 8'b01000000; // 7607 :  64 - 0x40
      13'h1DB8: dout  = 8'b00000000; // 7608 :   0 - 0x0
      13'h1DB9: dout  = 8'b10000000; // 7609 : 128 - 0x80
      13'h1DBA: dout  = 8'b10000000; // 7610 : 128 - 0x80
      13'h1DBB: dout  = 8'b10000000; // 7611 : 128 - 0x80
      13'h1DBC: dout  = 8'b10011000; // 7612 : 152 - 0x98
      13'h1DBD: dout  = 8'b10000000; // 7613 : 128 - 0x80
      13'h1DBE: dout  = 8'b10000000; // 7614 : 128 - 0x80
      13'h1DBF: dout  = 8'b10000000; // 7615 : 128 - 0x80
      13'h1DC0: dout  = 8'b00000000; // 7616 :   0 - 0x0 -- Background 0xdc
      13'h1DC1: dout  = 8'b00000000; // 7617 :   0 - 0x0
      13'h1DC2: dout  = 8'b00000000; // 7618 :   0 - 0x0
      13'h1DC3: dout  = 8'b00000110; // 7619 :   6 - 0x6
      13'h1DC4: dout  = 8'b00000111; // 7620 :   7 - 0x7
      13'h1DC5: dout  = 8'b00000111; // 7621 :   7 - 0x7
      13'h1DC6: dout  = 8'b00000111; // 7622 :   7 - 0x7
      13'h1DC7: dout  = 8'b00000011; // 7623 :   3 - 0x3
      13'h1DC8: dout  = 8'b00000000; // 7624 :   0 - 0x0
      13'h1DC9: dout  = 8'b00000000; // 7625 :   0 - 0x0
      13'h1DCA: dout  = 8'b00000000; // 7626 :   0 - 0x0
      13'h1DCB: dout  = 8'b00000000; // 7627 :   0 - 0x0
      13'h1DCC: dout  = 8'b00000010; // 7628 :   2 - 0x2
      13'h1DCD: dout  = 8'b00000011; // 7629 :   3 - 0x3
      13'h1DCE: dout  = 8'b00000011; // 7630 :   3 - 0x3
      13'h1DCF: dout  = 8'b00000001; // 7631 :   1 - 0x1
      13'h1DD0: dout  = 8'b00000000; // 7632 :   0 - 0x0 -- Background 0xdd
      13'h1DD1: dout  = 8'b00000000; // 7633 :   0 - 0x0
      13'h1DD2: dout  = 8'b00000000; // 7634 :   0 - 0x0
      13'h1DD3: dout  = 8'b10110000; // 7635 : 176 - 0xb0
      13'h1DD4: dout  = 8'b11110000; // 7636 : 240 - 0xf0
      13'h1DD5: dout  = 8'b11110000; // 7637 : 240 - 0xf0
      13'h1DD6: dout  = 8'b11110000; // 7638 : 240 - 0xf0
      13'h1DD7: dout  = 8'b11100000; // 7639 : 224 - 0xe0
      13'h1DD8: dout  = 8'b00000000; // 7640 :   0 - 0x0
      13'h1DD9: dout  = 8'b00000000; // 7641 :   0 - 0x0
      13'h1DDA: dout  = 8'b00000000; // 7642 :   0 - 0x0
      13'h1DDB: dout  = 8'b00000000; // 7643 :   0 - 0x0
      13'h1DDC: dout  = 8'b10100000; // 7644 : 160 - 0xa0
      13'h1DDD: dout  = 8'b11100000; // 7645 : 224 - 0xe0
      13'h1DDE: dout  = 8'b11100000; // 7646 : 224 - 0xe0
      13'h1DDF: dout  = 8'b11000000; // 7647 : 192 - 0xc0
      13'h1DE0: dout  = 8'b11001111; // 7648 : 207 - 0xcf -- Background 0xde
      13'h1DE1: dout  = 8'b10000000; // 7649 : 128 - 0x80
      13'h1DE2: dout  = 8'b11001111; // 7650 : 207 - 0xcf
      13'h1DE3: dout  = 8'b01001000; // 7651 :  72 - 0x48
      13'h1DE4: dout  = 8'b01001000; // 7652 :  72 - 0x48
      13'h1DE5: dout  = 8'b01001000; // 7653 :  72 - 0x48
      13'h1DE6: dout  = 8'b01001000; // 7654 :  72 - 0x48
      13'h1DE7: dout  = 8'b01001000; // 7655 :  72 - 0x48
      13'h1DE8: dout  = 8'b00110000; // 7656 :  48 - 0x30
      13'h1DE9: dout  = 8'b01111111; // 7657 : 127 - 0x7f
      13'h1DEA: dout  = 8'b00110000; // 7658 :  48 - 0x30
      13'h1DEB: dout  = 8'b00110000; // 7659 :  48 - 0x30
      13'h1DEC: dout  = 8'b00110000; // 7660 :  48 - 0x30
      13'h1DED: dout  = 8'b00110000; // 7661 :  48 - 0x30
      13'h1DEE: dout  = 8'b00110000; // 7662 :  48 - 0x30
      13'h1DEF: dout  = 8'b00110000; // 7663 :  48 - 0x30
      13'h1DF0: dout  = 8'b11110011; // 7664 : 243 - 0xf3 -- Background 0xdf
      13'h1DF1: dout  = 8'b00000001; // 7665 :   1 - 0x1
      13'h1DF2: dout  = 8'b11110011; // 7666 : 243 - 0xf3
      13'h1DF3: dout  = 8'b00010010; // 7667 :  18 - 0x12
      13'h1DF4: dout  = 8'b00010010; // 7668 :  18 - 0x12
      13'h1DF5: dout  = 8'b00010010; // 7669 :  18 - 0x12
      13'h1DF6: dout  = 8'b00010010; // 7670 :  18 - 0x12
      13'h1DF7: dout  = 8'b00010010; // 7671 :  18 - 0x12
      13'h1DF8: dout  = 8'b00001100; // 7672 :  12 - 0xc
      13'h1DF9: dout  = 8'b11111110; // 7673 : 254 - 0xfe
      13'h1DFA: dout  = 8'b00001100; // 7674 :  12 - 0xc
      13'h1DFB: dout  = 8'b00001100; // 7675 :  12 - 0xc
      13'h1DFC: dout  = 8'b00001100; // 7676 :  12 - 0xc
      13'h1DFD: dout  = 8'b00001100; // 7677 :  12 - 0xc
      13'h1DFE: dout  = 8'b00001100; // 7678 :  12 - 0xc
      13'h1DFF: dout  = 8'b00001100; // 7679 :  12 - 0xc
      13'h1E00: dout  = 8'b00000000; // 7680 :   0 - 0x0 -- Background 0xe0
      13'h1E01: dout  = 8'b00000000; // 7681 :   0 - 0x0
      13'h1E02: dout  = 8'b00000000; // 7682 :   0 - 0x0
      13'h1E03: dout  = 8'b00000000; // 7683 :   0 - 0x0
      13'h1E04: dout  = 8'b00000000; // 7684 :   0 - 0x0
      13'h1E05: dout  = 8'b00000000; // 7685 :   0 - 0x0
      13'h1E06: dout  = 8'b00000000; // 7686 :   0 - 0x0
      13'h1E07: dout  = 8'b00000000; // 7687 :   0 - 0x0
      13'h1E08: dout  = 8'b00000000; // 7688 :   0 - 0x0
      13'h1E09: dout  = 8'b00000000; // 7689 :   0 - 0x0
      13'h1E0A: dout  = 8'b00000000; // 7690 :   0 - 0x0
      13'h1E0B: dout  = 8'b00000000; // 7691 :   0 - 0x0
      13'h1E0C: dout  = 8'b00000000; // 7692 :   0 - 0x0
      13'h1E0D: dout  = 8'b00000000; // 7693 :   0 - 0x0
      13'h1E0E: dout  = 8'b00000000; // 7694 :   0 - 0x0
      13'h1E0F: dout  = 8'b00000000; // 7695 :   0 - 0x0
      13'h1E10: dout  = 8'b00000000; // 7696 :   0 - 0x0 -- Background 0xe1
      13'h1E11: dout  = 8'b00000000; // 7697 :   0 - 0x0
      13'h1E12: dout  = 8'b00000000; // 7698 :   0 - 0x0
      13'h1E13: dout  = 8'b00000000; // 7699 :   0 - 0x0
      13'h1E14: dout  = 8'b00000000; // 7700 :   0 - 0x0
      13'h1E15: dout  = 8'b00000000; // 7701 :   0 - 0x0
      13'h1E16: dout  = 8'b00000000; // 7702 :   0 - 0x0
      13'h1E17: dout  = 8'b00000000; // 7703 :   0 - 0x0
      13'h1E18: dout  = 8'b00000000; // 7704 :   0 - 0x0
      13'h1E19: dout  = 8'b00000000; // 7705 :   0 - 0x0
      13'h1E1A: dout  = 8'b00000000; // 7706 :   0 - 0x0
      13'h1E1B: dout  = 8'b00000000; // 7707 :   0 - 0x0
      13'h1E1C: dout  = 8'b00000000; // 7708 :   0 - 0x0
      13'h1E1D: dout  = 8'b00000000; // 7709 :   0 - 0x0
      13'h1E1E: dout  = 8'b00000000; // 7710 :   0 - 0x0
      13'h1E1F: dout  = 8'b00000000; // 7711 :   0 - 0x0
      13'h1E20: dout  = 8'b00000000; // 7712 :   0 - 0x0 -- Background 0xe2
      13'h1E21: dout  = 8'b00000000; // 7713 :   0 - 0x0
      13'h1E22: dout  = 8'b00000000; // 7714 :   0 - 0x0
      13'h1E23: dout  = 8'b00000000; // 7715 :   0 - 0x0
      13'h1E24: dout  = 8'b00000000; // 7716 :   0 - 0x0
      13'h1E25: dout  = 8'b00000000; // 7717 :   0 - 0x0
      13'h1E26: dout  = 8'b00000000; // 7718 :   0 - 0x0
      13'h1E27: dout  = 8'b00000000; // 7719 :   0 - 0x0
      13'h1E28: dout  = 8'b00000000; // 7720 :   0 - 0x0
      13'h1E29: dout  = 8'b00000000; // 7721 :   0 - 0x0
      13'h1E2A: dout  = 8'b00000000; // 7722 :   0 - 0x0
      13'h1E2B: dout  = 8'b00000000; // 7723 :   0 - 0x0
      13'h1E2C: dout  = 8'b00000000; // 7724 :   0 - 0x0
      13'h1E2D: dout  = 8'b00000000; // 7725 :   0 - 0x0
      13'h1E2E: dout  = 8'b00000000; // 7726 :   0 - 0x0
      13'h1E2F: dout  = 8'b00000000; // 7727 :   0 - 0x0
      13'h1E30: dout  = 8'b00000000; // 7728 :   0 - 0x0 -- Background 0xe3
      13'h1E31: dout  = 8'b00000000; // 7729 :   0 - 0x0
      13'h1E32: dout  = 8'b00000000; // 7730 :   0 - 0x0
      13'h1E33: dout  = 8'b00000000; // 7731 :   0 - 0x0
      13'h1E34: dout  = 8'b00000000; // 7732 :   0 - 0x0
      13'h1E35: dout  = 8'b00000000; // 7733 :   0 - 0x0
      13'h1E36: dout  = 8'b00000000; // 7734 :   0 - 0x0
      13'h1E37: dout  = 8'b00000000; // 7735 :   0 - 0x0
      13'h1E38: dout  = 8'b00000000; // 7736 :   0 - 0x0
      13'h1E39: dout  = 8'b00000000; // 7737 :   0 - 0x0
      13'h1E3A: dout  = 8'b00000000; // 7738 :   0 - 0x0
      13'h1E3B: dout  = 8'b00000000; // 7739 :   0 - 0x0
      13'h1E3C: dout  = 8'b00000000; // 7740 :   0 - 0x0
      13'h1E3D: dout  = 8'b00000000; // 7741 :   0 - 0x0
      13'h1E3E: dout  = 8'b00000000; // 7742 :   0 - 0x0
      13'h1E3F: dout  = 8'b00000000; // 7743 :   0 - 0x0
      13'h1E40: dout  = 8'b00000000; // 7744 :   0 - 0x0 -- Background 0xe4
      13'h1E41: dout  = 8'b00000000; // 7745 :   0 - 0x0
      13'h1E42: dout  = 8'b00000000; // 7746 :   0 - 0x0
      13'h1E43: dout  = 8'b00000000; // 7747 :   0 - 0x0
      13'h1E44: dout  = 8'b00000000; // 7748 :   0 - 0x0
      13'h1E45: dout  = 8'b00000000; // 7749 :   0 - 0x0
      13'h1E46: dout  = 8'b00000000; // 7750 :   0 - 0x0
      13'h1E47: dout  = 8'b00000000; // 7751 :   0 - 0x0
      13'h1E48: dout  = 8'b00000000; // 7752 :   0 - 0x0
      13'h1E49: dout  = 8'b00000000; // 7753 :   0 - 0x0
      13'h1E4A: dout  = 8'b00000000; // 7754 :   0 - 0x0
      13'h1E4B: dout  = 8'b00000000; // 7755 :   0 - 0x0
      13'h1E4C: dout  = 8'b00000000; // 7756 :   0 - 0x0
      13'h1E4D: dout  = 8'b00000000; // 7757 :   0 - 0x0
      13'h1E4E: dout  = 8'b00000000; // 7758 :   0 - 0x0
      13'h1E4F: dout  = 8'b00000000; // 7759 :   0 - 0x0
      13'h1E50: dout  = 8'b00000000; // 7760 :   0 - 0x0 -- Background 0xe5
      13'h1E51: dout  = 8'b00000000; // 7761 :   0 - 0x0
      13'h1E52: dout  = 8'b00000000; // 7762 :   0 - 0x0
      13'h1E53: dout  = 8'b00000000; // 7763 :   0 - 0x0
      13'h1E54: dout  = 8'b00000000; // 7764 :   0 - 0x0
      13'h1E55: dout  = 8'b00000000; // 7765 :   0 - 0x0
      13'h1E56: dout  = 8'b00000000; // 7766 :   0 - 0x0
      13'h1E57: dout  = 8'b00000000; // 7767 :   0 - 0x0
      13'h1E58: dout  = 8'b00000000; // 7768 :   0 - 0x0
      13'h1E59: dout  = 8'b00000000; // 7769 :   0 - 0x0
      13'h1E5A: dout  = 8'b00000000; // 7770 :   0 - 0x0
      13'h1E5B: dout  = 8'b00000000; // 7771 :   0 - 0x0
      13'h1E5C: dout  = 8'b00000000; // 7772 :   0 - 0x0
      13'h1E5D: dout  = 8'b00000000; // 7773 :   0 - 0x0
      13'h1E5E: dout  = 8'b00000000; // 7774 :   0 - 0x0
      13'h1E5F: dout  = 8'b00000000; // 7775 :   0 - 0x0
      13'h1E60: dout  = 8'b00000000; // 7776 :   0 - 0x0 -- Background 0xe6
      13'h1E61: dout  = 8'b00000000; // 7777 :   0 - 0x0
      13'h1E62: dout  = 8'b00000000; // 7778 :   0 - 0x0
      13'h1E63: dout  = 8'b00000000; // 7779 :   0 - 0x0
      13'h1E64: dout  = 8'b00000000; // 7780 :   0 - 0x0
      13'h1E65: dout  = 8'b00000000; // 7781 :   0 - 0x0
      13'h1E66: dout  = 8'b00000000; // 7782 :   0 - 0x0
      13'h1E67: dout  = 8'b00000000; // 7783 :   0 - 0x0
      13'h1E68: dout  = 8'b00000000; // 7784 :   0 - 0x0
      13'h1E69: dout  = 8'b00000000; // 7785 :   0 - 0x0
      13'h1E6A: dout  = 8'b00000000; // 7786 :   0 - 0x0
      13'h1E6B: dout  = 8'b00000000; // 7787 :   0 - 0x0
      13'h1E6C: dout  = 8'b00000000; // 7788 :   0 - 0x0
      13'h1E6D: dout  = 8'b00000000; // 7789 :   0 - 0x0
      13'h1E6E: dout  = 8'b00000000; // 7790 :   0 - 0x0
      13'h1E6F: dout  = 8'b00000000; // 7791 :   0 - 0x0
      13'h1E70: dout  = 8'b00000000; // 7792 :   0 - 0x0 -- Background 0xe7
      13'h1E71: dout  = 8'b00000000; // 7793 :   0 - 0x0
      13'h1E72: dout  = 8'b00000000; // 7794 :   0 - 0x0
      13'h1E73: dout  = 8'b00000000; // 7795 :   0 - 0x0
      13'h1E74: dout  = 8'b00000000; // 7796 :   0 - 0x0
      13'h1E75: dout  = 8'b00000000; // 7797 :   0 - 0x0
      13'h1E76: dout  = 8'b00000000; // 7798 :   0 - 0x0
      13'h1E77: dout  = 8'b00000000; // 7799 :   0 - 0x0
      13'h1E78: dout  = 8'b00000000; // 7800 :   0 - 0x0
      13'h1E79: dout  = 8'b00000000; // 7801 :   0 - 0x0
      13'h1E7A: dout  = 8'b00000000; // 7802 :   0 - 0x0
      13'h1E7B: dout  = 8'b00000000; // 7803 :   0 - 0x0
      13'h1E7C: dout  = 8'b00000000; // 7804 :   0 - 0x0
      13'h1E7D: dout  = 8'b00000000; // 7805 :   0 - 0x0
      13'h1E7E: dout  = 8'b00000000; // 7806 :   0 - 0x0
      13'h1E7F: dout  = 8'b00000000; // 7807 :   0 - 0x0
      13'h1E80: dout  = 8'b00000000; // 7808 :   0 - 0x0 -- Background 0xe8
      13'h1E81: dout  = 8'b00000000; // 7809 :   0 - 0x0
      13'h1E82: dout  = 8'b00000000; // 7810 :   0 - 0x0
      13'h1E83: dout  = 8'b00000000; // 7811 :   0 - 0x0
      13'h1E84: dout  = 8'b00000000; // 7812 :   0 - 0x0
      13'h1E85: dout  = 8'b00000000; // 7813 :   0 - 0x0
      13'h1E86: dout  = 8'b00000000; // 7814 :   0 - 0x0
      13'h1E87: dout  = 8'b00000000; // 7815 :   0 - 0x0
      13'h1E88: dout  = 8'b00000000; // 7816 :   0 - 0x0
      13'h1E89: dout  = 8'b00000000; // 7817 :   0 - 0x0
      13'h1E8A: dout  = 8'b00000000; // 7818 :   0 - 0x0
      13'h1E8B: dout  = 8'b00000000; // 7819 :   0 - 0x0
      13'h1E8C: dout  = 8'b00000000; // 7820 :   0 - 0x0
      13'h1E8D: dout  = 8'b00000000; // 7821 :   0 - 0x0
      13'h1E8E: dout  = 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout  = 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout  = 8'b00000000; // 7824 :   0 - 0x0 -- Background 0xe9
      13'h1E91: dout  = 8'b00000000; // 7825 :   0 - 0x0
      13'h1E92: dout  = 8'b00000000; // 7826 :   0 - 0x0
      13'h1E93: dout  = 8'b00000000; // 7827 :   0 - 0x0
      13'h1E94: dout  = 8'b00000000; // 7828 :   0 - 0x0
      13'h1E95: dout  = 8'b00000000; // 7829 :   0 - 0x0
      13'h1E96: dout  = 8'b00000000; // 7830 :   0 - 0x0
      13'h1E97: dout  = 8'b00000000; // 7831 :   0 - 0x0
      13'h1E98: dout  = 8'b00000000; // 7832 :   0 - 0x0
      13'h1E99: dout  = 8'b00000000; // 7833 :   0 - 0x0
      13'h1E9A: dout  = 8'b00000000; // 7834 :   0 - 0x0
      13'h1E9B: dout  = 8'b00000000; // 7835 :   0 - 0x0
      13'h1E9C: dout  = 8'b00000000; // 7836 :   0 - 0x0
      13'h1E9D: dout  = 8'b00000000; // 7837 :   0 - 0x0
      13'h1E9E: dout  = 8'b00000000; // 7838 :   0 - 0x0
      13'h1E9F: dout  = 8'b00000000; // 7839 :   0 - 0x0
      13'h1EA0: dout  = 8'b00000000; // 7840 :   0 - 0x0 -- Background 0xea
      13'h1EA1: dout  = 8'b00000000; // 7841 :   0 - 0x0
      13'h1EA2: dout  = 8'b00000000; // 7842 :   0 - 0x0
      13'h1EA3: dout  = 8'b00000000; // 7843 :   0 - 0x0
      13'h1EA4: dout  = 8'b00000000; // 7844 :   0 - 0x0
      13'h1EA5: dout  = 8'b00000000; // 7845 :   0 - 0x0
      13'h1EA6: dout  = 8'b00000000; // 7846 :   0 - 0x0
      13'h1EA7: dout  = 8'b00000000; // 7847 :   0 - 0x0
      13'h1EA8: dout  = 8'b00000000; // 7848 :   0 - 0x0
      13'h1EA9: dout  = 8'b00000000; // 7849 :   0 - 0x0
      13'h1EAA: dout  = 8'b00000000; // 7850 :   0 - 0x0
      13'h1EAB: dout  = 8'b00000000; // 7851 :   0 - 0x0
      13'h1EAC: dout  = 8'b00000000; // 7852 :   0 - 0x0
      13'h1EAD: dout  = 8'b00000000; // 7853 :   0 - 0x0
      13'h1EAE: dout  = 8'b00000000; // 7854 :   0 - 0x0
      13'h1EAF: dout  = 8'b00000000; // 7855 :   0 - 0x0
      13'h1EB0: dout  = 8'b00000000; // 7856 :   0 - 0x0 -- Background 0xeb
      13'h1EB1: dout  = 8'b00000000; // 7857 :   0 - 0x0
      13'h1EB2: dout  = 8'b00000000; // 7858 :   0 - 0x0
      13'h1EB3: dout  = 8'b00000000; // 7859 :   0 - 0x0
      13'h1EB4: dout  = 8'b00000000; // 7860 :   0 - 0x0
      13'h1EB5: dout  = 8'b00000000; // 7861 :   0 - 0x0
      13'h1EB6: dout  = 8'b00000000; // 7862 :   0 - 0x0
      13'h1EB7: dout  = 8'b00000000; // 7863 :   0 - 0x0
      13'h1EB8: dout  = 8'b00000000; // 7864 :   0 - 0x0
      13'h1EB9: dout  = 8'b00000000; // 7865 :   0 - 0x0
      13'h1EBA: dout  = 8'b00000000; // 7866 :   0 - 0x0
      13'h1EBB: dout  = 8'b00000000; // 7867 :   0 - 0x0
      13'h1EBC: dout  = 8'b00000000; // 7868 :   0 - 0x0
      13'h1EBD: dout  = 8'b00000000; // 7869 :   0 - 0x0
      13'h1EBE: dout  = 8'b00000000; // 7870 :   0 - 0x0
      13'h1EBF: dout  = 8'b00000000; // 7871 :   0 - 0x0
      13'h1EC0: dout  = 8'b00000000; // 7872 :   0 - 0x0 -- Background 0xec
      13'h1EC1: dout  = 8'b00000000; // 7873 :   0 - 0x0
      13'h1EC2: dout  = 8'b00000000; // 7874 :   0 - 0x0
      13'h1EC3: dout  = 8'b00000000; // 7875 :   0 - 0x0
      13'h1EC4: dout  = 8'b00000000; // 7876 :   0 - 0x0
      13'h1EC5: dout  = 8'b00000000; // 7877 :   0 - 0x0
      13'h1EC6: dout  = 8'b00000000; // 7878 :   0 - 0x0
      13'h1EC7: dout  = 8'b00000000; // 7879 :   0 - 0x0
      13'h1EC8: dout  = 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout  = 8'b00000000; // 7881 :   0 - 0x0
      13'h1ECA: dout  = 8'b00000000; // 7882 :   0 - 0x0
      13'h1ECB: dout  = 8'b00000000; // 7883 :   0 - 0x0
      13'h1ECC: dout  = 8'b00000000; // 7884 :   0 - 0x0
      13'h1ECD: dout  = 8'b00000000; // 7885 :   0 - 0x0
      13'h1ECE: dout  = 8'b00000000; // 7886 :   0 - 0x0
      13'h1ECF: dout  = 8'b00000000; // 7887 :   0 - 0x0
      13'h1ED0: dout  = 8'b00000000; // 7888 :   0 - 0x0 -- Background 0xed
      13'h1ED1: dout  = 8'b00000000; // 7889 :   0 - 0x0
      13'h1ED2: dout  = 8'b00000000; // 7890 :   0 - 0x0
      13'h1ED3: dout  = 8'b00000000; // 7891 :   0 - 0x0
      13'h1ED4: dout  = 8'b00000000; // 7892 :   0 - 0x0
      13'h1ED5: dout  = 8'b00000000; // 7893 :   0 - 0x0
      13'h1ED6: dout  = 8'b00000000; // 7894 :   0 - 0x0
      13'h1ED7: dout  = 8'b00000000; // 7895 :   0 - 0x0
      13'h1ED8: dout  = 8'b00000000; // 7896 :   0 - 0x0
      13'h1ED9: dout  = 8'b00000000; // 7897 :   0 - 0x0
      13'h1EDA: dout  = 8'b00000000; // 7898 :   0 - 0x0
      13'h1EDB: dout  = 8'b00000000; // 7899 :   0 - 0x0
      13'h1EDC: dout  = 8'b00000000; // 7900 :   0 - 0x0
      13'h1EDD: dout  = 8'b00000000; // 7901 :   0 - 0x0
      13'h1EDE: dout  = 8'b00000000; // 7902 :   0 - 0x0
      13'h1EDF: dout  = 8'b00000000; // 7903 :   0 - 0x0
      13'h1EE0: dout  = 8'b00000000; // 7904 :   0 - 0x0 -- Background 0xee
      13'h1EE1: dout  = 8'b00000000; // 7905 :   0 - 0x0
      13'h1EE2: dout  = 8'b00000000; // 7906 :   0 - 0x0
      13'h1EE3: dout  = 8'b00000000; // 7907 :   0 - 0x0
      13'h1EE4: dout  = 8'b00000000; // 7908 :   0 - 0x0
      13'h1EE5: dout  = 8'b00000000; // 7909 :   0 - 0x0
      13'h1EE6: dout  = 8'b00000000; // 7910 :   0 - 0x0
      13'h1EE7: dout  = 8'b00000000; // 7911 :   0 - 0x0
      13'h1EE8: dout  = 8'b00000000; // 7912 :   0 - 0x0
      13'h1EE9: dout  = 8'b00000000; // 7913 :   0 - 0x0
      13'h1EEA: dout  = 8'b00000000; // 7914 :   0 - 0x0
      13'h1EEB: dout  = 8'b00000000; // 7915 :   0 - 0x0
      13'h1EEC: dout  = 8'b00000000; // 7916 :   0 - 0x0
      13'h1EED: dout  = 8'b00000000; // 7917 :   0 - 0x0
      13'h1EEE: dout  = 8'b00000000; // 7918 :   0 - 0x0
      13'h1EEF: dout  = 8'b00000000; // 7919 :   0 - 0x0
      13'h1EF0: dout  = 8'b00000000; // 7920 :   0 - 0x0 -- Background 0xef
      13'h1EF1: dout  = 8'b00000000; // 7921 :   0 - 0x0
      13'h1EF2: dout  = 8'b00000000; // 7922 :   0 - 0x0
      13'h1EF3: dout  = 8'b00000000; // 7923 :   0 - 0x0
      13'h1EF4: dout  = 8'b00000000; // 7924 :   0 - 0x0
      13'h1EF5: dout  = 8'b00000000; // 7925 :   0 - 0x0
      13'h1EF6: dout  = 8'b00000000; // 7926 :   0 - 0x0
      13'h1EF7: dout  = 8'b00000000; // 7927 :   0 - 0x0
      13'h1EF8: dout  = 8'b00000000; // 7928 :   0 - 0x0
      13'h1EF9: dout  = 8'b00000000; // 7929 :   0 - 0x0
      13'h1EFA: dout  = 8'b00000000; // 7930 :   0 - 0x0
      13'h1EFB: dout  = 8'b00000000; // 7931 :   0 - 0x0
      13'h1EFC: dout  = 8'b00000000; // 7932 :   0 - 0x0
      13'h1EFD: dout  = 8'b00000000; // 7933 :   0 - 0x0
      13'h1EFE: dout  = 8'b00000000; // 7934 :   0 - 0x0
      13'h1EFF: dout  = 8'b00000000; // 7935 :   0 - 0x0
      13'h1F00: dout  = 8'b00000000; // 7936 :   0 - 0x0 -- Background 0xf0
      13'h1F01: dout  = 8'b00000000; // 7937 :   0 - 0x0
      13'h1F02: dout  = 8'b00000000; // 7938 :   0 - 0x0
      13'h1F03: dout  = 8'b00000000; // 7939 :   0 - 0x0
      13'h1F04: dout  = 8'b00000000; // 7940 :   0 - 0x0
      13'h1F05: dout  = 8'b00000000; // 7941 :   0 - 0x0
      13'h1F06: dout  = 8'b00000000; // 7942 :   0 - 0x0
      13'h1F07: dout  = 8'b00000000; // 7943 :   0 - 0x0
      13'h1F08: dout  = 8'b00000000; // 7944 :   0 - 0x0
      13'h1F09: dout  = 8'b00000000; // 7945 :   0 - 0x0
      13'h1F0A: dout  = 8'b00000000; // 7946 :   0 - 0x0
      13'h1F0B: dout  = 8'b00000000; // 7947 :   0 - 0x0
      13'h1F0C: dout  = 8'b00000000; // 7948 :   0 - 0x0
      13'h1F0D: dout  = 8'b00000000; // 7949 :   0 - 0x0
      13'h1F0E: dout  = 8'b00000000; // 7950 :   0 - 0x0
      13'h1F0F: dout  = 8'b00000000; // 7951 :   0 - 0x0
      13'h1F10: dout  = 8'b00000000; // 7952 :   0 - 0x0 -- Background 0xf1
      13'h1F11: dout  = 8'b00000000; // 7953 :   0 - 0x0
      13'h1F12: dout  = 8'b00000000; // 7954 :   0 - 0x0
      13'h1F13: dout  = 8'b00000000; // 7955 :   0 - 0x0
      13'h1F14: dout  = 8'b00000000; // 7956 :   0 - 0x0
      13'h1F15: dout  = 8'b00000000; // 7957 :   0 - 0x0
      13'h1F16: dout  = 8'b00000000; // 7958 :   0 - 0x0
      13'h1F17: dout  = 8'b00000000; // 7959 :   0 - 0x0
      13'h1F18: dout  = 8'b00000000; // 7960 :   0 - 0x0
      13'h1F19: dout  = 8'b00000000; // 7961 :   0 - 0x0
      13'h1F1A: dout  = 8'b00000000; // 7962 :   0 - 0x0
      13'h1F1B: dout  = 8'b00000000; // 7963 :   0 - 0x0
      13'h1F1C: dout  = 8'b00000000; // 7964 :   0 - 0x0
      13'h1F1D: dout  = 8'b00000000; // 7965 :   0 - 0x0
      13'h1F1E: dout  = 8'b00000000; // 7966 :   0 - 0x0
      13'h1F1F: dout  = 8'b00000000; // 7967 :   0 - 0x0
      13'h1F20: dout  = 8'b00000000; // 7968 :   0 - 0x0 -- Background 0xf2
      13'h1F21: dout  = 8'b00000000; // 7969 :   0 - 0x0
      13'h1F22: dout  = 8'b00000000; // 7970 :   0 - 0x0
      13'h1F23: dout  = 8'b00000000; // 7971 :   0 - 0x0
      13'h1F24: dout  = 8'b00000000; // 7972 :   0 - 0x0
      13'h1F25: dout  = 8'b00000000; // 7973 :   0 - 0x0
      13'h1F26: dout  = 8'b00000000; // 7974 :   0 - 0x0
      13'h1F27: dout  = 8'b00000000; // 7975 :   0 - 0x0
      13'h1F28: dout  = 8'b00000000; // 7976 :   0 - 0x0
      13'h1F29: dout  = 8'b00000000; // 7977 :   0 - 0x0
      13'h1F2A: dout  = 8'b00000000; // 7978 :   0 - 0x0
      13'h1F2B: dout  = 8'b00000000; // 7979 :   0 - 0x0
      13'h1F2C: dout  = 8'b00000000; // 7980 :   0 - 0x0
      13'h1F2D: dout  = 8'b00000000; // 7981 :   0 - 0x0
      13'h1F2E: dout  = 8'b00000000; // 7982 :   0 - 0x0
      13'h1F2F: dout  = 8'b00000000; // 7983 :   0 - 0x0
      13'h1F30: dout  = 8'b00000000; // 7984 :   0 - 0x0 -- Background 0xf3
      13'h1F31: dout  = 8'b00000000; // 7985 :   0 - 0x0
      13'h1F32: dout  = 8'b00000000; // 7986 :   0 - 0x0
      13'h1F33: dout  = 8'b00000000; // 7987 :   0 - 0x0
      13'h1F34: dout  = 8'b00000000; // 7988 :   0 - 0x0
      13'h1F35: dout  = 8'b00000000; // 7989 :   0 - 0x0
      13'h1F36: dout  = 8'b00000000; // 7990 :   0 - 0x0
      13'h1F37: dout  = 8'b00000000; // 7991 :   0 - 0x0
      13'h1F38: dout  = 8'b00000000; // 7992 :   0 - 0x0
      13'h1F39: dout  = 8'b00000000; // 7993 :   0 - 0x0
      13'h1F3A: dout  = 8'b00000000; // 7994 :   0 - 0x0
      13'h1F3B: dout  = 8'b00000000; // 7995 :   0 - 0x0
      13'h1F3C: dout  = 8'b00000000; // 7996 :   0 - 0x0
      13'h1F3D: dout  = 8'b00000000; // 7997 :   0 - 0x0
      13'h1F3E: dout  = 8'b00000000; // 7998 :   0 - 0x0
      13'h1F3F: dout  = 8'b00000000; // 7999 :   0 - 0x0
      13'h1F40: dout  = 8'b00000000; // 8000 :   0 - 0x0 -- Background 0xf4
      13'h1F41: dout  = 8'b00000000; // 8001 :   0 - 0x0
      13'h1F42: dout  = 8'b00000000; // 8002 :   0 - 0x0
      13'h1F43: dout  = 8'b00000000; // 8003 :   0 - 0x0
      13'h1F44: dout  = 8'b00000000; // 8004 :   0 - 0x0
      13'h1F45: dout  = 8'b00000000; // 8005 :   0 - 0x0
      13'h1F46: dout  = 8'b00000000; // 8006 :   0 - 0x0
      13'h1F47: dout  = 8'b00000000; // 8007 :   0 - 0x0
      13'h1F48: dout  = 8'b00000000; // 8008 :   0 - 0x0
      13'h1F49: dout  = 8'b00000000; // 8009 :   0 - 0x0
      13'h1F4A: dout  = 8'b00000000; // 8010 :   0 - 0x0
      13'h1F4B: dout  = 8'b00000000; // 8011 :   0 - 0x0
      13'h1F4C: dout  = 8'b00000000; // 8012 :   0 - 0x0
      13'h1F4D: dout  = 8'b00000000; // 8013 :   0 - 0x0
      13'h1F4E: dout  = 8'b00000000; // 8014 :   0 - 0x0
      13'h1F4F: dout  = 8'b00000000; // 8015 :   0 - 0x0
      13'h1F50: dout  = 8'b00000000; // 8016 :   0 - 0x0 -- Background 0xf5
      13'h1F51: dout  = 8'b00000000; // 8017 :   0 - 0x0
      13'h1F52: dout  = 8'b00000000; // 8018 :   0 - 0x0
      13'h1F53: dout  = 8'b00000000; // 8019 :   0 - 0x0
      13'h1F54: dout  = 8'b00000000; // 8020 :   0 - 0x0
      13'h1F55: dout  = 8'b00000000; // 8021 :   0 - 0x0
      13'h1F56: dout  = 8'b00000000; // 8022 :   0 - 0x0
      13'h1F57: dout  = 8'b00000000; // 8023 :   0 - 0x0
      13'h1F58: dout  = 8'b00000000; // 8024 :   0 - 0x0
      13'h1F59: dout  = 8'b00000000; // 8025 :   0 - 0x0
      13'h1F5A: dout  = 8'b00000000; // 8026 :   0 - 0x0
      13'h1F5B: dout  = 8'b00000000; // 8027 :   0 - 0x0
      13'h1F5C: dout  = 8'b00000000; // 8028 :   0 - 0x0
      13'h1F5D: dout  = 8'b00000000; // 8029 :   0 - 0x0
      13'h1F5E: dout  = 8'b00000000; // 8030 :   0 - 0x0
      13'h1F5F: dout  = 8'b00000000; // 8031 :   0 - 0x0
      13'h1F60: dout  = 8'b00000000; // 8032 :   0 - 0x0 -- Background 0xf6
      13'h1F61: dout  = 8'b00000000; // 8033 :   0 - 0x0
      13'h1F62: dout  = 8'b00000000; // 8034 :   0 - 0x0
      13'h1F63: dout  = 8'b00000000; // 8035 :   0 - 0x0
      13'h1F64: dout  = 8'b00000000; // 8036 :   0 - 0x0
      13'h1F65: dout  = 8'b00000000; // 8037 :   0 - 0x0
      13'h1F66: dout  = 8'b00000000; // 8038 :   0 - 0x0
      13'h1F67: dout  = 8'b00000000; // 8039 :   0 - 0x0
      13'h1F68: dout  = 8'b00000000; // 8040 :   0 - 0x0
      13'h1F69: dout  = 8'b00000000; // 8041 :   0 - 0x0
      13'h1F6A: dout  = 8'b00000000; // 8042 :   0 - 0x0
      13'h1F6B: dout  = 8'b00000000; // 8043 :   0 - 0x0
      13'h1F6C: dout  = 8'b00000000; // 8044 :   0 - 0x0
      13'h1F6D: dout  = 8'b00000000; // 8045 :   0 - 0x0
      13'h1F6E: dout  = 8'b00000000; // 8046 :   0 - 0x0
      13'h1F6F: dout  = 8'b00000000; // 8047 :   0 - 0x0
      13'h1F70: dout  = 8'b00000000; // 8048 :   0 - 0x0 -- Background 0xf7
      13'h1F71: dout  = 8'b00000000; // 8049 :   0 - 0x0
      13'h1F72: dout  = 8'b00000000; // 8050 :   0 - 0x0
      13'h1F73: dout  = 8'b00000000; // 8051 :   0 - 0x0
      13'h1F74: dout  = 8'b00000000; // 8052 :   0 - 0x0
      13'h1F75: dout  = 8'b00000000; // 8053 :   0 - 0x0
      13'h1F76: dout  = 8'b00000000; // 8054 :   0 - 0x0
      13'h1F77: dout  = 8'b00000000; // 8055 :   0 - 0x0
      13'h1F78: dout  = 8'b00000000; // 8056 :   0 - 0x0
      13'h1F79: dout  = 8'b00000000; // 8057 :   0 - 0x0
      13'h1F7A: dout  = 8'b00000000; // 8058 :   0 - 0x0
      13'h1F7B: dout  = 8'b00000000; // 8059 :   0 - 0x0
      13'h1F7C: dout  = 8'b00000000; // 8060 :   0 - 0x0
      13'h1F7D: dout  = 8'b00000000; // 8061 :   0 - 0x0
      13'h1F7E: dout  = 8'b00000000; // 8062 :   0 - 0x0
      13'h1F7F: dout  = 8'b00000000; // 8063 :   0 - 0x0
      13'h1F80: dout  = 8'b00000000; // 8064 :   0 - 0x0 -- Background 0xf8
      13'h1F81: dout  = 8'b00000000; // 8065 :   0 - 0x0
      13'h1F82: dout  = 8'b00000000; // 8066 :   0 - 0x0
      13'h1F83: dout  = 8'b00000000; // 8067 :   0 - 0x0
      13'h1F84: dout  = 8'b00000000; // 8068 :   0 - 0x0
      13'h1F85: dout  = 8'b00000000; // 8069 :   0 - 0x0
      13'h1F86: dout  = 8'b00000000; // 8070 :   0 - 0x0
      13'h1F87: dout  = 8'b00000000; // 8071 :   0 - 0x0
      13'h1F88: dout  = 8'b00000000; // 8072 :   0 - 0x0
      13'h1F89: dout  = 8'b00000000; // 8073 :   0 - 0x0
      13'h1F8A: dout  = 8'b00000000; // 8074 :   0 - 0x0
      13'h1F8B: dout  = 8'b00000000; // 8075 :   0 - 0x0
      13'h1F8C: dout  = 8'b00000000; // 8076 :   0 - 0x0
      13'h1F8D: dout  = 8'b00000000; // 8077 :   0 - 0x0
      13'h1F8E: dout  = 8'b00000000; // 8078 :   0 - 0x0
      13'h1F8F: dout  = 8'b00000000; // 8079 :   0 - 0x0
      13'h1F90: dout  = 8'b00000000; // 8080 :   0 - 0x0 -- Background 0xf9
      13'h1F91: dout  = 8'b00000000; // 8081 :   0 - 0x0
      13'h1F92: dout  = 8'b00000000; // 8082 :   0 - 0x0
      13'h1F93: dout  = 8'b00000000; // 8083 :   0 - 0x0
      13'h1F94: dout  = 8'b00000000; // 8084 :   0 - 0x0
      13'h1F95: dout  = 8'b00000000; // 8085 :   0 - 0x0
      13'h1F96: dout  = 8'b00000000; // 8086 :   0 - 0x0
      13'h1F97: dout  = 8'b00000000; // 8087 :   0 - 0x0
      13'h1F98: dout  = 8'b00000000; // 8088 :   0 - 0x0
      13'h1F99: dout  = 8'b00000000; // 8089 :   0 - 0x0
      13'h1F9A: dout  = 8'b00000000; // 8090 :   0 - 0x0
      13'h1F9B: dout  = 8'b00000000; // 8091 :   0 - 0x0
      13'h1F9C: dout  = 8'b00000000; // 8092 :   0 - 0x0
      13'h1F9D: dout  = 8'b00000000; // 8093 :   0 - 0x0
      13'h1F9E: dout  = 8'b00000000; // 8094 :   0 - 0x0
      13'h1F9F: dout  = 8'b00000000; // 8095 :   0 - 0x0
      13'h1FA0: dout  = 8'b00000000; // 8096 :   0 - 0x0 -- Background 0xfa
      13'h1FA1: dout  = 8'b00000000; // 8097 :   0 - 0x0
      13'h1FA2: dout  = 8'b00000000; // 8098 :   0 - 0x0
      13'h1FA3: dout  = 8'b00000000; // 8099 :   0 - 0x0
      13'h1FA4: dout  = 8'b00000000; // 8100 :   0 - 0x0
      13'h1FA5: dout  = 8'b00000000; // 8101 :   0 - 0x0
      13'h1FA6: dout  = 8'b00000000; // 8102 :   0 - 0x0
      13'h1FA7: dout  = 8'b00000000; // 8103 :   0 - 0x0
      13'h1FA8: dout  = 8'b00000000; // 8104 :   0 - 0x0
      13'h1FA9: dout  = 8'b00000000; // 8105 :   0 - 0x0
      13'h1FAA: dout  = 8'b00000000; // 8106 :   0 - 0x0
      13'h1FAB: dout  = 8'b00000000; // 8107 :   0 - 0x0
      13'h1FAC: dout  = 8'b00000000; // 8108 :   0 - 0x0
      13'h1FAD: dout  = 8'b00000000; // 8109 :   0 - 0x0
      13'h1FAE: dout  = 8'b00000000; // 8110 :   0 - 0x0
      13'h1FAF: dout  = 8'b00000000; // 8111 :   0 - 0x0
      13'h1FB0: dout  = 8'b00000000; // 8112 :   0 - 0x0 -- Background 0xfb
      13'h1FB1: dout  = 8'b00000000; // 8113 :   0 - 0x0
      13'h1FB2: dout  = 8'b00000000; // 8114 :   0 - 0x0
      13'h1FB3: dout  = 8'b00000000; // 8115 :   0 - 0x0
      13'h1FB4: dout  = 8'b00000000; // 8116 :   0 - 0x0
      13'h1FB5: dout  = 8'b00000000; // 8117 :   0 - 0x0
      13'h1FB6: dout  = 8'b00000000; // 8118 :   0 - 0x0
      13'h1FB7: dout  = 8'b00000000; // 8119 :   0 - 0x0
      13'h1FB8: dout  = 8'b00000000; // 8120 :   0 - 0x0
      13'h1FB9: dout  = 8'b00000000; // 8121 :   0 - 0x0
      13'h1FBA: dout  = 8'b00000000; // 8122 :   0 - 0x0
      13'h1FBB: dout  = 8'b00000000; // 8123 :   0 - 0x0
      13'h1FBC: dout  = 8'b00000000; // 8124 :   0 - 0x0
      13'h1FBD: dout  = 8'b00000000; // 8125 :   0 - 0x0
      13'h1FBE: dout  = 8'b00000000; // 8126 :   0 - 0x0
      13'h1FBF: dout  = 8'b00000000; // 8127 :   0 - 0x0
      13'h1FC0: dout  = 8'b00000000; // 8128 :   0 - 0x0 -- Background 0xfc
      13'h1FC1: dout  = 8'b00000000; // 8129 :   0 - 0x0
      13'h1FC2: dout  = 8'b10001110; // 8130 : 142 - 0x8e
      13'h1FC3: dout  = 8'b10001010; // 8131 : 138 - 0x8a
      13'h1FC4: dout  = 8'b10001010; // 8132 : 138 - 0x8a
      13'h1FC5: dout  = 8'b10001010; // 8133 : 138 - 0x8a
      13'h1FC6: dout  = 8'b10001010; // 8134 : 138 - 0x8a
      13'h1FC7: dout  = 8'b11101110; // 8135 : 238 - 0xee
      13'h1FC8: dout  = 8'b00000000; // 8136 :   0 - 0x0
      13'h1FC9: dout  = 8'b00000000; // 8137 :   0 - 0x0
      13'h1FCA: dout  = 8'b00000000; // 8138 :   0 - 0x0
      13'h1FCB: dout  = 8'b00000000; // 8139 :   0 - 0x0
      13'h1FCC: dout  = 8'b00000000; // 8140 :   0 - 0x0
      13'h1FCD: dout  = 8'b00000000; // 8141 :   0 - 0x0
      13'h1FCE: dout  = 8'b00000000; // 8142 :   0 - 0x0
      13'h1FCF: dout  = 8'b00000000; // 8143 :   0 - 0x0
      13'h1FD0: dout  = 8'b00000000; // 8144 :   0 - 0x0 -- Background 0xfd
      13'h1FD1: dout  = 8'b00000000; // 8145 :   0 - 0x0
      13'h1FD2: dout  = 8'b01001100; // 8146 :  76 - 0x4c
      13'h1FD3: dout  = 8'b10101010; // 8147 : 170 - 0xaa
      13'h1FD4: dout  = 8'b10101010; // 8148 : 170 - 0xaa
      13'h1FD5: dout  = 8'b11101010; // 8149 : 234 - 0xea
      13'h1FD6: dout  = 8'b10101010; // 8150 : 170 - 0xaa
      13'h1FD7: dout  = 8'b10101100; // 8151 : 172 - 0xac
      13'h1FD8: dout  = 8'b00000000; // 8152 :   0 - 0x0
      13'h1FD9: dout  = 8'b00000000; // 8153 :   0 - 0x0
      13'h1FDA: dout  = 8'b00000000; // 8154 :   0 - 0x0
      13'h1FDB: dout  = 8'b00000000; // 8155 :   0 - 0x0
      13'h1FDC: dout  = 8'b00000000; // 8156 :   0 - 0x0
      13'h1FDD: dout  = 8'b00000000; // 8157 :   0 - 0x0
      13'h1FDE: dout  = 8'b00000000; // 8158 :   0 - 0x0
      13'h1FDF: dout  = 8'b00000000; // 8159 :   0 - 0x0
      13'h1FE0: dout  = 8'b00000000; // 8160 :   0 - 0x0 -- Background 0xfe
      13'h1FE1: dout  = 8'b00000000; // 8161 :   0 - 0x0
      13'h1FE2: dout  = 8'b11101100; // 8162 : 236 - 0xec
      13'h1FE3: dout  = 8'b01001010; // 8163 :  74 - 0x4a
      13'h1FE4: dout  = 8'b01001010; // 8164 :  74 - 0x4a
      13'h1FE5: dout  = 8'b01001010; // 8165 :  74 - 0x4a
      13'h1FE6: dout  = 8'b01001010; // 8166 :  74 - 0x4a
      13'h1FE7: dout  = 8'b11101010; // 8167 : 234 - 0xea
      13'h1FE8: dout  = 8'b00000000; // 8168 :   0 - 0x0
      13'h1FE9: dout  = 8'b00000000; // 8169 :   0 - 0x0
      13'h1FEA: dout  = 8'b00000000; // 8170 :   0 - 0x0
      13'h1FEB: dout  = 8'b00000000; // 8171 :   0 - 0x0
      13'h1FEC: dout  = 8'b00000000; // 8172 :   0 - 0x0
      13'h1FED: dout  = 8'b00000000; // 8173 :   0 - 0x0
      13'h1FEE: dout  = 8'b00000000; // 8174 :   0 - 0x0
      13'h1FEF: dout  = 8'b00000000; // 8175 :   0 - 0x0
      13'h1FF0: dout  = 8'b00000000; // 8176 :   0 - 0x0 -- Background 0xff
      13'h1FF1: dout  = 8'b00000000; // 8177 :   0 - 0x0
      13'h1FF2: dout  = 8'b01100000; // 8178 :  96 - 0x60
      13'h1FF3: dout  = 8'b10001000; // 8179 : 136 - 0x88
      13'h1FF4: dout  = 8'b10100000; // 8180 : 160 - 0xa0
      13'h1FF5: dout  = 8'b10100000; // 8181 : 160 - 0xa0
      13'h1FF6: dout  = 8'b10101000; // 8182 : 168 - 0xa8
      13'h1FF7: dout  = 8'b01000000; // 8183 :  64 - 0x40
      13'h1FF8: dout  = 8'b00000000; // 8184 :   0 - 0x0
      13'h1FF9: dout  = 8'b00000000; // 8185 :   0 - 0x0
      13'h1FFA: dout  = 8'b00000000; // 8186 :   0 - 0x0
      13'h1FFB: dout  = 8'b00000000; // 8187 :   0 - 0x0
      13'h1FFC: dout  = 8'b00000000; // 8188 :   0 - 0x0
      13'h1FFD: dout  = 8'b00000000; // 8189 :   0 - 0x0
      13'h1FFE: dout  = 8'b00000000; // 8190 :   0 - 0x0
      13'h1FFF: dout  = 8'b00000000; // 8191 :   0 - 0x0
    endcase
  end

endmodule
