//- Autcmatically generated verilog ROM from a NES memory file----
//-   SPRITEs MEMORY (OAM)
// https://wiki.nesdev.com/w/index.php/PPU_OAM


//-  Original memory dump file name: smario_traspas_oam.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_OAM_SMARIO_TRASPAS
  (
     //input     clk,   // clock
     input      [8-1:0] addr,  //256 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
      8'h0: dout  = 8'b00011000; //    0 :  24 - 0x18 -- Sprite 0x0
      8'h1: dout  = 8'b11111111; //    1 : 255 - 0xff
      8'h2: dout  = 8'b00100011; //    2 :  35 - 0x23
      8'h3: dout  = 8'b01011000; //    3 :  88 - 0x58
      8'h4: dout  = 8'b10110000; //    4 : 176 - 0xb0 -- Sprite 0x1
      8'h5: dout  = 8'b11111100; //    5 : 252 - 0xfc
      8'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      8'h7: dout  = 8'b01110000; //    7 : 112 - 0x70
      8'h8: dout  = 8'b10110000; //    8 : 176 - 0xb0 -- Sprite 0x2
      8'h9: dout  = 8'b11111100; //    9 : 252 - 0xfc
      8'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      8'hB: dout  = 8'b01111000; //   11 : 120 - 0x78
      8'hC: dout  = 8'b10111000; //   12 : 184 - 0xb8 -- Sprite 0x3
      8'hD: dout  = 8'b11111100; //   13 : 252 - 0xfc
      8'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      8'hF: dout  = 8'b01110000; //   15 : 112 - 0x70
      8'h10: dout  = 8'b10111000; //   16 : 184 - 0xb8 -- Sprite 0x4
      8'h11: dout  = 8'b11111100; //   17 : 252 - 0xfc
      8'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      8'h13: dout  = 8'b01111000; //   19 : 120 - 0x78
      8'h14: dout  = 8'b11000000; //   20 : 192 - 0xc0 -- Sprite 0x5
      8'h15: dout  = 8'b00111010; //   21 :  58 - 0x3a
      8'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      8'h17: dout  = 8'b01110000; //   23 : 112 - 0x70
      8'h18: dout  = 8'b11000000; //   24 : 192 - 0xc0 -- Sprite 0x6
      8'h19: dout  = 8'b00110111; //   25 :  55 - 0x37
      8'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      8'h1B: dout  = 8'b01111000; //   27 : 120 - 0x78
      8'h1C: dout  = 8'b11001000; //   28 : 200 - 0xc8 -- Sprite 0x7
      8'h1D: dout  = 8'b01001111; //   29 :  79 - 0x4f
      8'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      8'h1F: dout  = 8'b01110000; //   31 : 112 - 0x70
      8'h20: dout  = 8'b11001000; //   32 : 200 - 0xc8 -- Sprite 0x8
      8'h21: dout  = 8'b01001111; //   33 :  79 - 0x4f
      8'h22: dout  = 8'b01000000; //   34 :  64 - 0x40
      8'h23: dout  = 8'b01111000; //   35 : 120 - 0x78
      8'h24: dout  = 8'b11111000; //   36 : 248 - 0xf8 -- Sprite 0x9
      8'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      8'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      8'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      8'h28: dout  = 8'b11111000; //   40 : 248 - 0xf8 -- Sprite 0xa
      8'h29: dout  = 8'b11111100; //   41 : 252 - 0xfc
      8'h2A: dout  = 8'b00000001; //   42 :   1 - 0x1
      8'h2B: dout  = 8'b01000010; //   43 :  66 - 0x42
      8'h2C: dout  = 8'b11111000; //   44 : 248 - 0xf8 -- Sprite 0xb
      8'h2D: dout  = 8'b11111100; //   45 : 252 - 0xfc
      8'h2E: dout  = 8'b01000001; //   46 :  65 - 0x41
      8'h2F: dout  = 8'b01001010; //   47 :  74 - 0x4a
      8'h30: dout  = 8'b11111000; //   48 : 248 - 0xf8 -- Sprite 0xc
      8'h31: dout  = 8'b01101111; //   49 : 111 - 0x6f
      8'h32: dout  = 8'b10000001; //   50 : 129 - 0x81
      8'h33: dout  = 8'b01000010; //   51 :  66 - 0x42
      8'h34: dout  = 8'b11111000; //   52 : 248 - 0xf8 -- Sprite 0xd
      8'h35: dout  = 8'b01101111; //   53 : 111 - 0x6f
      8'h36: dout  = 8'b11000001; //   54 : 193 - 0xc1
      8'h37: dout  = 8'b01001010; //   55 :  74 - 0x4a
      8'h38: dout  = 8'b11111000; //   56 : 248 - 0xf8 -- Sprite 0xe
      8'h39: dout  = 8'b01101110; //   57 : 110 - 0x6e
      8'h3A: dout  = 8'b10000001; //   58 : 129 - 0x81
      8'h3B: dout  = 8'b01000010; //   59 :  66 - 0x42
      8'h3C: dout  = 8'b11111000; //   60 : 248 - 0xf8 -- Sprite 0xf
      8'h3D: dout  = 8'b01101110; //   61 : 110 - 0x6e
      8'h3E: dout  = 8'b11000001; //   62 : 193 - 0xc1
      8'h3F: dout  = 8'b01001010; //   63 :  74 - 0x4a
      8'h40: dout  = 8'b11111000; //   64 : 248 - 0xf8 -- Sprite 0x10
      8'h41: dout  = 8'b01110011; //   65 : 115 - 0x73
      8'h42: dout  = 8'b01000011; //   66 :  67 - 0x43
      8'h43: dout  = 8'b10111101; //   67 : 189 - 0xbd
      8'h44: dout  = 8'b11111000; //   68 : 248 - 0xf8 -- Sprite 0x11
      8'h45: dout  = 8'b01110010; //   69 : 114 - 0x72
      8'h46: dout  = 8'b01000011; //   70 :  67 - 0x43
      8'h47: dout  = 8'b11000101; //   71 : 197 - 0xc5
      8'h48: dout  = 8'b11111000; //   72 : 248 - 0xf8 -- Sprite 0x12
      8'h49: dout  = 8'b11110110; //   73 : 246 - 0xf6
      8'h4A: dout  = 8'b00000010; //   74 :   2 - 0x2
      8'h4B: dout  = 8'b01011000; //   75 :  88 - 0x58
      8'h4C: dout  = 8'b11111000; //   76 : 248 - 0xf8 -- Sprite 0x13
      8'h4D: dout  = 8'b11111011; //   77 : 251 - 0xfb
      8'h4E: dout  = 8'b00000010; //   78 :   2 - 0x2
      8'h4F: dout  = 8'b01100000; //   79 :  96 - 0x60
      8'h50: dout  = 8'b11111000; //   80 : 248 - 0xf8 -- Sprite 0x14
      8'h51: dout  = 8'b11111100; //   81 : 252 - 0xfc
      8'h52: dout  = 8'b10000011; //   82 : 131 - 0x83
      8'h53: dout  = 8'b00101111; //   83 :  47 - 0x2f
      8'h54: dout  = 8'b11111000; //   84 : 248 - 0xf8 -- Sprite 0x15
      8'h55: dout  = 8'b11111100; //   85 : 252 - 0xfc
      8'h56: dout  = 8'b11000011; //   86 : 195 - 0xc3
      8'h57: dout  = 8'b00110111; //   87 :  55 - 0x37
      8'h58: dout  = 8'b11111000; //   88 : 248 - 0xf8 -- Sprite 0x16
      8'h59: dout  = 8'b11101111; //   89 : 239 - 0xef
      8'h5A: dout  = 8'b10000011; //   90 : 131 - 0x83
      8'h5B: dout  = 8'b00101111; //   91 :  47 - 0x2f
      8'h5C: dout  = 8'b11111000; //   92 : 248 - 0xf8 -- Sprite 0x17
      8'h5D: dout  = 8'b11101111; //   93 : 239 - 0xef
      8'h5E: dout  = 8'b11000011; //   94 : 195 - 0xc3
      8'h5F: dout  = 8'b00110111; //   95 :  55 - 0x37
      8'h60: dout  = 8'b11111000; //   96 : 248 - 0xf8 -- Sprite 0x18
      8'h61: dout  = 8'b11111100; //   97 : 252 - 0xfc
      8'h62: dout  = 8'b00000001; //   98 :   1 - 0x1
      8'h63: dout  = 8'b01000100; //   99 :  68 - 0x44
      8'h64: dout  = 8'b11111000; //  100 : 248 - 0xf8 -- Sprite 0x19
      8'h65: dout  = 8'b11111100; //  101 : 252 - 0xfc
      8'h66: dout  = 8'b01000001; //  102 :  65 - 0x41
      8'h67: dout  = 8'b01001100; //  103 :  76 - 0x4c
      8'h68: dout  = 8'b11111000; //  104 : 248 - 0xf8 -- Sprite 0x1a
      8'h69: dout  = 8'b01101111; //  105 : 111 - 0x6f
      8'h6A: dout  = 8'b10000001; //  106 : 129 - 0x81
      8'h6B: dout  = 8'b01000100; //  107 :  68 - 0x44
      8'h6C: dout  = 8'b11111000; //  108 : 248 - 0xf8 -- Sprite 0x1b
      8'h6D: dout  = 8'b01101111; //  109 : 111 - 0x6f
      8'h6E: dout  = 8'b11000001; //  110 : 193 - 0xc1
      8'h6F: dout  = 8'b01001100; //  111 :  76 - 0x4c
      8'h70: dout  = 8'b11111000; //  112 : 248 - 0xf8 -- Sprite 0x1c
      8'h71: dout  = 8'b01101110; //  113 : 110 - 0x6e
      8'h72: dout  = 8'b10000001; //  114 : 129 - 0x81
      8'h73: dout  = 8'b01000100; //  115 :  68 - 0x44
      8'h74: dout  = 8'b11111000; //  116 : 248 - 0xf8 -- Sprite 0x1d
      8'h75: dout  = 8'b01101110; //  117 : 110 - 0x6e
      8'h76: dout  = 8'b11000001; //  118 : 193 - 0xc1
      8'h77: dout  = 8'b01001100; //  119 :  76 - 0x4c
      8'h78: dout  = 8'b11111000; //  120 : 248 - 0xf8 -- Sprite 0x1e
      8'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      8'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      8'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      8'h7C: dout  = 8'b11111000; //  124 : 248 - 0xf8 -- Sprite 0x1f
      8'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      8'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      8'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      8'h80: dout  = 8'b11111000; //  128 : 248 - 0xf8 -- Sprite 0x20
      8'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      8'h82: dout  = 8'b00000000; //  130 :   0 - 0x0
      8'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      8'h84: dout  = 8'b11111000; //  132 : 248 - 0xf8 -- Sprite 0x21
      8'h85: dout  = 8'b00000000; //  133 :   0 - 0x0
      8'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      8'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      8'h88: dout  = 8'b11111000; //  136 : 248 - 0xf8 -- Sprite 0x22
      8'h89: dout  = 8'b11111100; //  137 : 252 - 0xfc
      8'h8A: dout  = 8'b01000011; //  138 :  67 - 0x43
      8'h8B: dout  = 8'b10111110; //  139 : 190 - 0xbe
      8'h8C: dout  = 8'b11111000; //  140 : 248 - 0xf8 -- Sprite 0x23
      8'h8D: dout  = 8'b11111100; //  141 : 252 - 0xfc
      8'h8E: dout  = 8'b01000011; //  142 :  67 - 0x43
      8'h8F: dout  = 8'b11000110; //  143 : 198 - 0xc6
      8'h90: dout  = 8'b11111000; //  144 : 248 - 0xf8 -- Sprite 0x24
      8'h91: dout  = 8'b01110001; //  145 : 113 - 0x71
      8'h92: dout  = 8'b01000011; //  146 :  67 - 0x43
      8'h93: dout  = 8'b10111110; //  147 : 190 - 0xbe
      8'h94: dout  = 8'b11111000; //  148 : 248 - 0xf8 -- Sprite 0x25
      8'h95: dout  = 8'b01110000; //  149 : 112 - 0x70
      8'h96: dout  = 8'b01000011; //  150 :  67 - 0x43
      8'h97: dout  = 8'b11000110; //  151 : 198 - 0xc6
      8'h98: dout  = 8'b11111000; //  152 : 248 - 0xf8 -- Sprite 0x26
      8'h99: dout  = 8'b01110011; //  153 : 115 - 0x73
      8'h9A: dout  = 8'b01000011; //  154 :  67 - 0x43
      8'h9B: dout  = 8'b10111110; //  155 : 190 - 0xbe
      8'h9C: dout  = 8'b11111000; //  156 : 248 - 0xf8 -- Sprite 0x27
      8'h9D: dout  = 8'b01110010; //  157 : 114 - 0x72
      8'h9E: dout  = 8'b01000011; //  158 :  67 - 0x43
      8'h9F: dout  = 8'b11000110; //  159 : 198 - 0xc6
      8'hA0: dout  = 8'b11111000; //  160 : 248 - 0xf8 -- Sprite 0x28
      8'hA1: dout  = 8'b11111100; //  161 : 252 - 0xfc
      8'hA2: dout  = 8'b00000011; //  162 :   3 - 0x3
      8'hA3: dout  = 8'b00101110; //  163 :  46 - 0x2e
      8'hA4: dout  = 8'b11111000; //  164 : 248 - 0xf8 -- Sprite 0x29
      8'hA5: dout  = 8'b11111100; //  165 : 252 - 0xfc
      8'hA6: dout  = 8'b01000011; //  166 :  67 - 0x43
      8'hA7: dout  = 8'b00110110; //  167 :  54 - 0x36
      8'hA8: dout  = 8'b11111000; //  168 : 248 - 0xf8 -- Sprite 0x2a
      8'hA9: dout  = 8'b11111100; //  169 : 252 - 0xfc
      8'hAA: dout  = 8'b10000011; //  170 : 131 - 0x83
      8'hAB: dout  = 8'b00101110; //  171 :  46 - 0x2e
      8'hAC: dout  = 8'b11111000; //  172 : 248 - 0xf8 -- Sprite 0x2b
      8'hAD: dout  = 8'b11111100; //  173 : 252 - 0xfc
      8'hAE: dout  = 8'b11000011; //  174 : 195 - 0xc3
      8'hAF: dout  = 8'b00110110; //  175 :  54 - 0x36
      8'hB0: dout  = 8'b11111000; //  176 : 248 - 0xf8 -- Sprite 0x2c
      8'hB1: dout  = 8'b11101111; //  177 : 239 - 0xef
      8'hB2: dout  = 8'b10000011; //  178 : 131 - 0x83
      8'hB3: dout  = 8'b00101110; //  179 :  46 - 0x2e
      8'hB4: dout  = 8'b11111000; //  180 : 248 - 0xf8 -- Sprite 0x2d
      8'hB5: dout  = 8'b11101111; //  181 : 239 - 0xef
      8'hB6: dout  = 8'b11000011; //  182 : 195 - 0xc3
      8'hB7: dout  = 8'b00110110; //  183 :  54 - 0x36
      8'hB8: dout  = 8'b11111000; //  184 : 248 - 0xf8 -- Sprite 0x2e
      8'hB9: dout  = 8'b11111100; //  185 : 252 - 0xfc
      8'hBA: dout  = 8'b00000001; //  186 :   1 - 0x1
      8'hBB: dout  = 8'b01000111; //  187 :  71 - 0x47
      8'hBC: dout  = 8'b11111000; //  188 : 248 - 0xf8 -- Sprite 0x2f
      8'hBD: dout  = 8'b11111100; //  189 : 252 - 0xfc
      8'hBE: dout  = 8'b01000001; //  190 :  65 - 0x41
      8'hBF: dout  = 8'b01001111; //  191 :  79 - 0x4f
      8'hC0: dout  = 8'b11111000; //  192 : 248 - 0xf8 -- Sprite 0x30
      8'hC1: dout  = 8'b01101111; //  193 : 111 - 0x6f
      8'hC2: dout  = 8'b10000001; //  194 : 129 - 0x81
      8'hC3: dout  = 8'b01000111; //  195 :  71 - 0x47
      8'hC4: dout  = 8'b11111000; //  196 : 248 - 0xf8 -- Sprite 0x31
      8'hC5: dout  = 8'b01101111; //  197 : 111 - 0x6f
      8'hC6: dout  = 8'b11000001; //  198 : 193 - 0xc1
      8'hC7: dout  = 8'b01001111; //  199 :  79 - 0x4f
      8'hC8: dout  = 8'b11111000; //  200 : 248 - 0xf8 -- Sprite 0x32
      8'hC9: dout  = 8'b01101110; //  201 : 110 - 0x6e
      8'hCA: dout  = 8'b10000001; //  202 : 129 - 0x81
      8'hCB: dout  = 8'b01000111; //  203 :  71 - 0x47
      8'hCC: dout  = 8'b11111000; //  204 : 248 - 0xf8 -- Sprite 0x33
      8'hCD: dout  = 8'b01101110; //  205 : 110 - 0x6e
      8'hCE: dout  = 8'b11000001; //  206 : 193 - 0xc1
      8'hCF: dout  = 8'b01001111; //  207 :  79 - 0x4f
      8'hD0: dout  = 8'b11111000; //  208 : 248 - 0xf8 -- Sprite 0x34
      8'hD1: dout  = 8'b11111100; //  209 : 252 - 0xfc
      8'hD2: dout  = 8'b01000011; //  210 :  67 - 0x43
      8'hD3: dout  = 8'b10111110; //  211 : 190 - 0xbe
      8'hD4: dout  = 8'b11111000; //  212 : 248 - 0xf8 -- Sprite 0x35
      8'hD5: dout  = 8'b11111100; //  213 : 252 - 0xfc
      8'hD6: dout  = 8'b01000011; //  214 :  67 - 0x43
      8'hD7: dout  = 8'b11000110; //  215 : 198 - 0xc6
      8'hD8: dout  = 8'b11111000; //  216 : 248 - 0xf8 -- Sprite 0x36
      8'hD9: dout  = 8'b01110001; //  217 : 113 - 0x71
      8'hDA: dout  = 8'b01000011; //  218 :  67 - 0x43
      8'hDB: dout  = 8'b10111110; //  219 : 190 - 0xbe
      8'hDC: dout  = 8'b11111000; //  220 : 248 - 0xf8 -- Sprite 0x37
      8'hDD: dout  = 8'b01110000; //  221 : 112 - 0x70
      8'hDE: dout  = 8'b01000011; //  222 :  67 - 0x43
      8'hDF: dout  = 8'b11000110; //  223 : 198 - 0xc6
      8'hE0: dout  = 8'b11111000; //  224 : 248 - 0xf8 -- Sprite 0x38
      8'hE1: dout  = 8'b01110011; //  225 : 115 - 0x73
      8'hE2: dout  = 8'b01000011; //  226 :  67 - 0x43
      8'hE3: dout  = 8'b10111110; //  227 : 190 - 0xbe
      8'hE4: dout  = 8'b11111000; //  228 : 248 - 0xf8 -- Sprite 0x39
      8'hE5: dout  = 8'b01110010; //  229 : 114 - 0x72
      8'hE6: dout  = 8'b01000011; //  230 :  67 - 0x43
      8'hE7: dout  = 8'b11000110; //  231 : 198 - 0xc6
      8'hE8: dout  = 8'b11111000; //  232 : 248 - 0xf8 -- Sprite 0x3a
      8'hE9: dout  = 8'b11110110; //  233 : 246 - 0xf6
      8'hEA: dout  = 8'b00000010; //  234 :   2 - 0x2
      8'hEB: dout  = 8'b01011000; //  235 :  88 - 0x58
      8'hEC: dout  = 8'b11111000; //  236 : 248 - 0xf8 -- Sprite 0x3b
      8'hED: dout  = 8'b11111011; //  237 : 251 - 0xfb
      8'hEE: dout  = 8'b00000010; //  238 :   2 - 0x2
      8'hEF: dout  = 8'b01100000; //  239 :  96 - 0x60
      8'hF0: dout  = 8'b11111000; //  240 : 248 - 0xf8 -- Sprite 0x3c
      8'hF1: dout  = 8'b11111100; //  241 : 252 - 0xfc
      8'hF2: dout  = 8'b10000011; //  242 : 131 - 0x83
      8'hF3: dout  = 8'b00110000; //  243 :  48 - 0x30
      8'hF4: dout  = 8'b11111000; //  244 : 248 - 0xf8 -- Sprite 0x3d
      8'hF5: dout  = 8'b11111100; //  245 : 252 - 0xfc
      8'hF6: dout  = 8'b11000011; //  246 : 195 - 0xc3
      8'hF7: dout  = 8'b00111000; //  247 :  56 - 0x38
      8'hF8: dout  = 8'b11111000; //  248 : 248 - 0xf8 -- Sprite 0x3e
      8'hF9: dout  = 8'b11101111; //  249 : 239 - 0xef
      8'hFA: dout  = 8'b10000011; //  250 : 131 - 0x83
      8'hFB: dout  = 8'b00110000; //  251 :  48 - 0x30
      8'hFC: dout  = 8'b11111000; //  252 : 248 - 0xf8 -- Sprite 0x3f
      8'hFD: dout  = 8'b11101111; //  253 : 239 - 0xef
      8'hFE: dout  = 8'b11000011; //  254 : 195 - 0xc3
      8'hFF: dout  = 8'b00111000; //  255 :  56 - 0x38
    endcase
  end

endmodule
