//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_DONKEYKONG_SPR
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      12'h2: dout <= 8'b00000111; //    2 :   7 - 0x7
      12'h3: dout <= 8'b00000111; //    3 :   7 - 0x7
      12'h4: dout <= 8'b00001001; //    4 :   9 - 0x9
      12'h5: dout <= 8'b00001001; //    5 :   9 - 0x9
      12'h6: dout <= 8'b00011100; //    6 :  28 - 0x1c
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b00000011; //    9 :   3 - 0x3
      12'hA: dout <= 8'b00000111; //   10 :   7 - 0x7
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000110; //   12 :   6 - 0x6
      12'hD: dout <= 8'b00000110; //   13 :   6 - 0x6
      12'hE: dout <= 8'b00000011; //   14 :   3 - 0x3
      12'hF: dout <= 8'b00000011; //   15 :   3 - 0x3
      12'h10: dout <= 8'b00001111; //   16 :  15 - 0xf -- Sprite 0x1
      12'h11: dout <= 8'b00001111; //   17 :  15 - 0xf
      12'h12: dout <= 8'b00001111; //   18 :  15 - 0xf
      12'h13: dout <= 8'b11111111; //   19 : 255 - 0xff
      12'h14: dout <= 8'b11111111; //   20 : 255 - 0xff
      12'h15: dout <= 8'b11111100; //   21 : 252 - 0xfc
      12'h16: dout <= 8'b10000001; //   22 : 129 - 0x81
      12'h17: dout <= 8'b00000001; //   23 :   1 - 0x1
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b00010000; //   25 :  16 - 0x10
      12'h1A: dout <= 8'b00111100; //   26 :  60 - 0x3c
      12'h1B: dout <= 8'b00111111; //   27 :  63 - 0x3f
      12'h1C: dout <= 8'b00111111; //   28 :  63 - 0x3f
      12'h1D: dout <= 8'b00111100; //   29 :  60 - 0x3c
      12'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      12'h21: dout <= 8'b11000000; //   33 : 192 - 0xc0
      12'h22: dout <= 8'b11111000; //   34 : 248 - 0xf8
      12'h23: dout <= 8'b10000000; //   35 : 128 - 0x80
      12'h24: dout <= 8'b00100000; //   36 :  32 - 0x20
      12'h25: dout <= 8'b10010000; //   37 : 144 - 0x90
      12'h26: dout <= 8'b00111100; //   38 :  60 - 0x3c
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b11000000; //   41 : 192 - 0xc0
      12'h2A: dout <= 8'b11111000; //   42 : 248 - 0xf8
      12'h2B: dout <= 8'b01100000; //   43 :  96 - 0x60
      12'h2C: dout <= 8'b11011100; //   44 : 220 - 0xdc
      12'h2D: dout <= 8'b01101110; //   45 : 110 - 0x6e
      12'h2E: dout <= 8'b11000000; //   46 : 192 - 0xc0
      12'h2F: dout <= 8'b11111000; //   47 : 248 - 0xf8
      12'h30: dout <= 8'b11000000; //   48 : 192 - 0xc0 -- Sprite 0x3
      12'h31: dout <= 8'b11000000; //   49 : 192 - 0xc0
      12'h32: dout <= 8'b11000000; //   50 : 192 - 0xc0
      12'h33: dout <= 8'b11110000; //   51 : 240 - 0xf0
      12'h34: dout <= 8'b11110000; //   52 : 240 - 0xf0
      12'h35: dout <= 8'b11100000; //   53 : 224 - 0xe0
      12'h36: dout <= 8'b11000000; //   54 : 192 - 0xc0
      12'h37: dout <= 8'b11100000; //   55 : 224 - 0xe0
      12'h38: dout <= 8'b01010000; //   56 :  80 - 0x50 -- plane 1
      12'h39: dout <= 8'b00111000; //   57 :  56 - 0x38
      12'h3A: dout <= 8'b00110000; //   58 :  48 - 0x30
      12'h3B: dout <= 8'b11110000; //   59 : 240 - 0xf0
      12'h3C: dout <= 8'b11110000; //   60 : 240 - 0xf0
      12'h3D: dout <= 8'b11100000; //   61 : 224 - 0xe0
      12'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b00000111; //   64 :   7 - 0x7 -- Sprite 0x4
      12'h41: dout <= 8'b00001111; //   65 :  15 - 0xf
      12'h42: dout <= 8'b00001111; //   66 :  15 - 0xf
      12'h43: dout <= 8'b00010010; //   67 :  18 - 0x12
      12'h44: dout <= 8'b00010011; //   68 :  19 - 0x13
      12'h45: dout <= 8'b00111000; //   69 :  56 - 0x38
      12'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout <= 8'b00001111; //   71 :  15 - 0xf
      12'h48: dout <= 8'b00000111; //   72 :   7 - 0x7 -- plane 1
      12'h49: dout <= 8'b00001111; //   73 :  15 - 0xf
      12'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout <= 8'b00001101; //   75 :  13 - 0xd
      12'h4C: dout <= 8'b00001100; //   76 :  12 - 0xc
      12'h4D: dout <= 8'b00000111; //   77 :   7 - 0x7
      12'h4E: dout <= 8'b00000111; //   78 :   7 - 0x7
      12'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout <= 8'b00011111; //   80 :  31 - 0x1f -- Sprite 0x5
      12'h51: dout <= 8'b00011111; //   81 :  31 - 0x1f
      12'h52: dout <= 8'b00011111; //   82 :  31 - 0x1f
      12'h53: dout <= 8'b00011000; //   83 :  24 - 0x18
      12'h54: dout <= 8'b00011001; //   84 :  25 - 0x19
      12'h55: dout <= 8'b00011110; //   85 :  30 - 0x1e
      12'h56: dout <= 8'b00011100; //   86 :  28 - 0x1c
      12'h57: dout <= 8'b00011110; //   87 :  30 - 0x1e
      12'h58: dout <= 8'b00000001; //   88 :   1 - 0x1 -- plane 1
      12'h59: dout <= 8'b00000011; //   89 :   3 - 0x3
      12'h5A: dout <= 8'b00000001; //   90 :   1 - 0x1
      12'h5B: dout <= 8'b00010111; //   91 :  23 - 0x17
      12'h5C: dout <= 8'b00011111; //   92 :  31 - 0x1f
      12'h5D: dout <= 8'b00011110; //   93 :  30 - 0x1e
      12'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b10000000; //   96 : 128 - 0x80 -- Sprite 0x6
      12'h61: dout <= 8'b11110000; //   97 : 240 - 0xf0
      12'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      12'h63: dout <= 8'b01000000; //   99 :  64 - 0x40
      12'h64: dout <= 8'b00100000; //  100 :  32 - 0x20
      12'h65: dout <= 8'b01111000; //  101 : 120 - 0x78
      12'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout <= 8'b11000000; //  103 : 192 - 0xc0
      12'h68: dout <= 8'b10000000; //  104 : 128 - 0x80 -- plane 1
      12'h69: dout <= 8'b11110000; //  105 : 240 - 0xf0
      12'h6A: dout <= 8'b11000000; //  106 : 192 - 0xc0
      12'h6B: dout <= 8'b10111000; //  107 : 184 - 0xb8
      12'h6C: dout <= 8'b11011100; //  108 : 220 - 0xdc
      12'h6D: dout <= 8'b10000000; //  109 : 128 - 0x80
      12'h6E: dout <= 8'b11110000; //  110 : 240 - 0xf0
      12'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout <= 8'b11100000; //  112 : 224 - 0xe0 -- Sprite 0x7
      12'h71: dout <= 8'b01100000; //  113 :  96 - 0x60
      12'h72: dout <= 8'b11110000; //  114 : 240 - 0xf0
      12'h73: dout <= 8'b11110000; //  115 : 240 - 0xf0
      12'h74: dout <= 8'b11110000; //  116 : 240 - 0xf0
      12'h75: dout <= 8'b11100000; //  117 : 224 - 0xe0
      12'h76: dout <= 8'b11100000; //  118 : 224 - 0xe0
      12'h77: dout <= 8'b11110000; //  119 : 240 - 0xf0
      12'h78: dout <= 8'b10000000; //  120 : 128 - 0x80 -- plane 1
      12'h79: dout <= 8'b11100000; //  121 : 224 - 0xe0
      12'h7A: dout <= 8'b11110000; //  122 : 240 - 0xf0
      12'h7B: dout <= 8'b11110000; //  123 : 240 - 0xf0
      12'h7C: dout <= 8'b11110000; //  124 : 240 - 0xf0
      12'h7D: dout <= 8'b11100000; //  125 : 224 - 0xe0
      12'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b00000111; //  128 :   7 - 0x7 -- Sprite 0x8
      12'h81: dout <= 8'b00001111; //  129 :  15 - 0xf
      12'h82: dout <= 8'b00001111; //  130 :  15 - 0xf
      12'h83: dout <= 8'b00010010; //  131 :  18 - 0x12
      12'h84: dout <= 8'b00010011; //  132 :  19 - 0x13
      12'h85: dout <= 8'b00111000; //  133 :  56 - 0x38
      12'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout <= 8'b00111111; //  135 :  63 - 0x3f
      12'h88: dout <= 8'b00000111; //  136 :   7 - 0x7 -- plane 1
      12'h89: dout <= 8'b00001111; //  137 :  15 - 0xf
      12'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout <= 8'b00001101; //  139 :  13 - 0xd
      12'h8C: dout <= 8'b00001100; //  140 :  12 - 0xc
      12'h8D: dout <= 8'b00000111; //  141 :   7 - 0x7
      12'h8E: dout <= 8'b00000111; //  142 :   7 - 0x7
      12'h8F: dout <= 8'b00000011; //  143 :   3 - 0x3
      12'h90: dout <= 8'b00111111; //  144 :  63 - 0x3f -- Sprite 0x9
      12'h91: dout <= 8'b00001110; //  145 :  14 - 0xe
      12'h92: dout <= 8'b00001111; //  146 :  15 - 0xf
      12'h93: dout <= 8'b00011111; //  147 :  31 - 0x1f
      12'h94: dout <= 8'b00111111; //  148 :  63 - 0x3f
      12'h95: dout <= 8'b01111100; //  149 : 124 - 0x7c
      12'h96: dout <= 8'b01110000; //  150 : 112 - 0x70
      12'h97: dout <= 8'b00111000; //  151 :  56 - 0x38
      12'h98: dout <= 8'b11000011; //  152 : 195 - 0xc3 -- plane 1
      12'h99: dout <= 8'b11100011; //  153 : 227 - 0xe3
      12'h9A: dout <= 8'b11001111; //  154 : 207 - 0xcf
      12'h9B: dout <= 8'b00011111; //  155 :  31 - 0x1f
      12'h9C: dout <= 8'b00111111; //  156 :  63 - 0x3f
      12'h9D: dout <= 8'b00001100; //  157 :  12 - 0xc
      12'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b10000000; //  160 : 128 - 0x80 -- Sprite 0xa
      12'hA1: dout <= 8'b11110000; //  161 : 240 - 0xf0
      12'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      12'hA3: dout <= 8'b01000000; //  163 :  64 - 0x40
      12'hA4: dout <= 8'b00100000; //  164 :  32 - 0x20
      12'hA5: dout <= 8'b01111000; //  165 : 120 - 0x78
      12'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout <= 8'b11000000; //  167 : 192 - 0xc0
      12'hA8: dout <= 8'b10000000; //  168 : 128 - 0x80 -- plane 1
      12'hA9: dout <= 8'b11110000; //  169 : 240 - 0xf0
      12'hAA: dout <= 8'b11000000; //  170 : 192 - 0xc0
      12'hAB: dout <= 8'b10111000; //  171 : 184 - 0xb8
      12'hAC: dout <= 8'b11011100; //  172 : 220 - 0xdc
      12'hAD: dout <= 8'b10000000; //  173 : 128 - 0x80
      12'hAE: dout <= 8'b11110000; //  174 : 240 - 0xf0
      12'hAF: dout <= 8'b00000110; //  175 :   6 - 0x6
      12'hB0: dout <= 8'b11110000; //  176 : 240 - 0xf0 -- Sprite 0xb
      12'hB1: dout <= 8'b11111000; //  177 : 248 - 0xf8
      12'hB2: dout <= 8'b11100100; //  178 : 228 - 0xe4
      12'hB3: dout <= 8'b11111100; //  179 : 252 - 0xfc
      12'hB4: dout <= 8'b11111100; //  180 : 252 - 0xfc
      12'hB5: dout <= 8'b01111100; //  181 : 124 - 0x7c
      12'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout <= 8'b10001110; //  184 : 142 - 0x8e -- plane 1
      12'hB9: dout <= 8'b11100110; //  185 : 230 - 0xe6
      12'hBA: dout <= 8'b11100000; //  186 : 224 - 0xe0
      12'hBB: dout <= 8'b11110000; //  187 : 240 - 0xf0
      12'hBC: dout <= 8'b11110000; //  188 : 240 - 0xf0
      12'hBD: dout <= 8'b01110000; //  189 : 112 - 0x70
      12'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      12'hC1: dout <= 8'b00000010; //  193 :   2 - 0x2
      12'hC2: dout <= 8'b00000110; //  194 :   6 - 0x6
      12'hC3: dout <= 8'b00000111; //  195 :   7 - 0x7
      12'hC4: dout <= 8'b00001001; //  196 :   9 - 0x9
      12'hC5: dout <= 8'b00001001; //  197 :   9 - 0x9
      12'hC6: dout <= 8'b00011101; //  198 :  29 - 0x1d
      12'hC7: dout <= 8'b00000011; //  199 :   3 - 0x3
      12'hC8: dout <= 8'b00000001; //  200 :   1 - 0x1 -- plane 1
      12'hC9: dout <= 8'b00000011; //  201 :   3 - 0x3
      12'hCA: dout <= 8'b00000111; //  202 :   7 - 0x7
      12'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout <= 8'b00000110; //  204 :   6 - 0x6
      12'hCD: dout <= 8'b00000110; //  205 :   6 - 0x6
      12'hCE: dout <= 8'b00000010; //  206 :   2 - 0x2
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b00001111; //  208 :  15 - 0xf -- Sprite 0xd
      12'hD1: dout <= 8'b00001111; //  209 :  15 - 0xf
      12'hD2: dout <= 8'b00001111; //  210 :  15 - 0xf
      12'hD3: dout <= 8'b11111111; //  211 : 255 - 0xff
      12'hD4: dout <= 8'b11111111; //  212 : 255 - 0xff
      12'hD5: dout <= 8'b11111100; //  213 : 252 - 0xfc
      12'hD6: dout <= 8'b10000001; //  214 : 129 - 0x81
      12'hD7: dout <= 8'b00000001; //  215 :   1 - 0x1
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- plane 1
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00001100; //  218 :  12 - 0xc
      12'hDB: dout <= 8'b00111111; //  219 :  63 - 0x3f
      12'hDC: dout <= 8'b00111111; //  220 :  63 - 0x3f
      12'hDD: dout <= 8'b00111100; //  221 :  60 - 0x3c
      12'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      12'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      12'hE2: dout <= 8'b00111000; //  226 :  56 - 0x38
      12'hE3: dout <= 8'b11000000; //  227 : 192 - 0xc0
      12'hE4: dout <= 8'b11100000; //  228 : 224 - 0xe0
      12'hE5: dout <= 8'b11010000; //  229 : 208 - 0xd0
      12'hE6: dout <= 8'b11111100; //  230 : 252 - 0xfc
      12'hE7: dout <= 8'b11000000; //  231 : 192 - 0xc0
      12'hE8: dout <= 8'b11000000; //  232 : 192 - 0xc0 -- plane 1
      12'hE9: dout <= 8'b11000000; //  233 : 192 - 0xc0
      12'hEA: dout <= 8'b11111000; //  234 : 248 - 0xf8
      12'hEB: dout <= 8'b00100000; //  235 :  32 - 0x20
      12'hEC: dout <= 8'b00011100; //  236 :  28 - 0x1c
      12'hED: dout <= 8'b00101110; //  237 :  46 - 0x2e
      12'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout <= 8'b00111000; //  239 :  56 - 0x38
      12'hF0: dout <= 8'b11100000; //  240 : 224 - 0xe0 -- Sprite 0xf
      12'hF1: dout <= 8'b11100000; //  241 : 224 - 0xe0
      12'hF2: dout <= 8'b10110000; //  242 : 176 - 0xb0
      12'hF3: dout <= 8'b11110000; //  243 : 240 - 0xf0
      12'hF4: dout <= 8'b11110000; //  244 : 240 - 0xf0
      12'hF5: dout <= 8'b11100000; //  245 : 224 - 0xe0
      12'hF6: dout <= 8'b11000000; //  246 : 192 - 0xc0
      12'hF7: dout <= 8'b11100000; //  247 : 224 - 0xe0
      12'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout <= 8'b01100000; //  249 :  96 - 0x60
      12'hFA: dout <= 8'b11110000; //  250 : 240 - 0xf0
      12'hFB: dout <= 8'b11110000; //  251 : 240 - 0xf0
      12'hFC: dout <= 8'b11110000; //  252 : 240 - 0xf0
      12'hFD: dout <= 8'b11100000; //  253 : 224 - 0xe0
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      12'h101: dout <= 8'b00000011; //  257 :   3 - 0x3
      12'h102: dout <= 8'b00000111; //  258 :   7 - 0x7
      12'h103: dout <= 8'b00000111; //  259 :   7 - 0x7
      12'h104: dout <= 8'b00001001; //  260 :   9 - 0x9
      12'h105: dout <= 8'b00001001; //  261 :   9 - 0x9
      12'h106: dout <= 8'b00011100; //  262 :  28 - 0x1c
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout <= 8'b00000011; //  265 :   3 - 0x3
      12'h10A: dout <= 8'b00000111; //  266 :   7 - 0x7
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000110; //  268 :   6 - 0x6
      12'h10D: dout <= 8'b00000110; //  269 :   6 - 0x6
      12'h10E: dout <= 8'b00000011; //  270 :   3 - 0x3
      12'h10F: dout <= 8'b00000011; //  271 :   3 - 0x3
      12'h110: dout <= 8'b00001111; //  272 :  15 - 0xf -- Sprite 0x11
      12'h111: dout <= 8'b00001111; //  273 :  15 - 0xf
      12'h112: dout <= 8'b00001111; //  274 :  15 - 0xf
      12'h113: dout <= 8'b11111111; //  275 : 255 - 0xff
      12'h114: dout <= 8'b11111111; //  276 : 255 - 0xff
      12'h115: dout <= 8'b11111100; //  277 : 252 - 0xfc
      12'h116: dout <= 8'b10000001; //  278 : 129 - 0x81
      12'h117: dout <= 8'b00000001; //  279 :   1 - 0x1
      12'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout <= 8'b00001100; //  282 :  12 - 0xc
      12'h11B: dout <= 8'b00111111; //  283 :  63 - 0x3f
      12'h11C: dout <= 8'b00111111; //  284 :  63 - 0x3f
      12'h11D: dout <= 8'b00111100; //  285 :  60 - 0x3c
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x12
      12'h121: dout <= 8'b11000000; //  289 : 192 - 0xc0
      12'h122: dout <= 8'b11111000; //  290 : 248 - 0xf8
      12'h123: dout <= 8'b10000000; //  291 : 128 - 0x80
      12'h124: dout <= 8'b00100000; //  292 :  32 - 0x20
      12'h125: dout <= 8'b10010000; //  293 : 144 - 0x90
      12'h126: dout <= 8'b00111100; //  294 :  60 - 0x3c
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout <= 8'b11000000; //  297 : 192 - 0xc0
      12'h12A: dout <= 8'b11111000; //  298 : 248 - 0xf8
      12'h12B: dout <= 8'b01100000; //  299 :  96 - 0x60
      12'h12C: dout <= 8'b11011100; //  300 : 220 - 0xdc
      12'h12D: dout <= 8'b01101110; //  301 : 110 - 0x6e
      12'h12E: dout <= 8'b11000000; //  302 : 192 - 0xc0
      12'h12F: dout <= 8'b11111000; //  303 : 248 - 0xf8
      12'h130: dout <= 8'b11100000; //  304 : 224 - 0xe0 -- Sprite 0x13
      12'h131: dout <= 8'b11110000; //  305 : 240 - 0xf0
      12'h132: dout <= 8'b11110000; //  306 : 240 - 0xf0
      12'h133: dout <= 8'b11110000; //  307 : 240 - 0xf0
      12'h134: dout <= 8'b11110000; //  308 : 240 - 0xf0
      12'h135: dout <= 8'b11100000; //  309 : 224 - 0xe0
      12'h136: dout <= 8'b11000000; //  310 : 192 - 0xc0
      12'h137: dout <= 8'b11100000; //  311 : 224 - 0xe0
      12'h138: dout <= 8'b01000111; //  312 :  71 - 0x47 -- plane 1
      12'h139: dout <= 8'b00001111; //  313 :  15 - 0xf
      12'h13A: dout <= 8'b00001110; //  314 :  14 - 0xe
      12'h13B: dout <= 8'b11110000; //  315 : 240 - 0xf0
      12'h13C: dout <= 8'b11110000; //  316 : 240 - 0xf0
      12'h13D: dout <= 8'b11100000; //  317 : 224 - 0xe0
      12'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b00000100; //  320 :   4 - 0x4 -- Sprite 0x14
      12'h141: dout <= 8'b00001100; //  321 :  12 - 0xc
      12'h142: dout <= 8'b00001100; //  322 :  12 - 0xc
      12'h143: dout <= 8'b00010011; //  323 :  19 - 0x13
      12'h144: dout <= 8'b00010011; //  324 :  19 - 0x13
      12'h145: dout <= 8'b00111011; //  325 :  59 - 0x3b
      12'h146: dout <= 8'b00000111; //  326 :   7 - 0x7
      12'h147: dout <= 8'b00001111; //  327 :  15 - 0xf
      12'h148: dout <= 8'b00000111; //  328 :   7 - 0x7 -- plane 1
      12'h149: dout <= 8'b00001111; //  329 :  15 - 0xf
      12'h14A: dout <= 8'b00000011; //  330 :   3 - 0x3
      12'h14B: dout <= 8'b00001100; //  331 :  12 - 0xc
      12'h14C: dout <= 8'b00001100; //  332 :  12 - 0xc
      12'h14D: dout <= 8'b00000100; //  333 :   4 - 0x4
      12'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout <= 8'b00001111; //  336 :  15 - 0xf -- Sprite 0x15
      12'h151: dout <= 8'b00001111; //  337 :  15 - 0xf
      12'h152: dout <= 8'b00001111; //  338 :  15 - 0xf
      12'h153: dout <= 8'b00011111; //  339 :  31 - 0x1f
      12'h154: dout <= 8'b00011111; //  340 :  31 - 0x1f
      12'h155: dout <= 8'b00011110; //  341 :  30 - 0x1e
      12'h156: dout <= 8'b00011100; //  342 :  28 - 0x1c
      12'h157: dout <= 8'b00011110; //  343 :  30 - 0x1e
      12'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- plane 1
      12'h159: dout <= 8'b00000001; //  345 :   1 - 0x1
      12'h15A: dout <= 8'b00001111; //  346 :  15 - 0xf
      12'h15B: dout <= 8'b00011111; //  347 :  31 - 0x1f
      12'h15C: dout <= 8'b00011111; //  348 :  31 - 0x1f
      12'h15D: dout <= 8'b00011110; //  349 :  30 - 0x1e
      12'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      12'h161: dout <= 8'b01110000; //  353 : 112 - 0x70
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b11000000; //  355 : 192 - 0xc0
      12'h164: dout <= 8'b10100000; //  356 : 160 - 0xa0
      12'h165: dout <= 8'b11111000; //  357 : 248 - 0xf8
      12'h166: dout <= 8'b10000000; //  358 : 128 - 0x80
      12'h167: dout <= 8'b11000000; //  359 : 192 - 0xc0
      12'h168: dout <= 8'b10000000; //  360 : 128 - 0x80 -- plane 1
      12'h169: dout <= 8'b11110000; //  361 : 240 - 0xf0
      12'h16A: dout <= 8'b11000000; //  362 : 192 - 0xc0
      12'h16B: dout <= 8'b00111000; //  363 :  56 - 0x38
      12'h16C: dout <= 8'b01011100; //  364 :  92 - 0x5c
      12'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout <= 8'b01110000; //  366 : 112 - 0x70
      12'h16F: dout <= 8'b01000000; //  367 :  64 - 0x40
      12'h170: dout <= 8'b11100000; //  368 : 224 - 0xe0 -- Sprite 0x17
      12'h171: dout <= 8'b01100000; //  369 :  96 - 0x60
      12'h172: dout <= 8'b11110000; //  370 : 240 - 0xf0
      12'h173: dout <= 8'b11110000; //  371 : 240 - 0xf0
      12'h174: dout <= 8'b11110000; //  372 : 240 - 0xf0
      12'h175: dout <= 8'b11100000; //  373 : 224 - 0xe0
      12'h176: dout <= 8'b11100000; //  374 : 224 - 0xe0
      12'h177: dout <= 8'b11110000; //  375 : 240 - 0xf0
      12'h178: dout <= 8'b11000000; //  376 : 192 - 0xc0 -- plane 1
      12'h179: dout <= 8'b11100000; //  377 : 224 - 0xe0
      12'h17A: dout <= 8'b11110000; //  378 : 240 - 0xf0
      12'h17B: dout <= 8'b11110000; //  379 : 240 - 0xf0
      12'h17C: dout <= 8'b11110000; //  380 : 240 - 0xf0
      12'h17D: dout <= 8'b11100000; //  381 : 224 - 0xe0
      12'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00000111; //  384 :   7 - 0x7 -- Sprite 0x18
      12'h181: dout <= 8'b00001111; //  385 :  15 - 0xf
      12'h182: dout <= 8'b00001111; //  386 :  15 - 0xf
      12'h183: dout <= 8'b00010010; //  387 :  18 - 0x12
      12'h184: dout <= 8'b00010011; //  388 :  19 - 0x13
      12'h185: dout <= 8'b00111000; //  389 :  56 - 0x38
      12'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      12'h187: dout <= 8'b00001111; //  391 :  15 - 0xf
      12'h188: dout <= 8'b00000111; //  392 :   7 - 0x7 -- plane 1
      12'h189: dout <= 8'b00001111; //  393 :  15 - 0xf
      12'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout <= 8'b00001101; //  395 :  13 - 0xd
      12'h18C: dout <= 8'b00001100; //  396 :  12 - 0xc
      12'h18D: dout <= 8'b00000111; //  397 :   7 - 0x7
      12'h18E: dout <= 8'b00000111; //  398 :   7 - 0x7
      12'h18F: dout <= 8'b00000001; //  399 :   1 - 0x1
      12'h190: dout <= 8'b00011111; //  400 :  31 - 0x1f -- Sprite 0x19
      12'h191: dout <= 8'b00011111; //  401 :  31 - 0x1f
      12'h192: dout <= 8'b00011111; //  402 :  31 - 0x1f
      12'h193: dout <= 8'b00011111; //  403 :  31 - 0x1f
      12'h194: dout <= 8'b00011111; //  404 :  31 - 0x1f
      12'h195: dout <= 8'b00011110; //  405 :  30 - 0x1e
      12'h196: dout <= 8'b00011100; //  406 :  28 - 0x1c
      12'h197: dout <= 8'b00011110; //  407 :  30 - 0x1e
      12'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout <= 8'b00010011; //  410 :  19 - 0x13
      12'h19B: dout <= 8'b00011111; //  411 :  31 - 0x1f
      12'h19C: dout <= 8'b00011111; //  412 :  31 - 0x1f
      12'h19D: dout <= 8'b00011110; //  413 :  30 - 0x1e
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b10000000; //  416 : 128 - 0x80 -- Sprite 0x1a
      12'h1A1: dout <= 8'b11110000; //  417 : 240 - 0xf0
      12'h1A2: dout <= 8'b00000000; //  418 :   0 - 0x0
      12'h1A3: dout <= 8'b01000000; //  419 :  64 - 0x40
      12'h1A4: dout <= 8'b00100000; //  420 :  32 - 0x20
      12'h1A5: dout <= 8'b01111000; //  421 : 120 - 0x78
      12'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      12'h1A7: dout <= 8'b11000000; //  423 : 192 - 0xc0
      12'h1A8: dout <= 8'b10000000; //  424 : 128 - 0x80 -- plane 1
      12'h1A9: dout <= 8'b11110000; //  425 : 240 - 0xf0
      12'h1AA: dout <= 8'b11000000; //  426 : 192 - 0xc0
      12'h1AB: dout <= 8'b10111000; //  427 : 184 - 0xb8
      12'h1AC: dout <= 8'b11011100; //  428 : 220 - 0xdc
      12'h1AD: dout <= 8'b10000000; //  429 : 128 - 0x80
      12'h1AE: dout <= 8'b11110000; //  430 : 240 - 0xf0
      12'h1AF: dout <= 8'b10000000; //  431 : 128 - 0x80
      12'h1B0: dout <= 8'b11111000; //  432 : 248 - 0xf8 -- Sprite 0x1b
      12'h1B1: dout <= 8'b11111000; //  433 : 248 - 0xf8
      12'h1B2: dout <= 8'b11110000; //  434 : 240 - 0xf0
      12'h1B3: dout <= 8'b11110000; //  435 : 240 - 0xf0
      12'h1B4: dout <= 8'b11110000; //  436 : 240 - 0xf0
      12'h1B5: dout <= 8'b11100000; //  437 : 224 - 0xe0
      12'h1B6: dout <= 8'b11100000; //  438 : 224 - 0xe0
      12'h1B7: dout <= 8'b11110000; //  439 : 240 - 0xf0
      12'h1B8: dout <= 8'b00000111; //  440 :   7 - 0x7 -- plane 1
      12'h1B9: dout <= 8'b00000111; //  441 :   7 - 0x7
      12'h1BA: dout <= 8'b11111110; //  442 : 254 - 0xfe
      12'h1BB: dout <= 8'b11110000; //  443 : 240 - 0xf0
      12'h1BC: dout <= 8'b11110000; //  444 : 240 - 0xf0
      12'h1BD: dout <= 8'b11100000; //  445 : 224 - 0xe0
      12'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b00000100; //  448 :   4 - 0x4 -- Sprite 0x1c
      12'h1C1: dout <= 8'b00001100; //  449 :  12 - 0xc
      12'h1C2: dout <= 8'b00001100; //  450 :  12 - 0xc
      12'h1C3: dout <= 8'b00010011; //  451 :  19 - 0x13
      12'h1C4: dout <= 8'b00010011; //  452 :  19 - 0x13
      12'h1C5: dout <= 8'b00111111; //  453 :  63 - 0x3f
      12'h1C6: dout <= 8'b00000111; //  454 :   7 - 0x7
      12'h1C7: dout <= 8'b00001111; //  455 :  15 - 0xf
      12'h1C8: dout <= 8'b00000111; //  456 :   7 - 0x7 -- plane 1
      12'h1C9: dout <= 8'b00001111; //  457 :  15 - 0xf
      12'h1CA: dout <= 8'b00000011; //  458 :   3 - 0x3
      12'h1CB: dout <= 8'b00001100; //  459 :  12 - 0xc
      12'h1CC: dout <= 8'b00001100; //  460 :  12 - 0xc
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00001111; //  464 :  15 - 0xf -- Sprite 0x1d
      12'h1D1: dout <= 8'b00001111; //  465 :  15 - 0xf
      12'h1D2: dout <= 8'b00001111; //  466 :  15 - 0xf
      12'h1D3: dout <= 8'b00011111; //  467 :  31 - 0x1f
      12'h1D4: dout <= 8'b00111111; //  468 :  63 - 0x3f
      12'h1D5: dout <= 8'b01111100; //  469 : 124 - 0x7c
      12'h1D6: dout <= 8'b01110000; //  470 : 112 - 0x70
      12'h1D7: dout <= 8'b00111000; //  471 :  56 - 0x38
      12'h1D8: dout <= 8'b00000001; //  472 :   1 - 0x1 -- plane 1
      12'h1D9: dout <= 8'b00000001; //  473 :   1 - 0x1
      12'h1DA: dout <= 8'b00001111; //  474 :  15 - 0xf
      12'h1DB: dout <= 8'b00011111; //  475 :  31 - 0x1f
      12'h1DC: dout <= 8'b00111111; //  476 :  63 - 0x3f
      12'h1DD: dout <= 8'b00011100; //  477 :  28 - 0x1c
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x1e
      12'h1E1: dout <= 8'b01110000; //  481 : 112 - 0x70
      12'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout <= 8'b11000000; //  483 : 192 - 0xc0
      12'h1E4: dout <= 8'b10100000; //  484 : 160 - 0xa0
      12'h1E5: dout <= 8'b11111000; //  485 : 248 - 0xf8
      12'h1E6: dout <= 8'b10000000; //  486 : 128 - 0x80
      12'h1E7: dout <= 8'b11000000; //  487 : 192 - 0xc0
      12'h1E8: dout <= 8'b10000000; //  488 : 128 - 0x80 -- plane 1
      12'h1E9: dout <= 8'b11110000; //  489 : 240 - 0xf0
      12'h1EA: dout <= 8'b11000000; //  490 : 192 - 0xc0
      12'h1EB: dout <= 8'b00111000; //  491 :  56 - 0x38
      12'h1EC: dout <= 8'b01011100; //  492 :  92 - 0x5c
      12'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout <= 8'b01110000; //  494 : 112 - 0x70
      12'h1EF: dout <= 8'b01000000; //  495 :  64 - 0x40
      12'h1F0: dout <= 8'b11000000; //  496 : 192 - 0xc0 -- Sprite 0x1f
      12'h1F1: dout <= 8'b01100000; //  497 :  96 - 0x60
      12'h1F2: dout <= 8'b11100100; //  498 : 228 - 0xe4
      12'h1F3: dout <= 8'b11111100; //  499 : 252 - 0xfc
      12'h1F4: dout <= 8'b11111100; //  500 : 252 - 0xfc
      12'h1F5: dout <= 8'b01111100; //  501 : 124 - 0x7c
      12'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout <= 8'b11000000; //  504 : 192 - 0xc0 -- plane 1
      12'h1F9: dout <= 8'b11100000; //  505 : 224 - 0xe0
      12'h1FA: dout <= 8'b11100000; //  506 : 224 - 0xe0
      12'h1FB: dout <= 8'b11110000; //  507 : 240 - 0xf0
      12'h1FC: dout <= 8'b11110000; //  508 : 240 - 0xf0
      12'h1FD: dout <= 8'b01110000; //  509 : 112 - 0x70
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000111; //  512 :   7 - 0x7 -- Sprite 0x20
      12'h201: dout <= 8'b00001111; //  513 :  15 - 0xf
      12'h202: dout <= 8'b00001111; //  514 :  15 - 0xf
      12'h203: dout <= 8'b00010010; //  515 :  18 - 0x12
      12'h204: dout <= 8'b00010011; //  516 :  19 - 0x13
      12'h205: dout <= 8'b00111000; //  517 :  56 - 0x38
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000111; //  519 :   7 - 0x7
      12'h208: dout <= 8'b00000111; //  520 :   7 - 0x7 -- plane 1
      12'h209: dout <= 8'b00001111; //  521 :  15 - 0xf
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00001101; //  523 :  13 - 0xd
      12'h20C: dout <= 8'b00001100; //  524 :  12 - 0xc
      12'h20D: dout <= 8'b00000111; //  525 :   7 - 0x7
      12'h20E: dout <= 8'b00000111; //  526 :   7 - 0x7
      12'h20F: dout <= 8'b00000001; //  527 :   1 - 0x1
      12'h210: dout <= 8'b00001111; //  528 :  15 - 0xf -- Sprite 0x21
      12'h211: dout <= 8'b00001111; //  529 :  15 - 0xf
      12'h212: dout <= 8'b00001111; //  530 :  15 - 0xf
      12'h213: dout <= 8'b00011111; //  531 :  31 - 0x1f
      12'h214: dout <= 8'b00111111; //  532 :  63 - 0x3f
      12'h215: dout <= 8'b01111100; //  533 : 124 - 0x7c
      12'h216: dout <= 8'b01110000; //  534 : 112 - 0x70
      12'h217: dout <= 8'b00111000; //  535 :  56 - 0x38
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout <= 8'b00001001; //  538 :   9 - 0x9
      12'h21B: dout <= 8'b00011111; //  539 :  31 - 0x1f
      12'h21C: dout <= 8'b00111111; //  540 :  63 - 0x3f
      12'h21D: dout <= 8'b00011100; //  541 :  28 - 0x1c
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b10000000; //  544 : 128 - 0x80 -- Sprite 0x22
      12'h221: dout <= 8'b11110000; //  545 : 240 - 0xf0
      12'h222: dout <= 8'b00000000; //  546 :   0 - 0x0
      12'h223: dout <= 8'b01000000; //  547 :  64 - 0x40
      12'h224: dout <= 8'b00100000; //  548 :  32 - 0x20
      12'h225: dout <= 8'b01111000; //  549 : 120 - 0x78
      12'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      12'h227: dout <= 8'b11000000; //  551 : 192 - 0xc0
      12'h228: dout <= 8'b10000000; //  552 : 128 - 0x80 -- plane 1
      12'h229: dout <= 8'b11110000; //  553 : 240 - 0xf0
      12'h22A: dout <= 8'b11000000; //  554 : 192 - 0xc0
      12'h22B: dout <= 8'b10111000; //  555 : 184 - 0xb8
      12'h22C: dout <= 8'b11011100; //  556 : 220 - 0xdc
      12'h22D: dout <= 8'b10000000; //  557 : 128 - 0x80
      12'h22E: dout <= 8'b11110000; //  558 : 240 - 0xf0
      12'h22F: dout <= 8'b10000000; //  559 : 128 - 0x80
      12'h230: dout <= 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x23
      12'h231: dout <= 8'b11111000; //  561 : 248 - 0xf8
      12'h232: dout <= 8'b11100000; //  562 : 224 - 0xe0
      12'h233: dout <= 8'b11111100; //  563 : 252 - 0xfc
      12'h234: dout <= 8'b11111100; //  564 : 252 - 0xfc
      12'h235: dout <= 8'b01111100; //  565 : 124 - 0x7c
      12'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00000111; //  568 :   7 - 0x7 -- plane 1
      12'h239: dout <= 8'b00000111; //  569 :   7 - 0x7
      12'h23A: dout <= 8'b11101110; //  570 : 238 - 0xee
      12'h23B: dout <= 8'b11110000; //  571 : 240 - 0xf0
      12'h23C: dout <= 8'b11110000; //  572 : 240 - 0xf0
      12'h23D: dout <= 8'b01110000; //  573 : 112 - 0x70
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      12'h241: dout <= 8'b00000111; //  577 :   7 - 0x7
      12'h242: dout <= 8'b00000111; //  578 :   7 - 0x7
      12'h243: dout <= 8'b00001111; //  579 :  15 - 0xf
      12'h244: dout <= 8'b00001111; //  580 :  15 - 0xf
      12'h245: dout <= 8'b00111000; //  581 :  56 - 0x38
      12'h246: dout <= 8'b01111111; //  582 : 127 - 0x7f
      12'h247: dout <= 8'b01111111; //  583 : 127 - 0x7f
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- plane 1
      12'h249: dout <= 8'b00000111; //  585 :   7 - 0x7
      12'h24A: dout <= 8'b00000011; //  586 :   3 - 0x3
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000111; //  589 :   7 - 0x7
      12'h24E: dout <= 8'b00000100; //  590 :   4 - 0x4
      12'h24F: dout <= 8'b00000100; //  591 :   4 - 0x4
      12'h250: dout <= 8'b00011111; //  592 :  31 - 0x1f -- Sprite 0x25
      12'h251: dout <= 8'b00011111; //  593 :  31 - 0x1f
      12'h252: dout <= 8'b00011111; //  594 :  31 - 0x1f
      12'h253: dout <= 8'b00011111; //  595 :  31 - 0x1f
      12'h254: dout <= 8'b00001111; //  596 :  15 - 0xf
      12'h255: dout <= 8'b00001111; //  597 :  15 - 0xf
      12'h256: dout <= 8'b00001111; //  598 :  15 - 0xf
      12'h257: dout <= 8'b00000111; //  599 :   7 - 0x7
      12'h258: dout <= 8'b00011110; //  600 :  30 - 0x1e -- plane 1
      12'h259: dout <= 8'b00011111; //  601 :  31 - 0x1f
      12'h25A: dout <= 8'b00011111; //  602 :  31 - 0x1f
      12'h25B: dout <= 8'b00011111; //  603 :  31 - 0x1f
      12'h25C: dout <= 8'b00001111; //  604 :  15 - 0xf
      12'h25D: dout <= 8'b00001000; //  605 :   8 - 0x8
      12'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      12'h261: dout <= 8'b11100000; //  609 : 224 - 0xe0
      12'h262: dout <= 8'b11111000; //  610 : 248 - 0xf8
      12'h263: dout <= 8'b11111100; //  611 : 252 - 0xfc
      12'h264: dout <= 8'b11111100; //  612 : 252 - 0xfc
      12'h265: dout <= 8'b00011100; //  613 :  28 - 0x1c
      12'h266: dout <= 8'b11111000; //  614 : 248 - 0xf8
      12'h267: dout <= 8'b11111000; //  615 : 248 - 0xf8
      12'h268: dout <= 8'b00111000; //  616 :  56 - 0x38 -- plane 1
      12'h269: dout <= 8'b11111000; //  617 : 248 - 0xf8
      12'h26A: dout <= 8'b11000000; //  618 : 192 - 0xc0
      12'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b11100000; //  621 : 224 - 0xe0
      12'h26E: dout <= 8'b00100000; //  622 :  32 - 0x20
      12'h26F: dout <= 8'b00100000; //  623 :  32 - 0x20
      12'h270: dout <= 8'b11111000; //  624 : 248 - 0xf8 -- Sprite 0x27
      12'h271: dout <= 8'b11111100; //  625 : 252 - 0xfc
      12'h272: dout <= 8'b11111100; //  626 : 252 - 0xfc
      12'h273: dout <= 8'b11111000; //  627 : 248 - 0xf8
      12'h274: dout <= 8'b01111000; //  628 : 120 - 0x78
      12'h275: dout <= 8'b10000000; //  629 : 128 - 0x80
      12'h276: dout <= 8'b11000000; //  630 : 192 - 0xc0
      12'h277: dout <= 8'b11000000; //  631 : 192 - 0xc0
      12'h278: dout <= 8'b01111000; //  632 : 120 - 0x78 -- plane 1
      12'h279: dout <= 8'b11111100; //  633 : 252 - 0xfc
      12'h27A: dout <= 8'b11111100; //  634 : 252 - 0xfc
      12'h27B: dout <= 8'b11111000; //  635 : 248 - 0xf8
      12'h27C: dout <= 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout <= 8'b10000000; //  637 : 128 - 0x80
      12'h27E: dout <= 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      12'h281: dout <= 8'b00000011; //  641 :   3 - 0x3
      12'h282: dout <= 8'b00000111; //  642 :   7 - 0x7
      12'h283: dout <= 8'b00000111; //  643 :   7 - 0x7
      12'h284: dout <= 8'b00001001; //  644 :   9 - 0x9
      12'h285: dout <= 8'b00001001; //  645 :   9 - 0x9
      12'h286: dout <= 8'b00011100; //  646 :  28 - 0x1c
      12'h287: dout <= 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout <= 8'b00000011; //  649 :   3 - 0x3
      12'h28A: dout <= 8'b00000111; //  650 :   7 - 0x7
      12'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout <= 8'b00000110; //  652 :   6 - 0x6
      12'h28D: dout <= 8'b00000110; //  653 :   6 - 0x6
      12'h28E: dout <= 8'b00000011; //  654 :   3 - 0x3
      12'h28F: dout <= 8'b01100011; //  655 :  99 - 0x63
      12'h290: dout <= 8'b00011111; //  656 :  31 - 0x1f -- Sprite 0x29
      12'h291: dout <= 8'b00001111; //  657 :  15 - 0xf
      12'h292: dout <= 8'b00000111; //  658 :   7 - 0x7
      12'h293: dout <= 8'b00110111; //  659 :  55 - 0x37
      12'h294: dout <= 8'b01111111; //  660 : 127 - 0x7f
      12'h295: dout <= 8'b11011111; //  661 : 223 - 0xdf
      12'h296: dout <= 8'b00001111; //  662 :  15 - 0xf
      12'h297: dout <= 8'b00000110; //  663 :   6 - 0x6
      12'h298: dout <= 8'b11100000; //  664 : 224 - 0xe0 -- plane 1
      12'h299: dout <= 8'b00100001; //  665 :  33 - 0x21
      12'h29A: dout <= 8'b00000001; //  666 :   1 - 0x1
      12'h29B: dout <= 8'b00000111; //  667 :   7 - 0x7
      12'h29C: dout <= 8'b00000111; //  668 :   7 - 0x7
      12'h29D: dout <= 8'b00011111; //  669 :  31 - 0x1f
      12'h29E: dout <= 8'b00001111; //  670 :  15 - 0xf
      12'h29F: dout <= 8'b00000110; //  671 :   6 - 0x6
      12'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x2a
      12'h2A1: dout <= 8'b11000000; //  673 : 192 - 0xc0
      12'h2A2: dout <= 8'b11111000; //  674 : 248 - 0xf8
      12'h2A3: dout <= 8'b10000000; //  675 : 128 - 0x80
      12'h2A4: dout <= 8'b00100000; //  676 :  32 - 0x20
      12'h2A5: dout <= 8'b10010000; //  677 : 144 - 0x90
      12'h2A6: dout <= 8'b00111100; //  678 :  60 - 0x3c
      12'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- plane 1
      12'h2A9: dout <= 8'b11000000; //  681 : 192 - 0xc0
      12'h2AA: dout <= 8'b11111000; //  682 : 248 - 0xf8
      12'h2AB: dout <= 8'b01100000; //  683 :  96 - 0x60
      12'h2AC: dout <= 8'b11011100; //  684 : 220 - 0xdc
      12'h2AD: dout <= 8'b01101110; //  685 : 110 - 0x6e
      12'h2AE: dout <= 8'b11000000; //  686 : 192 - 0xc0
      12'h2AF: dout <= 8'b11111011; //  687 : 251 - 0xfb
      12'h2B0: dout <= 8'b11100100; //  688 : 228 - 0xe4 -- Sprite 0x2b
      12'h2B1: dout <= 8'b11111110; //  689 : 254 - 0xfe
      12'h2B2: dout <= 8'b01110000; //  690 : 112 - 0x70
      12'h2B3: dout <= 8'b11110001; //  691 : 241 - 0xf1
      12'h2B4: dout <= 8'b11111111; //  692 : 255 - 0xff
      12'h2B5: dout <= 8'b11111111; //  693 : 255 - 0xff
      12'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout <= 8'b10000011; //  696 : 131 - 0x83 -- plane 1
      12'h2B9: dout <= 8'b11000000; //  697 : 192 - 0xc0
      12'h2BA: dout <= 8'b11110000; //  698 : 240 - 0xf0
      12'h2BB: dout <= 8'b11110000; //  699 : 240 - 0xf0
      12'h2BC: dout <= 8'b11111100; //  700 : 252 - 0xfc
      12'h2BD: dout <= 8'b11111100; //  701 : 252 - 0xfc
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b00000111; //  704 :   7 - 0x7 -- Sprite 0x2c
      12'h2C1: dout <= 8'b00001111; //  705 :  15 - 0xf
      12'h2C2: dout <= 8'b00001111; //  706 :  15 - 0xf
      12'h2C3: dout <= 8'b00010010; //  707 :  18 - 0x12
      12'h2C4: dout <= 8'b00010011; //  708 :  19 - 0x13
      12'h2C5: dout <= 8'b00111000; //  709 :  56 - 0x38
      12'h2C6: dout <= 8'b01110000; //  710 : 112 - 0x70
      12'h2C7: dout <= 8'b11111111; //  711 : 255 - 0xff
      12'h2C8: dout <= 8'b00000111; //  712 :   7 - 0x7 -- plane 1
      12'h2C9: dout <= 8'b00001111; //  713 :  15 - 0xf
      12'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout <= 8'b00001101; //  715 :  13 - 0xd
      12'h2CC: dout <= 8'b00001100; //  716 :  12 - 0xc
      12'h2CD: dout <= 8'b00000111; //  717 :   7 - 0x7
      12'h2CE: dout <= 8'b00001111; //  718 :  15 - 0xf
      12'h2CF: dout <= 8'b00000010; //  719 :   2 - 0x2
      12'h2D0: dout <= 8'b11011111; //  720 : 223 - 0xdf -- Sprite 0x2d
      12'h2D1: dout <= 8'b00011110; //  721 :  30 - 0x1e
      12'h2D2: dout <= 8'b00011111; //  722 :  31 - 0x1f
      12'h2D3: dout <= 8'b00011111; //  723 :  31 - 0x1f
      12'h2D4: dout <= 8'b00011111; //  724 :  31 - 0x1f
      12'h2D5: dout <= 8'b00001111; //  725 :  15 - 0xf
      12'h2D6: dout <= 8'b00000111; //  726 :   7 - 0x7
      12'h2D7: dout <= 8'b00000001; //  727 :   1 - 0x1
      12'h2D8: dout <= 8'b00000001; //  728 :   1 - 0x1 -- plane 1
      12'h2D9: dout <= 8'b11110011; //  729 : 243 - 0xf3
      12'h2DA: dout <= 8'b01011111; //  730 :  95 - 0x5f
      12'h2DB: dout <= 8'b00011111; //  731 :  31 - 0x1f
      12'h2DC: dout <= 8'b00011111; //  732 :  31 - 0x1f
      12'h2DD: dout <= 8'b01001111; //  733 :  79 - 0x4f
      12'h2DE: dout <= 8'b00110111; //  734 :  55 - 0x37
      12'h2DF: dout <= 8'b11000000; //  735 : 192 - 0xc0
      12'h2E0: dout <= 8'b10000000; //  736 : 128 - 0x80 -- Sprite 0x2e
      12'h2E1: dout <= 8'b11110000; //  737 : 240 - 0xf0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b01000000; //  739 :  64 - 0x40
      12'h2E4: dout <= 8'b00100000; //  740 :  32 - 0x20
      12'h2E5: dout <= 8'b01111000; //  741 : 120 - 0x78
      12'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout <= 8'b11111100; //  743 : 252 - 0xfc
      12'h2E8: dout <= 8'b10000000; //  744 : 128 - 0x80 -- plane 1
      12'h2E9: dout <= 8'b11110000; //  745 : 240 - 0xf0
      12'h2EA: dout <= 8'b11000000; //  746 : 192 - 0xc0
      12'h2EB: dout <= 8'b10111000; //  747 : 184 - 0xb8
      12'h2EC: dout <= 8'b11011100; //  748 : 220 - 0xdc
      12'h2ED: dout <= 8'b10000000; //  749 : 128 - 0x80
      12'h2EE: dout <= 8'b11110000; //  750 : 240 - 0xf0
      12'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout <= 8'b11110000; //  752 : 240 - 0xf0 -- Sprite 0x2f
      12'h2F1: dout <= 8'b11100000; //  753 : 224 - 0xe0
      12'h2F2: dout <= 8'b11100000; //  754 : 224 - 0xe0
      12'h2F3: dout <= 8'b11110000; //  755 : 240 - 0xf0
      12'h2F4: dout <= 8'b11111010; //  756 : 250 - 0xfa
      12'h2F5: dout <= 8'b11111110; //  757 : 254 - 0xfe
      12'h2F6: dout <= 8'b11111100; //  758 : 252 - 0xfc
      12'h2F7: dout <= 8'b11011000; //  759 : 216 - 0xd8
      12'h2F8: dout <= 8'b10001111; //  760 : 143 - 0x8f -- plane 1
      12'h2F9: dout <= 8'b11100111; //  761 : 231 - 0xe7
      12'h2FA: dout <= 8'b11100000; //  762 : 224 - 0xe0
      12'h2FB: dout <= 8'b11110000; //  763 : 240 - 0xf0
      12'h2FC: dout <= 8'b11001000; //  764 : 200 - 0xc8
      12'h2FD: dout <= 8'b10001000; //  765 : 136 - 0x88
      12'h2FE: dout <= 8'b00010000; //  766 :  16 - 0x10
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x30
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b00000111; //  770 :   7 - 0x7
      12'h303: dout <= 8'b00001000; //  771 :   8 - 0x8
      12'h304: dout <= 8'b00010000; //  772 :  16 - 0x10
      12'h305: dout <= 8'b00100000; //  773 :  32 - 0x20
      12'h306: dout <= 8'b01000000; //  774 :  64 - 0x40
      12'h307: dout <= 8'b01000000; //  775 :  64 - 0x40
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- plane 1
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      12'h30B: dout <= 8'b00000111; //  779 :   7 - 0x7
      12'h30C: dout <= 8'b00001000; //  780 :   8 - 0x8
      12'h30D: dout <= 8'b00010000; //  781 :  16 - 0x10
      12'h30E: dout <= 8'b00100000; //  782 :  32 - 0x20
      12'h30F: dout <= 8'b00100000; //  783 :  32 - 0x20
      12'h310: dout <= 8'b01000000; //  784 :  64 - 0x40 -- Sprite 0x31
      12'h311: dout <= 8'b01000000; //  785 :  64 - 0x40
      12'h312: dout <= 8'b00100000; //  786 :  32 - 0x20
      12'h313: dout <= 8'b00010000; //  787 :  16 - 0x10
      12'h314: dout <= 8'b00001000; //  788 :   8 - 0x8
      12'h315: dout <= 8'b00000111; //  789 :   7 - 0x7
      12'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b00100000; //  792 :  32 - 0x20 -- plane 1
      12'h319: dout <= 8'b00100000; //  793 :  32 - 0x20
      12'h31A: dout <= 8'b00010000; //  794 :  16 - 0x10
      12'h31B: dout <= 8'b00001000; //  795 :   8 - 0x8
      12'h31C: dout <= 8'b00000111; //  796 :   7 - 0x7
      12'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      12'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout <= 8'b11100000; //  802 : 224 - 0xe0
      12'h323: dout <= 8'b00010000; //  803 :  16 - 0x10
      12'h324: dout <= 8'b00001000; //  804 :   8 - 0x8
      12'h325: dout <= 8'b00000100; //  805 :   4 - 0x4
      12'h326: dout <= 8'b00000010; //  806 :   2 - 0x2
      12'h327: dout <= 8'b00000010; //  807 :   2 - 0x2
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b11100000; //  811 : 224 - 0xe0
      12'h32C: dout <= 8'b00010000; //  812 :  16 - 0x10
      12'h32D: dout <= 8'b00001000; //  813 :   8 - 0x8
      12'h32E: dout <= 8'b00000100; //  814 :   4 - 0x4
      12'h32F: dout <= 8'b00000100; //  815 :   4 - 0x4
      12'h330: dout <= 8'b00000010; //  816 :   2 - 0x2 -- Sprite 0x33
      12'h331: dout <= 8'b00000010; //  817 :   2 - 0x2
      12'h332: dout <= 8'b00000100; //  818 :   4 - 0x4
      12'h333: dout <= 8'b00001000; //  819 :   8 - 0x8
      12'h334: dout <= 8'b00010000; //  820 :  16 - 0x10
      12'h335: dout <= 8'b11100000; //  821 : 224 - 0xe0
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b00000100; //  824 :   4 - 0x4 -- plane 1
      12'h339: dout <= 8'b00000100; //  825 :   4 - 0x4
      12'h33A: dout <= 8'b00001000; //  826 :   8 - 0x8
      12'h33B: dout <= 8'b00010000; //  827 :  16 - 0x10
      12'h33C: dout <= 8'b11100000; //  828 : 224 - 0xe0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout <= 8'b00000011; //  836 :   3 - 0x3
      12'h345: dout <= 8'b00000100; //  837 :   4 - 0x4
      12'h346: dout <= 8'b00001000; //  838 :   8 - 0x8
      12'h347: dout <= 8'b00010000; //  839 :  16 - 0x10
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000011; //  845 :   3 - 0x3
      12'h34E: dout <= 8'b00000100; //  846 :   4 - 0x4
      12'h34F: dout <= 8'b00001000; //  847 :   8 - 0x8
      12'h350: dout <= 8'b00010000; //  848 :  16 - 0x10 -- Sprite 0x35
      12'h351: dout <= 8'b00001000; //  849 :   8 - 0x8
      12'h352: dout <= 8'b00000100; //  850 :   4 - 0x4
      12'h353: dout <= 8'b00000011; //  851 :   3 - 0x3
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00001000; //  856 :   8 - 0x8 -- plane 1
      12'h359: dout <= 8'b00000100; //  857 :   4 - 0x4
      12'h35A: dout <= 8'b00000011; //  858 :   3 - 0x3
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      12'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout <= 8'b11000000; //  868 : 192 - 0xc0
      12'h365: dout <= 8'b00100000; //  869 :  32 - 0x20
      12'h366: dout <= 8'b00010000; //  870 :  16 - 0x10
      12'h367: dout <= 8'b00001000; //  871 :   8 - 0x8
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b11000000; //  877 : 192 - 0xc0
      12'h36E: dout <= 8'b00100000; //  878 :  32 - 0x20
      12'h36F: dout <= 8'b00010000; //  879 :  16 - 0x10
      12'h370: dout <= 8'b00001000; //  880 :   8 - 0x8 -- Sprite 0x37
      12'h371: dout <= 8'b00010000; //  881 :  16 - 0x10
      12'h372: dout <= 8'b00100000; //  882 :  32 - 0x20
      12'h373: dout <= 8'b11000000; //  883 : 192 - 0xc0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b00010000; //  888 :  16 - 0x10 -- plane 1
      12'h379: dout <= 8'b00100000; //  889 :  32 - 0x20
      12'h37A: dout <= 8'b11000000; //  890 : 192 - 0xc0
      12'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      12'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b00000001; //  903 :   1 - 0x1
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b00000010; //  912 :   2 - 0x2 -- Sprite 0x39
      12'h391: dout <= 8'b00000001; //  913 :   1 - 0x1
      12'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b00000001; //  920 :   1 - 0x1 -- plane 1
      12'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b10000000; //  944 : 128 - 0x80 -- Sprite 0x3b
      12'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000001; //  963 :   1 - 0x1
      12'h3C4: dout <= 8'b00100001; //  964 :  33 - 0x21
      12'h3C5: dout <= 8'b00010000; //  965 :  16 - 0x10
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000001; //  969 :   1 - 0x1
      12'h3CA: dout <= 8'b00000001; //  970 :   1 - 0x1
      12'h3CB: dout <= 8'b01000000; //  971 :  64 - 0x40
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b01100000; //  976 :  96 - 0x60 -- Sprite 0x3d
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00010000; //  979 :  16 - 0x10
      12'h3D4: dout <= 8'b00100001; //  980 :  33 - 0x21
      12'h3D5: dout <= 8'b00000001; //  981 :   1 - 0x1
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b10000000; //  984 : 128 - 0x80 -- plane 1
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b01000000; //  989 :  64 - 0x40
      12'h3DE: dout <= 8'b00000001; //  990 :   1 - 0x1
      12'h3DF: dout <= 8'b00000001; //  991 :   1 - 0x1
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      12'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout <= 8'b00001000; //  996 :   8 - 0x8
      12'h3E5: dout <= 8'b00010000; //  997 :  16 - 0x10
      12'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout <= 8'b00000100; // 1003 :   4 - 0x4
      12'h3EC: dout <= 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout <= 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout <= 8'b00001100; // 1008 :  12 - 0xc -- Sprite 0x3f
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00010000; // 1011 :  16 - 0x10
      12'h3F4: dout <= 8'b00001000; // 1012 :   8 - 0x8
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b00000010; // 1016 :   2 - 0x2 -- plane 1
      12'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout <= 8'b00000100; // 1021 :   4 - 0x4
      12'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b00000100; // 1024 :   4 - 0x4 -- Sprite 0x40
      12'h401: dout <= 8'b00000010; // 1025 :   2 - 0x2
      12'h402: dout <= 8'b00000001; // 1026 :   1 - 0x1
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout <= 8'b00001111; // 1032 :  15 - 0xf -- plane 1
      12'h409: dout <= 8'b00000111; // 1033 :   7 - 0x7
      12'h40A: dout <= 8'b00000011; // 1034 :   3 - 0x3
      12'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000001; // 1037 :   1 - 0x1
      12'h40E: dout <= 8'b00000001; // 1038 :   1 - 0x1
      12'h40F: dout <= 8'b00000001; // 1039 :   1 - 0x1
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      12'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      12'h415: dout <= 8'b00000000; // 1045 :   0 - 0x0
      12'h416: dout <= 8'b00000001; // 1046 :   1 - 0x1
      12'h417: dout <= 8'b00000011; // 1047 :   3 - 0x3
      12'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000001; // 1054 :   1 - 0x1
      12'h41F: dout <= 8'b00000011; // 1055 :   3 - 0x3
      12'h420: dout <= 8'b00000111; // 1056 :   7 - 0x7 -- Sprite 0x42
      12'h421: dout <= 8'b00000111; // 1057 :   7 - 0x7
      12'h422: dout <= 8'b00000111; // 1058 :   7 - 0x7
      12'h423: dout <= 8'b00000011; // 1059 :   3 - 0x3
      12'h424: dout <= 8'b00000001; // 1060 :   1 - 0x1
      12'h425: dout <= 8'b00000000; // 1061 :   0 - 0x0
      12'h426: dout <= 8'b00000000; // 1062 :   0 - 0x0
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000111; // 1064 :   7 - 0x7 -- plane 1
      12'h429: dout <= 8'b00000111; // 1065 :   7 - 0x7
      12'h42A: dout <= 8'b00000111; // 1066 :   7 - 0x7
      12'h42B: dout <= 8'b00000111; // 1067 :   7 - 0x7
      12'h42C: dout <= 8'b00000011; // 1068 :   3 - 0x3
      12'h42D: dout <= 8'b00000001; // 1069 :   1 - 0x1
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- plane 1
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      12'h441: dout <= 8'b01000010; // 1089 :  66 - 0x42
      12'h442: dout <= 8'b00111001; // 1090 :  57 - 0x39
      12'h443: dout <= 8'b11111111; // 1091 : 255 - 0xff
      12'h444: dout <= 8'b11111111; // 1092 : 255 - 0xff
      12'h445: dout <= 8'b11111111; // 1093 : 255 - 0xff
      12'h446: dout <= 8'b11111111; // 1094 : 255 - 0xff
      12'h447: dout <= 8'b11111111; // 1095 : 255 - 0xff
      12'h448: dout <= 8'b11111111; // 1096 : 255 - 0xff -- plane 1
      12'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      12'h44A: dout <= 8'b11111111; // 1098 : 255 - 0xff
      12'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      12'h44C: dout <= 8'b11111111; // 1100 : 255 - 0xff
      12'h44D: dout <= 8'b11111111; // 1101 : 255 - 0xff
      12'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      12'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      12'h450: dout <= 8'b01111111; // 1104 : 127 - 0x7f -- Sprite 0x45
      12'h451: dout <= 8'b00111111; // 1105 :  63 - 0x3f
      12'h452: dout <= 8'b00011111; // 1106 :  31 - 0x1f
      12'h453: dout <= 8'b00001111; // 1107 :  15 - 0xf
      12'h454: dout <= 8'b00011111; // 1108 :  31 - 0x1f
      12'h455: dout <= 8'b11111111; // 1109 : 255 - 0xff
      12'h456: dout <= 8'b11111111; // 1110 : 255 - 0xff
      12'h457: dout <= 8'b11111111; // 1111 : 255 - 0xff
      12'h458: dout <= 8'b11111111; // 1112 : 255 - 0xff -- plane 1
      12'h459: dout <= 8'b01111111; // 1113 : 127 - 0x7f
      12'h45A: dout <= 8'b00111111; // 1114 :  63 - 0x3f
      12'h45B: dout <= 8'b00011111; // 1115 :  31 - 0x1f
      12'h45C: dout <= 8'b00011111; // 1116 :  31 - 0x1f
      12'h45D: dout <= 8'b11111111; // 1117 : 255 - 0xff
      12'h45E: dout <= 8'b11111111; // 1118 : 255 - 0xff
      12'h45F: dout <= 8'b11111111; // 1119 : 255 - 0xff
      12'h460: dout <= 8'b11111000; // 1120 : 248 - 0xf8 -- Sprite 0x46
      12'h461: dout <= 8'b11110111; // 1121 : 247 - 0xf7
      12'h462: dout <= 8'b11101111; // 1122 : 239 - 0xef
      12'h463: dout <= 8'b11111111; // 1123 : 255 - 0xff
      12'h464: dout <= 8'b11111111; // 1124 : 255 - 0xff
      12'h465: dout <= 8'b11111110; // 1125 : 254 - 0xfe
      12'h466: dout <= 8'b01111110; // 1126 : 126 - 0x7e
      12'h467: dout <= 8'b00111110; // 1127 :  62 - 0x3e
      12'h468: dout <= 8'b11111111; // 1128 : 255 - 0xff -- plane 1
      12'h469: dout <= 8'b11111111; // 1129 : 255 - 0xff
      12'h46A: dout <= 8'b11111111; // 1130 : 255 - 0xff
      12'h46B: dout <= 8'b11111111; // 1131 : 255 - 0xff
      12'h46C: dout <= 8'b11111111; // 1132 : 255 - 0xff
      12'h46D: dout <= 8'b11111111; // 1133 : 255 - 0xff
      12'h46E: dout <= 8'b11111111; // 1134 : 255 - 0xff
      12'h46F: dout <= 8'b01111111; // 1135 : 127 - 0x7f
      12'h470: dout <= 8'b00000111; // 1136 :   7 - 0x7 -- Sprite 0x47
      12'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      12'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout <= 8'b00000000; // 1140 :   0 - 0x0
      12'h475: dout <= 8'b00000000; // 1141 :   0 - 0x0
      12'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b00000111; // 1144 :   7 - 0x7 -- plane 1
      12'h479: dout <= 8'b00000011; // 1145 :   3 - 0x3
      12'h47A: dout <= 8'b00000011; // 1146 :   3 - 0x3
      12'h47B: dout <= 8'b00000001; // 1147 :   1 - 0x1
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b11000000; // 1155 : 192 - 0xc0
      12'h484: dout <= 8'b11100000; // 1156 : 224 - 0xe0
      12'h485: dout <= 8'b11110000; // 1157 : 240 - 0xf0
      12'h486: dout <= 8'b11011011; // 1158 : 219 - 0xdb
      12'h487: dout <= 8'b11110110; // 1159 : 246 - 0xf6
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b10000000; // 1161 : 128 - 0x80
      12'h48A: dout <= 8'b10000000; // 1162 : 128 - 0x80
      12'h48B: dout <= 8'b11000000; // 1163 : 192 - 0xc0
      12'h48C: dout <= 8'b11100000; // 1164 : 224 - 0xe0
      12'h48D: dout <= 8'b11110000; // 1165 : 240 - 0xf0
      12'h48E: dout <= 8'b11111111; // 1166 : 255 - 0xff
      12'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      12'h490: dout <= 8'b11001011; // 1168 : 203 - 0xcb -- Sprite 0x49
      12'h491: dout <= 8'b11100000; // 1169 : 224 - 0xe0
      12'h492: dout <= 8'b11000100; // 1170 : 196 - 0xc4
      12'h493: dout <= 8'b00000010; // 1171 :   2 - 0x2
      12'h494: dout <= 8'b11010001; // 1172 : 209 - 0xd1
      12'h495: dout <= 8'b11100001; // 1173 : 225 - 0xe1
      12'h496: dout <= 8'b11010001; // 1174 : 209 - 0xd1
      12'h497: dout <= 8'b10000011; // 1175 : 131 - 0x83
      12'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- plane 1
      12'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      12'h49A: dout <= 8'b11111111; // 1178 : 255 - 0xff
      12'h49B: dout <= 8'b11111111; // 1179 : 255 - 0xff
      12'h49C: dout <= 8'b11111111; // 1180 : 255 - 0xff
      12'h49D: dout <= 8'b11111111; // 1181 : 255 - 0xff
      12'h49E: dout <= 8'b11111111; // 1182 : 255 - 0xff
      12'h49F: dout <= 8'b11111111; // 1183 : 255 - 0xff
      12'h4A0: dout <= 8'b00001111; // 1184 :  15 - 0xf -- Sprite 0x4a
      12'h4A1: dout <= 8'b11111111; // 1185 : 255 - 0xff
      12'h4A2: dout <= 8'b11100000; // 1186 : 224 - 0xe0
      12'h4A3: dout <= 8'b10001111; // 1187 : 143 - 0x8f
      12'h4A4: dout <= 8'b01101110; // 1188 : 110 - 0x6e
      12'h4A5: dout <= 8'b01000100; // 1189 :  68 - 0x44
      12'h4A6: dout <= 8'b11101110; // 1190 : 238 - 0xee
      12'h4A7: dout <= 8'b01100000; // 1191 :  96 - 0x60
      12'h4A8: dout <= 8'b11111111; // 1192 : 255 - 0xff -- plane 1
      12'h4A9: dout <= 8'b11111111; // 1193 : 255 - 0xff
      12'h4AA: dout <= 8'b11111111; // 1194 : 255 - 0xff
      12'h4AB: dout <= 8'b11110000; // 1195 : 240 - 0xf0
      12'h4AC: dout <= 8'b10000000; // 1196 : 128 - 0x80
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout <= 8'b10011111; // 1199 : 159 - 0x9f
      12'h4B0: dout <= 8'b10000011; // 1200 : 131 - 0x83 -- Sprite 0x4b
      12'h4B1: dout <= 8'b11100000; // 1201 : 224 - 0xe0
      12'h4B2: dout <= 8'b11100100; // 1202 : 228 - 0xe4
      12'h4B3: dout <= 8'b11000110; // 1203 : 198 - 0xc6
      12'h4B4: dout <= 8'b01100001; // 1204 :  97 - 0x61
      12'h4B5: dout <= 8'b00110011; // 1205 :  51 - 0x33
      12'h4B6: dout <= 8'b00011111; // 1206 :  31 - 0x1f
      12'h4B7: dout <= 8'b00001111; // 1207 :  15 - 0xf
      12'h4B8: dout <= 8'b11111111; // 1208 : 255 - 0xff -- plane 1
      12'h4B9: dout <= 8'b11111111; // 1209 : 255 - 0xff
      12'h4BA: dout <= 8'b11111001; // 1210 : 249 - 0xf9
      12'h4BB: dout <= 8'b11111001; // 1211 : 249 - 0xf9
      12'h4BC: dout <= 8'b01111111; // 1212 : 127 - 0x7f
      12'h4BD: dout <= 8'b00111111; // 1213 :  63 - 0x3f
      12'h4BE: dout <= 8'b00011111; // 1214 :  31 - 0x1f
      12'h4BF: dout <= 8'b00001111; // 1215 :  15 - 0xf
      12'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x4c
      12'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout <= 8'b00000011; // 1219 :   3 - 0x3
      12'h4C4: dout <= 8'b00000111; // 1220 :   7 - 0x7
      12'h4C5: dout <= 8'b00001111; // 1221 :  15 - 0xf
      12'h4C6: dout <= 8'b01011011; // 1222 :  91 - 0x5b
      12'h4C7: dout <= 8'b10100111; // 1223 : 167 - 0xa7
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00000001; // 1225 :   1 - 0x1
      12'h4CA: dout <= 8'b00000001; // 1226 :   1 - 0x1
      12'h4CB: dout <= 8'b00000011; // 1227 :   3 - 0x3
      12'h4CC: dout <= 8'b00000111; // 1228 :   7 - 0x7
      12'h4CD: dout <= 8'b00001111; // 1229 :  15 - 0xf
      12'h4CE: dout <= 8'b11111111; // 1230 : 255 - 0xff
      12'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      12'h4D0: dout <= 8'b01110011; // 1232 : 115 - 0x73 -- Sprite 0x4d
      12'h4D1: dout <= 8'b00000111; // 1233 :   7 - 0x7
      12'h4D2: dout <= 8'b00100111; // 1234 :  39 - 0x27
      12'h4D3: dout <= 8'b01000000; // 1235 :  64 - 0x40
      12'h4D4: dout <= 8'b10001011; // 1236 : 139 - 0x8b
      12'h4D5: dout <= 8'b10000111; // 1237 : 135 - 0x87
      12'h4D6: dout <= 8'b10001011; // 1238 : 139 - 0x8b
      12'h4D7: dout <= 8'b11000001; // 1239 : 193 - 0xc1
      12'h4D8: dout <= 8'b11111111; // 1240 : 255 - 0xff -- plane 1
      12'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      12'h4DA: dout <= 8'b11111111; // 1242 : 255 - 0xff
      12'h4DB: dout <= 8'b11111111; // 1243 : 255 - 0xff
      12'h4DC: dout <= 8'b11111111; // 1244 : 255 - 0xff
      12'h4DD: dout <= 8'b11111111; // 1245 : 255 - 0xff
      12'h4DE: dout <= 8'b11111111; // 1246 : 255 - 0xff
      12'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      12'h4E0: dout <= 8'b11110000; // 1248 : 240 - 0xf0 -- Sprite 0x4e
      12'h4E1: dout <= 8'b11111111; // 1249 : 255 - 0xff
      12'h4E2: dout <= 8'b00001111; // 1250 :  15 - 0xf
      12'h4E3: dout <= 8'b11100001; // 1251 : 225 - 0xe1
      12'h4E4: dout <= 8'b11101100; // 1252 : 236 - 0xec
      12'h4E5: dout <= 8'b01000100; // 1253 :  68 - 0x44
      12'h4E6: dout <= 8'b11101110; // 1254 : 238 - 0xee
      12'h4E7: dout <= 8'b00001100; // 1255 :  12 - 0xc
      12'h4E8: dout <= 8'b11111111; // 1256 : 255 - 0xff -- plane 1
      12'h4E9: dout <= 8'b11111111; // 1257 : 255 - 0xff
      12'h4EA: dout <= 8'b11111111; // 1258 : 255 - 0xff
      12'h4EB: dout <= 8'b00011111; // 1259 :  31 - 0x1f
      12'h4EC: dout <= 8'b00000011; // 1260 :   3 - 0x3
      12'h4ED: dout <= 8'b00000001; // 1261 :   1 - 0x1
      12'h4EE: dout <= 8'b00000001; // 1262 :   1 - 0x1
      12'h4EF: dout <= 8'b11110011; // 1263 : 243 - 0xf3
      12'h4F0: dout <= 8'b10000000; // 1264 : 128 - 0x80 -- Sprite 0x4f
      12'h4F1: dout <= 8'b00001110; // 1265 :  14 - 0xe
      12'h4F2: dout <= 8'b01001110; // 1266 :  78 - 0x4e
      12'h4F3: dout <= 8'b11000110; // 1267 : 198 - 0xc6
      12'h4F4: dout <= 8'b00001100; // 1268 :  12 - 0xc
      12'h4F5: dout <= 8'b10011000; // 1269 : 152 - 0x98
      12'h4F6: dout <= 8'b11110000; // 1270 : 240 - 0xf0
      12'h4F7: dout <= 8'b11100000; // 1271 : 224 - 0xe0
      12'h4F8: dout <= 8'b11111111; // 1272 : 255 - 0xff -- plane 1
      12'h4F9: dout <= 8'b11111111; // 1273 : 255 - 0xff
      12'h4FA: dout <= 8'b00111111; // 1274 :  63 - 0x3f
      12'h4FB: dout <= 8'b00111111; // 1275 :  63 - 0x3f
      12'h4FC: dout <= 8'b11111100; // 1276 : 252 - 0xfc
      12'h4FD: dout <= 8'b11111000; // 1277 : 248 - 0xf8
      12'h4FE: dout <= 8'b11110000; // 1278 : 240 - 0xf0
      12'h4FF: dout <= 8'b11100000; // 1279 : 224 - 0xe0
      12'h500: dout <= 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0x50
      12'h501: dout <= 8'b01000010; // 1281 :  66 - 0x42
      12'h502: dout <= 8'b10011100; // 1282 : 156 - 0x9c
      12'h503: dout <= 8'b11111111; // 1283 : 255 - 0xff
      12'h504: dout <= 8'b11111111; // 1284 : 255 - 0xff
      12'h505: dout <= 8'b11111111; // 1285 : 255 - 0xff
      12'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      12'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      12'h508: dout <= 8'b11111111; // 1288 : 255 - 0xff -- plane 1
      12'h509: dout <= 8'b11111111; // 1289 : 255 - 0xff
      12'h50A: dout <= 8'b11111111; // 1290 : 255 - 0xff
      12'h50B: dout <= 8'b11111111; // 1291 : 255 - 0xff
      12'h50C: dout <= 8'b11111111; // 1292 : 255 - 0xff
      12'h50D: dout <= 8'b11111111; // 1293 : 255 - 0xff
      12'h50E: dout <= 8'b11111111; // 1294 : 255 - 0xff
      12'h50F: dout <= 8'b11111111; // 1295 : 255 - 0xff
      12'h510: dout <= 8'b11111110; // 1296 : 254 - 0xfe -- Sprite 0x51
      12'h511: dout <= 8'b11111100; // 1297 : 252 - 0xfc
      12'h512: dout <= 8'b11111000; // 1298 : 248 - 0xf8
      12'h513: dout <= 8'b11110000; // 1299 : 240 - 0xf0
      12'h514: dout <= 8'b11111000; // 1300 : 248 - 0xf8
      12'h515: dout <= 8'b11111111; // 1301 : 255 - 0xff
      12'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      12'h517: dout <= 8'b11111111; // 1303 : 255 - 0xff
      12'h518: dout <= 8'b11111111; // 1304 : 255 - 0xff -- plane 1
      12'h519: dout <= 8'b11111110; // 1305 : 254 - 0xfe
      12'h51A: dout <= 8'b11111100; // 1306 : 252 - 0xfc
      12'h51B: dout <= 8'b11111000; // 1307 : 248 - 0xf8
      12'h51C: dout <= 8'b11111000; // 1308 : 248 - 0xf8
      12'h51D: dout <= 8'b11111111; // 1309 : 255 - 0xff
      12'h51E: dout <= 8'b11111111; // 1310 : 255 - 0xff
      12'h51F: dout <= 8'b11111111; // 1311 : 255 - 0xff
      12'h520: dout <= 8'b00011111; // 1312 :  31 - 0x1f -- Sprite 0x52
      12'h521: dout <= 8'b11101111; // 1313 : 239 - 0xef
      12'h522: dout <= 8'b11110111; // 1314 : 247 - 0xf7
      12'h523: dout <= 8'b11111111; // 1315 : 255 - 0xff
      12'h524: dout <= 8'b11111111; // 1316 : 255 - 0xff
      12'h525: dout <= 8'b11111110; // 1317 : 254 - 0xfe
      12'h526: dout <= 8'b01111100; // 1318 : 124 - 0x7c
      12'h527: dout <= 8'b01110000; // 1319 : 112 - 0x70
      12'h528: dout <= 8'b11111111; // 1320 : 255 - 0xff -- plane 1
      12'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      12'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      12'h52B: dout <= 8'b11111111; // 1323 : 255 - 0xff
      12'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      12'h52D: dout <= 8'b11111111; // 1325 : 255 - 0xff
      12'h52E: dout <= 8'b11111110; // 1326 : 254 - 0xfe
      12'h52F: dout <= 8'b11111100; // 1327 : 252 - 0xfc
      12'h530: dout <= 8'b11100000; // 1328 : 224 - 0xe0 -- Sprite 0x53
      12'h531: dout <= 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout <= 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout <= 8'b00000000; // 1331 :   0 - 0x0
      12'h534: dout <= 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      12'h536: dout <= 8'b00000000; // 1334 :   0 - 0x0
      12'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout <= 8'b11100000; // 1336 : 224 - 0xe0 -- plane 1
      12'h539: dout <= 8'b10000000; // 1337 : 128 - 0x80
      12'h53A: dout <= 8'b10000000; // 1338 : 128 - 0x80
      12'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout <= 8'b00100000; // 1344 :  32 - 0x20 -- Sprite 0x54
      12'h541: dout <= 8'b01000000; // 1345 :  64 - 0x40
      12'h542: dout <= 8'b10000000; // 1346 : 128 - 0x80
      12'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout <= 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout <= 8'b11110000; // 1352 : 240 - 0xf0 -- plane 1
      12'h549: dout <= 8'b11100000; // 1353 : 224 - 0xe0
      12'h54A: dout <= 8'b11000000; // 1354 : 192 - 0xc0
      12'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout <= 8'b10000000; // 1357 : 128 - 0x80
      12'h54E: dout <= 8'b10000000; // 1358 : 128 - 0x80
      12'h54F: dout <= 8'b10000000; // 1359 : 128 - 0x80
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      12'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout <= 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout <= 8'b10000000; // 1366 : 128 - 0x80
      12'h557: dout <= 8'b11000000; // 1367 : 192 - 0xc0
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b10000000; // 1374 : 128 - 0x80
      12'h55F: dout <= 8'b11000000; // 1375 : 192 - 0xc0
      12'h560: dout <= 8'b11100000; // 1376 : 224 - 0xe0 -- Sprite 0x56
      12'h561: dout <= 8'b11100000; // 1377 : 224 - 0xe0
      12'h562: dout <= 8'b11100000; // 1378 : 224 - 0xe0
      12'h563: dout <= 8'b11000000; // 1379 : 192 - 0xc0
      12'h564: dout <= 8'b10000000; // 1380 : 128 - 0x80
      12'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b11100000; // 1384 : 224 - 0xe0 -- plane 1
      12'h569: dout <= 8'b11100000; // 1385 : 224 - 0xe0
      12'h56A: dout <= 8'b11100000; // 1386 : 224 - 0xe0
      12'h56B: dout <= 8'b11100000; // 1387 : 224 - 0xe0
      12'h56C: dout <= 8'b11000000; // 1388 : 192 - 0xc0
      12'h56D: dout <= 8'b10000000; // 1389 : 128 - 0x80
      12'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0x57
      12'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      12'h581: dout <= 8'b11111111; // 1409 : 255 - 0xff
      12'h582: dout <= 8'b11111111; // 1410 : 255 - 0xff
      12'h583: dout <= 8'b11111111; // 1411 : 255 - 0xff
      12'h584: dout <= 8'b11111111; // 1412 : 255 - 0xff
      12'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      12'h586: dout <= 8'b11111111; // 1414 : 255 - 0xff
      12'h587: dout <= 8'b11111111; // 1415 : 255 - 0xff
      12'h588: dout <= 8'b11111111; // 1416 : 255 - 0xff -- plane 1
      12'h589: dout <= 8'b11111111; // 1417 : 255 - 0xff
      12'h58A: dout <= 8'b11111111; // 1418 : 255 - 0xff
      12'h58B: dout <= 8'b11111111; // 1419 : 255 - 0xff
      12'h58C: dout <= 8'b11111111; // 1420 : 255 - 0xff
      12'h58D: dout <= 8'b11111111; // 1421 : 255 - 0xff
      12'h58E: dout <= 8'b11111111; // 1422 : 255 - 0xff
      12'h58F: dout <= 8'b11111111; // 1423 : 255 - 0xff
      12'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0x59
      12'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      12'h592: dout <= 8'b11111111; // 1426 : 255 - 0xff
      12'h593: dout <= 8'b11111111; // 1427 : 255 - 0xff
      12'h594: dout <= 8'b11111111; // 1428 : 255 - 0xff
      12'h595: dout <= 8'b11111111; // 1429 : 255 - 0xff
      12'h596: dout <= 8'b11111111; // 1430 : 255 - 0xff
      12'h597: dout <= 8'b11111111; // 1431 : 255 - 0xff
      12'h598: dout <= 8'b11111111; // 1432 : 255 - 0xff -- plane 1
      12'h599: dout <= 8'b11111111; // 1433 : 255 - 0xff
      12'h59A: dout <= 8'b11111111; // 1434 : 255 - 0xff
      12'h59B: dout <= 8'b11111111; // 1435 : 255 - 0xff
      12'h59C: dout <= 8'b11111111; // 1436 : 255 - 0xff
      12'h59D: dout <= 8'b11111111; // 1437 : 255 - 0xff
      12'h59E: dout <= 8'b11111111; // 1438 : 255 - 0xff
      12'h59F: dout <= 8'b11111111; // 1439 : 255 - 0xff
      12'h5A0: dout <= 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      12'h5A1: dout <= 8'b11111111; // 1441 : 255 - 0xff
      12'h5A2: dout <= 8'b11111111; // 1442 : 255 - 0xff
      12'h5A3: dout <= 8'b11111111; // 1443 : 255 - 0xff
      12'h5A4: dout <= 8'b11111111; // 1444 : 255 - 0xff
      12'h5A5: dout <= 8'b11111111; // 1445 : 255 - 0xff
      12'h5A6: dout <= 8'b11111111; // 1446 : 255 - 0xff
      12'h5A7: dout <= 8'b11111111; // 1447 : 255 - 0xff
      12'h5A8: dout <= 8'b11111111; // 1448 : 255 - 0xff -- plane 1
      12'h5A9: dout <= 8'b11111111; // 1449 : 255 - 0xff
      12'h5AA: dout <= 8'b11111111; // 1450 : 255 - 0xff
      12'h5AB: dout <= 8'b11111111; // 1451 : 255 - 0xff
      12'h5AC: dout <= 8'b11111111; // 1452 : 255 - 0xff
      12'h5AD: dout <= 8'b11111111; // 1453 : 255 - 0xff
      12'h5AE: dout <= 8'b11111111; // 1454 : 255 - 0xff
      12'h5AF: dout <= 8'b11111111; // 1455 : 255 - 0xff
      12'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0x5b
      12'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      12'h5B2: dout <= 8'b11111111; // 1458 : 255 - 0xff
      12'h5B3: dout <= 8'b11111111; // 1459 : 255 - 0xff
      12'h5B4: dout <= 8'b11111111; // 1460 : 255 - 0xff
      12'h5B5: dout <= 8'b11111111; // 1461 : 255 - 0xff
      12'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      12'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      12'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- plane 1
      12'h5B9: dout <= 8'b11111111; // 1465 : 255 - 0xff
      12'h5BA: dout <= 8'b11111111; // 1466 : 255 - 0xff
      12'h5BB: dout <= 8'b11111111; // 1467 : 255 - 0xff
      12'h5BC: dout <= 8'b11111111; // 1468 : 255 - 0xff
      12'h5BD: dout <= 8'b11111111; // 1469 : 255 - 0xff
      12'h5BE: dout <= 8'b11111111; // 1470 : 255 - 0xff
      12'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      12'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0x5c
      12'h5C1: dout <= 8'b11111111; // 1473 : 255 - 0xff
      12'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      12'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      12'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      12'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      12'h5C6: dout <= 8'b11111111; // 1478 : 255 - 0xff
      12'h5C7: dout <= 8'b11111111; // 1479 : 255 - 0xff
      12'h5C8: dout <= 8'b11111111; // 1480 : 255 - 0xff -- plane 1
      12'h5C9: dout <= 8'b11111111; // 1481 : 255 - 0xff
      12'h5CA: dout <= 8'b11111111; // 1482 : 255 - 0xff
      12'h5CB: dout <= 8'b11111111; // 1483 : 255 - 0xff
      12'h5CC: dout <= 8'b11111111; // 1484 : 255 - 0xff
      12'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      12'h5CE: dout <= 8'b11111111; // 1486 : 255 - 0xff
      12'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      12'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      12'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      12'h5D2: dout <= 8'b11111111; // 1490 : 255 - 0xff
      12'h5D3: dout <= 8'b11111111; // 1491 : 255 - 0xff
      12'h5D4: dout <= 8'b11111111; // 1492 : 255 - 0xff
      12'h5D5: dout <= 8'b11111111; // 1493 : 255 - 0xff
      12'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      12'h5D7: dout <= 8'b11111111; // 1495 : 255 - 0xff
      12'h5D8: dout <= 8'b11111111; // 1496 : 255 - 0xff -- plane 1
      12'h5D9: dout <= 8'b11111111; // 1497 : 255 - 0xff
      12'h5DA: dout <= 8'b11111111; // 1498 : 255 - 0xff
      12'h5DB: dout <= 8'b11111111; // 1499 : 255 - 0xff
      12'h5DC: dout <= 8'b11111111; // 1500 : 255 - 0xff
      12'h5DD: dout <= 8'b11111111; // 1501 : 255 - 0xff
      12'h5DE: dout <= 8'b11111111; // 1502 : 255 - 0xff
      12'h5DF: dout <= 8'b11111111; // 1503 : 255 - 0xff
      12'h5E0: dout <= 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0x5e
      12'h5E1: dout <= 8'b11111111; // 1505 : 255 - 0xff
      12'h5E2: dout <= 8'b11111111; // 1506 : 255 - 0xff
      12'h5E3: dout <= 8'b11111111; // 1507 : 255 - 0xff
      12'h5E4: dout <= 8'b11111111; // 1508 : 255 - 0xff
      12'h5E5: dout <= 8'b11111111; // 1509 : 255 - 0xff
      12'h5E6: dout <= 8'b11111111; // 1510 : 255 - 0xff
      12'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      12'h5E8: dout <= 8'b11111111; // 1512 : 255 - 0xff -- plane 1
      12'h5E9: dout <= 8'b11111111; // 1513 : 255 - 0xff
      12'h5EA: dout <= 8'b11111111; // 1514 : 255 - 0xff
      12'h5EB: dout <= 8'b11111111; // 1515 : 255 - 0xff
      12'h5EC: dout <= 8'b11111111; // 1516 : 255 - 0xff
      12'h5ED: dout <= 8'b11111111; // 1517 : 255 - 0xff
      12'h5EE: dout <= 8'b11111111; // 1518 : 255 - 0xff
      12'h5EF: dout <= 8'b11111111; // 1519 : 255 - 0xff
      12'h5F0: dout <= 8'b11111111; // 1520 : 255 - 0xff -- Sprite 0x5f
      12'h5F1: dout <= 8'b11111111; // 1521 : 255 - 0xff
      12'h5F2: dout <= 8'b11111111; // 1522 : 255 - 0xff
      12'h5F3: dout <= 8'b11111111; // 1523 : 255 - 0xff
      12'h5F4: dout <= 8'b11111111; // 1524 : 255 - 0xff
      12'h5F5: dout <= 8'b11111111; // 1525 : 255 - 0xff
      12'h5F6: dout <= 8'b11111111; // 1526 : 255 - 0xff
      12'h5F7: dout <= 8'b11111111; // 1527 : 255 - 0xff
      12'h5F8: dout <= 8'b11111111; // 1528 : 255 - 0xff -- plane 1
      12'h5F9: dout <= 8'b11111111; // 1529 : 255 - 0xff
      12'h5FA: dout <= 8'b11111111; // 1530 : 255 - 0xff
      12'h5FB: dout <= 8'b11111111; // 1531 : 255 - 0xff
      12'h5FC: dout <= 8'b11111111; // 1532 : 255 - 0xff
      12'h5FD: dout <= 8'b11111111; // 1533 : 255 - 0xff
      12'h5FE: dout <= 8'b11111111; // 1534 : 255 - 0xff
      12'h5FF: dout <= 8'b11111111; // 1535 : 255 - 0xff
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00011111; // 1538 :  31 - 0x1f
      12'h603: dout <= 8'b00111111; // 1539 :  63 - 0x3f
      12'h604: dout <= 8'b00111111; // 1540 :  63 - 0x3f
      12'h605: dout <= 8'b01111111; // 1541 : 127 - 0x7f
      12'h606: dout <= 8'b01111111; // 1542 : 127 - 0x7f
      12'h607: dout <= 8'b01111111; // 1543 : 127 - 0x7f
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout <= 8'b00001111; // 1545 :  15 - 0xf
      12'h60A: dout <= 8'b00101000; // 1546 :  40 - 0x28
      12'h60B: dout <= 8'b01011100; // 1547 :  92 - 0x5c
      12'h60C: dout <= 8'b00111111; // 1548 :  63 - 0x3f
      12'h60D: dout <= 8'b01111111; // 1549 : 127 - 0x7f
      12'h60E: dout <= 8'b01111111; // 1550 : 127 - 0x7f
      12'h60F: dout <= 8'b01111111; // 1551 : 127 - 0x7f
      12'h610: dout <= 8'b01111111; // 1552 : 127 - 0x7f -- Sprite 0x61
      12'h611: dout <= 8'b00111110; // 1553 :  62 - 0x3e
      12'h612: dout <= 8'b00011111; // 1554 :  31 - 0x1f
      12'h613: dout <= 8'b00011111; // 1555 :  31 - 0x1f
      12'h614: dout <= 8'b00001111; // 1556 :  15 - 0xf
      12'h615: dout <= 8'b00001111; // 1557 :  15 - 0xf
      12'h616: dout <= 8'b00001111; // 1558 :  15 - 0xf
      12'h617: dout <= 8'b00000111; // 1559 :   7 - 0x7
      12'h618: dout <= 8'b01111111; // 1560 : 127 - 0x7f -- plane 1
      12'h619: dout <= 8'b00111110; // 1561 :  62 - 0x3e
      12'h61A: dout <= 8'b00011111; // 1562 :  31 - 0x1f
      12'h61B: dout <= 8'b00011111; // 1563 :  31 - 0x1f
      12'h61C: dout <= 8'b00001000; // 1564 :   8 - 0x8
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0x62
      12'h621: dout <= 8'b01100000; // 1569 :  96 - 0x60
      12'h622: dout <= 8'b11110000; // 1570 : 240 - 0xf0
      12'h623: dout <= 8'b11111000; // 1571 : 248 - 0xf8
      12'h624: dout <= 8'b11111000; // 1572 : 248 - 0xf8
      12'h625: dout <= 8'b11111000; // 1573 : 248 - 0xf8
      12'h626: dout <= 8'b11111100; // 1574 : 252 - 0xfc
      12'h627: dout <= 8'b11111100; // 1575 : 252 - 0xfc
      12'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout <= 8'b10000000; // 1577 : 128 - 0x80
      12'h62A: dout <= 8'b01000000; // 1578 :  64 - 0x40
      12'h62B: dout <= 8'b11000100; // 1579 : 196 - 0xc4
      12'h62C: dout <= 8'b11110110; // 1580 : 246 - 0xf6
      12'h62D: dout <= 8'b11111110; // 1581 : 254 - 0xfe
      12'h62E: dout <= 8'b11111100; // 1582 : 252 - 0xfc
      12'h62F: dout <= 8'b11111100; // 1583 : 252 - 0xfc
      12'h630: dout <= 8'b11111000; // 1584 : 248 - 0xf8 -- Sprite 0x63
      12'h631: dout <= 8'b11110000; // 1585 : 240 - 0xf0
      12'h632: dout <= 8'b11110000; // 1586 : 240 - 0xf0
      12'h633: dout <= 8'b11100000; // 1587 : 224 - 0xe0
      12'h634: dout <= 8'b10000000; // 1588 : 128 - 0x80
      12'h635: dout <= 8'b10000000; // 1589 : 128 - 0x80
      12'h636: dout <= 8'b11000000; // 1590 : 192 - 0xc0
      12'h637: dout <= 8'b11000000; // 1591 : 192 - 0xc0
      12'h638: dout <= 8'b11111000; // 1592 : 248 - 0xf8 -- plane 1
      12'h639: dout <= 8'b11110000; // 1593 : 240 - 0xf0
      12'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout <= 8'b10000000; // 1596 : 128 - 0x80
      12'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      12'h641: dout <= 8'b00011111; // 1601 :  31 - 0x1f
      12'h642: dout <= 8'b00111111; // 1602 :  63 - 0x3f
      12'h643: dout <= 8'b01111111; // 1603 : 127 - 0x7f
      12'h644: dout <= 8'b11111111; // 1604 : 255 - 0xff
      12'h645: dout <= 8'b11111111; // 1605 : 255 - 0xff
      12'h646: dout <= 8'b00111110; // 1606 :  62 - 0x3e
      12'h647: dout <= 8'b00001111; // 1607 :  15 - 0xf
      12'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout <= 8'b00011100; // 1609 :  28 - 0x1c
      12'h64A: dout <= 8'b00111111; // 1610 :  63 - 0x3f
      12'h64B: dout <= 8'b01111111; // 1611 : 127 - 0x7f
      12'h64C: dout <= 8'b11111111; // 1612 : 255 - 0xff
      12'h64D: dout <= 8'b11111111; // 1613 : 255 - 0xff
      12'h64E: dout <= 8'b00111110; // 1614 :  62 - 0x3e
      12'h64F: dout <= 8'b01110000; // 1615 : 112 - 0x70
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00000001; // 1619 :   1 - 0x1
      12'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout <= 8'b00000000; // 1622 :   0 - 0x0
      12'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0x66
      12'h661: dout <= 8'b11100000; // 1633 : 224 - 0xe0
      12'h662: dout <= 8'b11110000; // 1634 : 240 - 0xf0
      12'h663: dout <= 8'b11111100; // 1635 : 252 - 0xfc
      12'h664: dout <= 8'b11111110; // 1636 : 254 - 0xfe
      12'h665: dout <= 8'b11111110; // 1637 : 254 - 0xfe
      12'h666: dout <= 8'b11111111; // 1638 : 255 - 0xff
      12'h667: dout <= 8'b11111100; // 1639 : 252 - 0xfc
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout <= 8'b01100000; // 1641 :  96 - 0x60
      12'h66A: dout <= 8'b11110000; // 1642 : 240 - 0xf0
      12'h66B: dout <= 8'b11111000; // 1643 : 248 - 0xf8
      12'h66C: dout <= 8'b11111100; // 1644 : 252 - 0xfc
      12'h66D: dout <= 8'b11111100; // 1645 : 252 - 0xfc
      12'h66E: dout <= 8'b11111100; // 1646 : 252 - 0xfc
      12'h66F: dout <= 8'b11111111; // 1647 : 255 - 0xff
      12'h670: dout <= 8'b01111100; // 1648 : 124 - 0x7c -- Sprite 0x67
      12'h671: dout <= 8'b11111100; // 1649 : 252 - 0xfc
      12'h672: dout <= 8'b11111000; // 1650 : 248 - 0xf8
      12'h673: dout <= 8'b11110000; // 1651 : 240 - 0xf0
      12'h674: dout <= 8'b11100000; // 1652 : 224 - 0xe0
      12'h675: dout <= 8'b00000000; // 1653 :   0 - 0x0
      12'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b01111100; // 1656 : 124 - 0x7c -- plane 1
      12'h679: dout <= 8'b11111100; // 1657 : 252 - 0xfc
      12'h67A: dout <= 8'b10001000; // 1658 : 136 - 0x88
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      12'h681: dout <= 8'b00000111; // 1665 :   7 - 0x7
      12'h682: dout <= 8'b00000111; // 1666 :   7 - 0x7
      12'h683: dout <= 8'b00001111; // 1667 :  15 - 0xf
      12'h684: dout <= 8'b00001111; // 1668 :  15 - 0xf
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00011111; // 1670 :  31 - 0x1f
      12'h687: dout <= 8'b00111111; // 1671 :  63 - 0x3f
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout <= 8'b00000111; // 1673 :   7 - 0x7
      12'h68A: dout <= 8'b00000011; // 1674 :   3 - 0x3
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000111; // 1677 :   7 - 0x7
      12'h68E: dout <= 8'b00000100; // 1678 :   4 - 0x4
      12'h68F: dout <= 8'b00000100; // 1679 :   4 - 0x4
      12'h690: dout <= 8'b01111111; // 1680 : 127 - 0x7f -- Sprite 0x69
      12'h691: dout <= 8'b01111111; // 1681 : 127 - 0x7f
      12'h692: dout <= 8'b00011111; // 1682 :  31 - 0x1f
      12'h693: dout <= 8'b00011111; // 1683 :  31 - 0x1f
      12'h694: dout <= 8'b00011111; // 1684 :  31 - 0x1f
      12'h695: dout <= 8'b00011110; // 1685 :  30 - 0x1e
      12'h696: dout <= 8'b00001111; // 1686 :  15 - 0xf
      12'h697: dout <= 8'b00011111; // 1687 :  31 - 0x1f
      12'h698: dout <= 8'b00001100; // 1688 :  12 - 0xc -- plane 1
      12'h699: dout <= 8'b10011110; // 1689 : 158 - 0x9e
      12'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      12'h69B: dout <= 8'b00011111; // 1691 :  31 - 0x1f
      12'h69C: dout <= 8'b00011111; // 1692 :  31 - 0x1f
      12'h69D: dout <= 8'b00011110; // 1693 :  30 - 0x1e
      12'h69E: dout <= 8'b00001111; // 1694 :  15 - 0xf
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      12'h6A1: dout <= 8'b11100000; // 1697 : 224 - 0xe0
      12'h6A2: dout <= 8'b11100000; // 1698 : 224 - 0xe0
      12'h6A3: dout <= 8'b11110000; // 1699 : 240 - 0xf0
      12'h6A4: dout <= 8'b11110000; // 1700 : 240 - 0xf0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b11111000; // 1702 : 248 - 0xf8
      12'h6A7: dout <= 8'b11111100; // 1703 : 252 - 0xfc
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout <= 8'b11100000; // 1705 : 224 - 0xe0
      12'h6AA: dout <= 8'b11000000; // 1706 : 192 - 0xc0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b11100000; // 1709 : 224 - 0xe0
      12'h6AE: dout <= 8'b00100000; // 1710 :  32 - 0x20
      12'h6AF: dout <= 8'b00100000; // 1711 :  32 - 0x20
      12'h6B0: dout <= 8'b11111110; // 1712 : 254 - 0xfe -- Sprite 0x6b
      12'h6B1: dout <= 8'b11111110; // 1713 : 254 - 0xfe
      12'h6B2: dout <= 8'b11111000; // 1714 : 248 - 0xf8
      12'h6B3: dout <= 8'b11111000; // 1715 : 248 - 0xf8
      12'h6B4: dout <= 8'b11111000; // 1716 : 248 - 0xf8
      12'h6B5: dout <= 8'b01111000; // 1717 : 120 - 0x78
      12'h6B6: dout <= 8'b11110000; // 1718 : 240 - 0xf0
      12'h6B7: dout <= 8'b11111000; // 1719 : 248 - 0xf8
      12'h6B8: dout <= 8'b00110000; // 1720 :  48 - 0x30 -- plane 1
      12'h6B9: dout <= 8'b01111001; // 1721 : 121 - 0x79
      12'h6BA: dout <= 8'b11111111; // 1722 : 255 - 0xff
      12'h6BB: dout <= 8'b11111000; // 1723 : 248 - 0xf8
      12'h6BC: dout <= 8'b11111000; // 1724 : 248 - 0xf8
      12'h6BD: dout <= 8'b01111000; // 1725 : 120 - 0x78
      12'h6BE: dout <= 8'b11110000; // 1726 : 240 - 0xf0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b00000011; // 1728 :   3 - 0x3 -- Sprite 0x6c
      12'h6C1: dout <= 8'b00000111; // 1729 :   7 - 0x7
      12'h6C2: dout <= 8'b00000101; // 1730 :   5 - 0x5
      12'h6C3: dout <= 8'b00001000; // 1731 :   8 - 0x8
      12'h6C4: dout <= 8'b00011011; // 1732 :  27 - 0x1b
      12'h6C5: dout <= 8'b00011001; // 1733 :  25 - 0x19
      12'h6C6: dout <= 8'b00000101; // 1734 :   5 - 0x5
      12'h6C7: dout <= 8'b00111111; // 1735 :  63 - 0x3f
      12'h6C8: dout <= 8'b00000011; // 1736 :   3 - 0x3 -- plane 1
      12'h6C9: dout <= 8'b00000111; // 1737 :   7 - 0x7
      12'h6CA: dout <= 8'b00000010; // 1738 :   2 - 0x2
      12'h6CB: dout <= 8'b00000111; // 1739 :   7 - 0x7
      12'h6CC: dout <= 8'b00000100; // 1740 :   4 - 0x4
      12'h6CD: dout <= 8'b01000110; // 1741 :  70 - 0x46
      12'h6CE: dout <= 8'b11100011; // 1742 : 227 - 0xe3
      12'h6CF: dout <= 8'b11000010; // 1743 : 194 - 0xc2
      12'h6D0: dout <= 8'b00111111; // 1744 :  63 - 0x3f -- Sprite 0x6d
      12'h6D1: dout <= 8'b00001111; // 1745 :  15 - 0xf
      12'h6D2: dout <= 8'b00000101; // 1746 :   5 - 0x5
      12'h6D3: dout <= 8'b00110111; // 1747 :  55 - 0x37
      12'h6D4: dout <= 8'b00111111; // 1748 :  63 - 0x3f
      12'h6D5: dout <= 8'b00111111; // 1749 :  63 - 0x3f
      12'h6D6: dout <= 8'b00111110; // 1750 :  62 - 0x3e
      12'h6D7: dout <= 8'b00011100; // 1751 :  28 - 0x1c
      12'h6D8: dout <= 8'b01000010; // 1752 :  66 - 0x42 -- plane 1
      12'h6D9: dout <= 8'b00000111; // 1753 :   7 - 0x7
      12'h6DA: dout <= 8'b00000111; // 1754 :   7 - 0x7
      12'h6DB: dout <= 8'b00000111; // 1755 :   7 - 0x7
      12'h6DC: dout <= 8'b00000111; // 1756 :   7 - 0x7
      12'h6DD: dout <= 8'b00000011; // 1757 :   3 - 0x3
      12'h6DE: dout <= 8'b00000010; // 1758 :   2 - 0x2
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b11100000; // 1760 : 224 - 0xe0 -- Sprite 0x6e
      12'h6E1: dout <= 8'b11110000; // 1761 : 240 - 0xf0
      12'h6E2: dout <= 8'b01010000; // 1762 :  80 - 0x50
      12'h6E3: dout <= 8'b00001000; // 1763 :   8 - 0x8
      12'h6E4: dout <= 8'b01101100; // 1764 : 108 - 0x6c
      12'h6E5: dout <= 8'b11001100; // 1765 : 204 - 0xcc
      12'h6E6: dout <= 8'b11010000; // 1766 : 208 - 0xd0
      12'h6E7: dout <= 8'b11111110; // 1767 : 254 - 0xfe
      12'h6E8: dout <= 8'b11100000; // 1768 : 224 - 0xe0 -- plane 1
      12'h6E9: dout <= 8'b11110000; // 1769 : 240 - 0xf0
      12'h6EA: dout <= 8'b10100000; // 1770 : 160 - 0xa0
      12'h6EB: dout <= 8'b11110000; // 1771 : 240 - 0xf0
      12'h6EC: dout <= 8'b10010000; // 1772 : 144 - 0x90
      12'h6ED: dout <= 8'b00110010; // 1773 :  50 - 0x32
      12'h6EE: dout <= 8'b11100011; // 1774 : 227 - 0xe3
      12'h6EF: dout <= 8'b00100001; // 1775 :  33 - 0x21
      12'h6F0: dout <= 8'b11111110; // 1776 : 254 - 0xfe -- Sprite 0x6f
      12'h6F1: dout <= 8'b11111000; // 1777 : 248 - 0xf8
      12'h6F2: dout <= 8'b11010000; // 1778 : 208 - 0xd0
      12'h6F3: dout <= 8'b11111011; // 1779 : 251 - 0xfb
      12'h6F4: dout <= 8'b11111111; // 1780 : 255 - 0xff
      12'h6F5: dout <= 8'b11111111; // 1781 : 255 - 0xff
      12'h6F6: dout <= 8'b00111110; // 1782 :  62 - 0x3e
      12'h6F7: dout <= 8'b00001100; // 1783 :  12 - 0xc
      12'h6F8: dout <= 8'b00100000; // 1784 :  32 - 0x20 -- plane 1
      12'h6F9: dout <= 8'b01110000; // 1785 : 112 - 0x70
      12'h6FA: dout <= 8'b11110000; // 1786 : 240 - 0xf0
      12'h6FB: dout <= 8'b11111000; // 1787 : 248 - 0xf8
      12'h6FC: dout <= 8'b11111000; // 1788 : 248 - 0xf8
      12'h6FD: dout <= 8'b11110000; // 1789 : 240 - 0xf0
      12'h6FE: dout <= 8'b00110000; // 1790 :  48 - 0x30
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      12'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout <= 8'b01111001; // 1794 : 121 - 0x79
      12'h703: dout <= 8'b11111001; // 1795 : 249 - 0xf9
      12'h704: dout <= 8'b11110011; // 1796 : 243 - 0xf3
      12'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout <= 8'b01111011; // 1798 : 123 - 0x7b
      12'h707: dout <= 8'b00111111; // 1799 :  63 - 0x3f
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout <= 8'b00000001; // 1801 :   1 - 0x1
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b00011110; // 1805 :  30 - 0x1e
      12'h70E: dout <= 8'b01111111; // 1806 : 127 - 0x7f
      12'h70F: dout <= 8'b00111110; // 1807 :  62 - 0x3e
      12'h710: dout <= 8'b00111111; // 1808 :  63 - 0x3f -- Sprite 0x71
      12'h711: dout <= 8'b00111111; // 1809 :  63 - 0x3f
      12'h712: dout <= 8'b01111011; // 1810 : 123 - 0x7b
      12'h713: dout <= 8'b01111111; // 1811 : 127 - 0x7f
      12'h714: dout <= 8'b11111011; // 1812 : 251 - 0xfb
      12'h715: dout <= 8'b11110001; // 1813 : 241 - 0xf1
      12'h716: dout <= 8'b01111001; // 1814 : 121 - 0x79
      12'h717: dout <= 8'b00111000; // 1815 :  56 - 0x38
      12'h718: dout <= 8'b00111100; // 1816 :  60 - 0x3c -- plane 1
      12'h719: dout <= 8'b00111110; // 1817 :  62 - 0x3e
      12'h71A: dout <= 8'b01111111; // 1818 : 127 - 0x7f
      12'h71B: dout <= 8'b01111110; // 1819 : 126 - 0x7e
      12'h71C: dout <= 8'b00011000; // 1820 :  24 - 0x18
      12'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0x72
      12'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout <= 8'b10000000; // 1826 : 128 - 0x80
      12'h723: dout <= 8'b10110000; // 1827 : 176 - 0xb0
      12'h724: dout <= 8'b10111000; // 1828 : 184 - 0xb8
      12'h725: dout <= 8'b11000110; // 1829 : 198 - 0xc6
      12'h726: dout <= 8'b10010011; // 1830 : 147 - 0x93
      12'h727: dout <= 8'b11110111; // 1831 : 247 - 0xf7
      12'h728: dout <= 8'b11000000; // 1832 : 192 - 0xc0 -- plane 1
      12'h729: dout <= 8'b11100000; // 1833 : 224 - 0xe0
      12'h72A: dout <= 8'b01000000; // 1834 :  64 - 0x40
      12'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout <= 8'b00111010; // 1837 :  58 - 0x3a
      12'h72E: dout <= 8'b11101111; // 1838 : 239 - 0xef
      12'h72F: dout <= 8'b01001011; // 1839 :  75 - 0x4b
      12'h730: dout <= 8'b11100011; // 1840 : 227 - 0xe3 -- Sprite 0x73
      12'h731: dout <= 8'b11110111; // 1841 : 247 - 0xf7
      12'h732: dout <= 8'b10010011; // 1842 : 147 - 0x93
      12'h733: dout <= 8'b11000110; // 1843 : 198 - 0xc6
      12'h734: dout <= 8'b10111000; // 1844 : 184 - 0xb8
      12'h735: dout <= 8'b10110000; // 1845 : 176 - 0xb0
      12'h736: dout <= 8'b10000000; // 1846 : 128 - 0x80
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b01011111; // 1848 :  95 - 0x5f -- plane 1
      12'h739: dout <= 8'b01001011; // 1849 :  75 - 0x4b
      12'h73A: dout <= 8'b11101111; // 1850 : 239 - 0xef
      12'h73B: dout <= 8'b00111010; // 1851 :  58 - 0x3a
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout <= 8'b01100000; // 1854 :  96 - 0x60
      12'h73F: dout <= 8'b11000000; // 1855 : 192 - 0xc0
      12'h740: dout <= 8'b00110000; // 1856 :  48 - 0x30 -- Sprite 0x74
      12'h741: dout <= 8'b01111100; // 1857 : 124 - 0x7c
      12'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      12'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout <= 8'b11011111; // 1860 : 223 - 0xdf
      12'h745: dout <= 8'b00001011; // 1861 :  11 - 0xb
      12'h746: dout <= 8'b00011111; // 1862 :  31 - 0x1f
      12'h747: dout <= 8'b01111111; // 1863 : 127 - 0x7f
      12'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout <= 8'b00001100; // 1865 :  12 - 0xc
      12'h74A: dout <= 8'b00001111; // 1866 :  15 - 0xf
      12'h74B: dout <= 8'b00011111; // 1867 :  31 - 0x1f
      12'h74C: dout <= 8'b00011111; // 1868 :  31 - 0x1f
      12'h74D: dout <= 8'b00001111; // 1869 :  15 - 0xf
      12'h74E: dout <= 8'b00001110; // 1870 :  14 - 0xe
      12'h74F: dout <= 8'b00000100; // 1871 :   4 - 0x4
      12'h750: dout <= 8'b01111111; // 1872 : 127 - 0x7f -- Sprite 0x75
      12'h751: dout <= 8'b00001011; // 1873 :  11 - 0xb
      12'h752: dout <= 8'b00110011; // 1874 :  51 - 0x33
      12'h753: dout <= 8'b00110110; // 1875 :  54 - 0x36
      12'h754: dout <= 8'b00010000; // 1876 :  16 - 0x10
      12'h755: dout <= 8'b00001010; // 1877 :  10 - 0xa
      12'h756: dout <= 8'b00001111; // 1878 :  15 - 0xf
      12'h757: dout <= 8'b00000111; // 1879 :   7 - 0x7
      12'h758: dout <= 8'b10000100; // 1880 : 132 - 0x84 -- plane 1
      12'h759: dout <= 8'b11000111; // 1881 : 199 - 0xc7
      12'h75A: dout <= 8'b01001100; // 1882 :  76 - 0x4c
      12'h75B: dout <= 8'b00001001; // 1883 :   9 - 0x9
      12'h75C: dout <= 8'b00001111; // 1884 :  15 - 0xf
      12'h75D: dout <= 8'b00000101; // 1885 :   5 - 0x5
      12'h75E: dout <= 8'b00001111; // 1886 :  15 - 0xf
      12'h75F: dout <= 8'b00000111; // 1887 :   7 - 0x7
      12'h760: dout <= 8'b00111000; // 1888 :  56 - 0x38 -- Sprite 0x76
      12'h761: dout <= 8'b01111100; // 1889 : 124 - 0x7c
      12'h762: dout <= 8'b11111100; // 1890 : 252 - 0xfc
      12'h763: dout <= 8'b11111100; // 1891 : 252 - 0xfc
      12'h764: dout <= 8'b11101100; // 1892 : 236 - 0xec
      12'h765: dout <= 8'b10100000; // 1893 : 160 - 0xa0
      12'h766: dout <= 8'b11110000; // 1894 : 240 - 0xf0
      12'h767: dout <= 8'b11111100; // 1895 : 252 - 0xfc
      12'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- plane 1
      12'h769: dout <= 8'b01000000; // 1897 :  64 - 0x40
      12'h76A: dout <= 8'b11000000; // 1898 : 192 - 0xc0
      12'h76B: dout <= 8'b11100000; // 1899 : 224 - 0xe0
      12'h76C: dout <= 8'b11100000; // 1900 : 224 - 0xe0
      12'h76D: dout <= 8'b11100000; // 1901 : 224 - 0xe0
      12'h76E: dout <= 8'b11100000; // 1902 : 224 - 0xe0
      12'h76F: dout <= 8'b01000010; // 1903 :  66 - 0x42
      12'h770: dout <= 8'b11111100; // 1904 : 252 - 0xfc -- Sprite 0x77
      12'h771: dout <= 8'b10100000; // 1905 : 160 - 0xa0
      12'h772: dout <= 8'b10011000; // 1906 : 152 - 0x98
      12'h773: dout <= 8'b11011000; // 1907 : 216 - 0xd8
      12'h774: dout <= 8'b00010000; // 1908 :  16 - 0x10
      12'h775: dout <= 8'b10100000; // 1909 : 160 - 0xa0
      12'h776: dout <= 8'b11100000; // 1910 : 224 - 0xe0
      12'h777: dout <= 8'b11000000; // 1911 : 192 - 0xc0
      12'h778: dout <= 8'b01000011; // 1912 :  67 - 0x43 -- plane 1
      12'h779: dout <= 8'b11000111; // 1913 : 199 - 0xc7
      12'h77A: dout <= 8'b01100010; // 1914 :  98 - 0x62
      12'h77B: dout <= 8'b00100000; // 1915 :  32 - 0x20
      12'h77C: dout <= 8'b11100000; // 1916 : 224 - 0xe0
      12'h77D: dout <= 8'b01000000; // 1917 :  64 - 0x40
      12'h77E: dout <= 8'b11100000; // 1918 : 224 - 0xe0
      12'h77F: dout <= 8'b11000000; // 1919 : 192 - 0xc0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      12'h781: dout <= 8'b00000001; // 1921 :   1 - 0x1
      12'h782: dout <= 8'b00001101; // 1922 :  13 - 0xd
      12'h783: dout <= 8'b00011101; // 1923 :  29 - 0x1d
      12'h784: dout <= 8'b01100011; // 1924 :  99 - 0x63
      12'h785: dout <= 8'b11001001; // 1925 : 201 - 0xc9
      12'h786: dout <= 8'b11101111; // 1926 : 239 - 0xef
      12'h787: dout <= 8'b11000111; // 1927 : 199 - 0xc7
      12'h788: dout <= 8'b00000011; // 1928 :   3 - 0x3 -- plane 1
      12'h789: dout <= 8'b00000100; // 1929 :   4 - 0x4
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b01011100; // 1932 :  92 - 0x5c
      12'h78D: dout <= 8'b11110111; // 1933 : 247 - 0xf7
      12'h78E: dout <= 8'b11010010; // 1934 : 210 - 0xd2
      12'h78F: dout <= 8'b11111010; // 1935 : 250 - 0xfa
      12'h790: dout <= 8'b11101111; // 1936 : 239 - 0xef -- Sprite 0x79
      12'h791: dout <= 8'b11001001; // 1937 : 201 - 0xc9
      12'h792: dout <= 8'b01100011; // 1938 :  99 - 0x63
      12'h793: dout <= 8'b00011101; // 1939 :  29 - 0x1d
      12'h794: dout <= 8'b00001101; // 1940 :  13 - 0xd
      12'h795: dout <= 8'b00000001; // 1941 :   1 - 0x1
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b11010010; // 1944 : 210 - 0xd2 -- plane 1
      12'h799: dout <= 8'b11110111; // 1945 : 247 - 0xf7
      12'h79A: dout <= 8'b01011100; // 1946 :  92 - 0x5c
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000010; // 1949 :   2 - 0x2
      12'h79E: dout <= 8'b00000111; // 1950 :   7 - 0x7
      12'h79F: dout <= 8'b00000011; // 1951 :   3 - 0x3
      12'h7A0: dout <= 8'b00011100; // 1952 :  28 - 0x1c -- Sprite 0x7a
      12'h7A1: dout <= 8'b10011110; // 1953 : 158 - 0x9e
      12'h7A2: dout <= 8'b10001111; // 1954 : 143 - 0x8f
      12'h7A3: dout <= 8'b11011111; // 1955 : 223 - 0xdf
      12'h7A4: dout <= 8'b11111110; // 1956 : 254 - 0xfe
      12'h7A5: dout <= 8'b11011110; // 1957 : 222 - 0xde
      12'h7A6: dout <= 8'b11111100; // 1958 : 252 - 0xfc
      12'h7A7: dout <= 8'b11111100; // 1959 : 252 - 0xfc
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- plane 1
      12'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00011000; // 1963 :  24 - 0x18
      12'h7AC: dout <= 8'b01111110; // 1964 : 126 - 0x7e
      12'h7AD: dout <= 8'b11111110; // 1965 : 254 - 0xfe
      12'h7AE: dout <= 8'b01111100; // 1966 : 124 - 0x7c
      12'h7AF: dout <= 8'b00111100; // 1967 :  60 - 0x3c
      12'h7B0: dout <= 8'b11111100; // 1968 : 252 - 0xfc -- Sprite 0x7b
      12'h7B1: dout <= 8'b11011110; // 1969 : 222 - 0xde
      12'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      12'h7B3: dout <= 8'b11001111; // 1971 : 207 - 0xcf
      12'h7B4: dout <= 8'b10011111; // 1972 : 159 - 0x9f
      12'h7B5: dout <= 8'b10011110; // 1973 : 158 - 0x9e
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b01111100; // 1976 : 124 - 0x7c -- plane 1
      12'h7B9: dout <= 8'b11111110; // 1977 : 254 - 0xfe
      12'h7BA: dout <= 8'b01111000; // 1978 : 120 - 0x78
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b10000000; // 1982 : 128 - 0x80
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      12'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout <= 8'b00011110; // 1988 :  30 - 0x1e
      12'h7C5: dout <= 8'b00111111; // 1989 :  63 - 0x3f
      12'h7C6: dout <= 8'b01111101; // 1990 : 125 - 0x7d
      12'h7C7: dout <= 8'b01111000; // 1991 : 120 - 0x78
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout <= 8'b00000001; // 1994 :   1 - 0x1
      12'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout <= 8'b00100000; // 1997 :  32 - 0x20
      12'h7CE: dout <= 8'b01111100; // 1998 : 124 - 0x7c
      12'h7CF: dout <= 8'b01111000; // 1999 : 120 - 0x78
      12'h7D0: dout <= 8'b01111100; // 2000 : 124 - 0x7c -- Sprite 0x7d
      12'h7D1: dout <= 8'b11111011; // 2001 : 251 - 0xfb
      12'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout <= 8'b01011111; // 2004 :  95 - 0x5f
      12'h7D5: dout <= 8'b00011111; // 2005 :  31 - 0x1f
      12'h7D6: dout <= 8'b00011111; // 2006 :  31 - 0x1f
      12'h7D7: dout <= 8'b00011111; // 2007 :  31 - 0x1f
      12'h7D8: dout <= 8'b01111100; // 2008 : 124 - 0x7c -- plane 1
      12'h7D9: dout <= 8'b11111110; // 2009 : 254 - 0xfe
      12'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout <= 8'b11111110; // 2011 : 254 - 0xfe
      12'h7DC: dout <= 8'b01111100; // 2012 : 124 - 0x7c
      12'h7DD: dout <= 8'b01100000; // 2013 :  96 - 0x60
      12'h7DE: dout <= 8'b11100000; // 2014 : 224 - 0xe0
      12'h7DF: dout <= 8'b11100001; // 2015 : 225 - 0xe1
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout <= 8'b10000000; // 2021 : 128 - 0x80
      12'h7E6: dout <= 8'b10000000; // 2022 : 128 - 0x80
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b01111100; // 2024 : 124 - 0x7c -- plane 1
      12'h7E9: dout <= 8'b10000010; // 2025 : 130 - 0x82
      12'h7EA: dout <= 8'b00000001; // 2026 :   1 - 0x1
      12'h7EB: dout <= 8'b10000010; // 2027 : 130 - 0x82
      12'h7EC: dout <= 8'b01111100; // 2028 : 124 - 0x7c
      12'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      12'h7F1: dout <= 8'b00100001; // 2033 :  33 - 0x21
      12'h7F2: dout <= 8'b10100010; // 2034 : 162 - 0xa2
      12'h7F3: dout <= 8'b10100011; // 2035 : 163 - 0xa3
      12'h7F4: dout <= 8'b10110011; // 2036 : 179 - 0xb3
      12'h7F5: dout <= 8'b10001111; // 2037 : 143 - 0x8f
      12'h7F6: dout <= 8'b00100111; // 2038 :  39 - 0x27
      12'h7F7: dout <= 8'b11111110; // 2039 : 254 - 0xfe
      12'h7F8: dout <= 8'b00010000; // 2040 :  16 - 0x10 -- plane 1
      12'h7F9: dout <= 8'b00011001; // 2041 :  25 - 0x19
      12'h7FA: dout <= 8'b01011010; // 2042 :  90 - 0x5a
      12'h7FB: dout <= 8'b11011111; // 2043 : 223 - 0xdf
      12'h7FC: dout <= 8'b01001111; // 2044 :  79 - 0x4f
      12'h7FD: dout <= 8'b01110011; // 2045 : 115 - 0x73
      12'h7FE: dout <= 8'b11011011; // 2046 : 219 - 0xdb
      12'h7FF: dout <= 8'b00000010; // 2047 :   2 - 0x2
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Sprite 0x80
      12'h801: dout <= 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout <= 8'b00000000; // 2050 :   0 - 0x0
      12'h803: dout <= 8'b00000000; // 2051 :   0 - 0x0
      12'h804: dout <= 8'b00000011; // 2052 :   3 - 0x3
      12'h805: dout <= 8'b00001111; // 2053 :  15 - 0xf
      12'h806: dout <= 8'b00011111; // 2054 :  31 - 0x1f
      12'h807: dout <= 8'b00011111; // 2055 :  31 - 0x1f
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- plane 1
      12'h809: dout <= 8'b00000000; // 2057 :   0 - 0x0
      12'h80A: dout <= 8'b00000000; // 2058 :   0 - 0x0
      12'h80B: dout <= 8'b00000011; // 2059 :   3 - 0x3
      12'h80C: dout <= 8'b00001100; // 2060 :  12 - 0xc
      12'h80D: dout <= 8'b00010000; // 2061 :  16 - 0x10
      12'h80E: dout <= 8'b00100010; // 2062 :  34 - 0x22
      12'h80F: dout <= 8'b00100000; // 2063 :  32 - 0x20
      12'h810: dout <= 8'b00011111; // 2064 :  31 - 0x1f -- Sprite 0x81
      12'h811: dout <= 8'b00011111; // 2065 :  31 - 0x1f
      12'h812: dout <= 8'b00001111; // 2066 :  15 - 0xf
      12'h813: dout <= 8'b00000011; // 2067 :   3 - 0x3
      12'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b00100001; // 2072 :  33 - 0x21 -- plane 1
      12'h819: dout <= 8'b00100011; // 2073 :  35 - 0x23
      12'h81A: dout <= 8'b00010000; // 2074 :  16 - 0x10
      12'h81B: dout <= 8'b00001100; // 2075 :  12 - 0xc
      12'h81C: dout <= 8'b00000011; // 2076 :   3 - 0x3
      12'h81D: dout <= 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b00000000; // 2080 :   0 - 0x0 -- Sprite 0x82
      12'h821: dout <= 8'b00000000; // 2081 :   0 - 0x0
      12'h822: dout <= 8'b00000000; // 2082 :   0 - 0x0
      12'h823: dout <= 8'b00000000; // 2083 :   0 - 0x0
      12'h824: dout <= 8'b11000000; // 2084 : 192 - 0xc0
      12'h825: dout <= 8'b11110000; // 2085 : 240 - 0xf0
      12'h826: dout <= 8'b11111000; // 2086 : 248 - 0xf8
      12'h827: dout <= 8'b11111000; // 2087 : 248 - 0xf8
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout <= 8'b11000000; // 2091 : 192 - 0xc0
      12'h82C: dout <= 8'b00110000; // 2092 :  48 - 0x30
      12'h82D: dout <= 8'b00001000; // 2093 :   8 - 0x8
      12'h82E: dout <= 8'b01100100; // 2094 : 100 - 0x64
      12'h82F: dout <= 8'b11000100; // 2095 : 196 - 0xc4
      12'h830: dout <= 8'b11111000; // 2096 : 248 - 0xf8 -- Sprite 0x83
      12'h831: dout <= 8'b11111000; // 2097 : 248 - 0xf8
      12'h832: dout <= 8'b11110000; // 2098 : 240 - 0xf0
      12'h833: dout <= 8'b11000000; // 2099 : 192 - 0xc0
      12'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b10000100; // 2104 : 132 - 0x84 -- plane 1
      12'h839: dout <= 8'b00000100; // 2105 :   4 - 0x4
      12'h83A: dout <= 8'b00001000; // 2106 :   8 - 0x8
      12'h83B: dout <= 8'b00110000; // 2107 :  48 - 0x30
      12'h83C: dout <= 8'b11000000; // 2108 : 192 - 0xc0
      12'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout <= 8'b00000000; // 2112 :   0 - 0x0 -- Sprite 0x84
      12'h841: dout <= 8'b00000000; // 2113 :   0 - 0x0
      12'h842: dout <= 8'b00000000; // 2114 :   0 - 0x0
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000011; // 2116 :   3 - 0x3
      12'h845: dout <= 8'b00001111; // 2117 :  15 - 0xf
      12'h846: dout <= 8'b00011111; // 2118 :  31 - 0x1f
      12'h847: dout <= 8'b00011111; // 2119 :  31 - 0x1f
      12'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0 -- plane 1
      12'h849: dout <= 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout <= 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout <= 8'b00000011; // 2123 :   3 - 0x3
      12'h84C: dout <= 8'b00001100; // 2124 :  12 - 0xc
      12'h84D: dout <= 8'b00010000; // 2125 :  16 - 0x10
      12'h84E: dout <= 8'b00100110; // 2126 :  38 - 0x26
      12'h84F: dout <= 8'b00100011; // 2127 :  35 - 0x23
      12'h850: dout <= 8'b00011111; // 2128 :  31 - 0x1f -- Sprite 0x85
      12'h851: dout <= 8'b00011111; // 2129 :  31 - 0x1f
      12'h852: dout <= 8'b00001111; // 2130 :  15 - 0xf
      12'h853: dout <= 8'b00000011; // 2131 :   3 - 0x3
      12'h854: dout <= 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b00100001; // 2136 :  33 - 0x21 -- plane 1
      12'h859: dout <= 8'b00100000; // 2137 :  32 - 0x20
      12'h85A: dout <= 8'b00010000; // 2138 :  16 - 0x10
      12'h85B: dout <= 8'b00001100; // 2139 :  12 - 0xc
      12'h85C: dout <= 8'b00000011; // 2140 :   3 - 0x3
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b00000000; // 2144 :   0 - 0x0 -- Sprite 0x86
      12'h861: dout <= 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout <= 8'b11000000; // 2148 : 192 - 0xc0
      12'h865: dout <= 8'b11110000; // 2149 : 240 - 0xf0
      12'h866: dout <= 8'b11111000; // 2150 : 248 - 0xf8
      12'h867: dout <= 8'b11111000; // 2151 : 248 - 0xf8
      12'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b11000000; // 2155 : 192 - 0xc0
      12'h86C: dout <= 8'b00110000; // 2156 :  48 - 0x30
      12'h86D: dout <= 8'b00001000; // 2157 :   8 - 0x8
      12'h86E: dout <= 8'b01000100; // 2158 :  68 - 0x44
      12'h86F: dout <= 8'b00000100; // 2159 :   4 - 0x4
      12'h870: dout <= 8'b11111000; // 2160 : 248 - 0xf8 -- Sprite 0x87
      12'h871: dout <= 8'b11111000; // 2161 : 248 - 0xf8
      12'h872: dout <= 8'b11110000; // 2162 : 240 - 0xf0
      12'h873: dout <= 8'b11000000; // 2163 : 192 - 0xc0
      12'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout <= 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout <= 8'b10000100; // 2168 : 132 - 0x84 -- plane 1
      12'h879: dout <= 8'b11000100; // 2169 : 196 - 0xc4
      12'h87A: dout <= 8'b00001000; // 2170 :   8 - 0x8
      12'h87B: dout <= 8'b00110000; // 2171 :  48 - 0x30
      12'h87C: dout <= 8'b11000000; // 2172 : 192 - 0xc0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout <= 8'b00000000; // 2176 :   0 - 0x0 -- Sprite 0x88
      12'h881: dout <= 8'b00000000; // 2177 :   0 - 0x0
      12'h882: dout <= 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout <= 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout <= 8'b00000011; // 2180 :   3 - 0x3
      12'h885: dout <= 8'b00001111; // 2181 :  15 - 0xf
      12'h886: dout <= 8'b00011111; // 2182 :  31 - 0x1f
      12'h887: dout <= 8'b00011111; // 2183 :  31 - 0x1f
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout <= 8'b00000000; // 2185 :   0 - 0x0
      12'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout <= 8'b00000011; // 2187 :   3 - 0x3
      12'h88C: dout <= 8'b00001100; // 2188 :  12 - 0xc
      12'h88D: dout <= 8'b00010000; // 2189 :  16 - 0x10
      12'h88E: dout <= 8'b00100000; // 2190 :  32 - 0x20
      12'h88F: dout <= 8'b00100001; // 2191 :  33 - 0x21
      12'h890: dout <= 8'b00011111; // 2192 :  31 - 0x1f -- Sprite 0x89
      12'h891: dout <= 8'b00011111; // 2193 :  31 - 0x1f
      12'h892: dout <= 8'b00001111; // 2194 :  15 - 0xf
      12'h893: dout <= 8'b00000011; // 2195 :   3 - 0x3
      12'h894: dout <= 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout <= 8'b00000000; // 2197 :   0 - 0x0
      12'h896: dout <= 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00100011; // 2200 :  35 - 0x23 -- plane 1
      12'h899: dout <= 8'b00100110; // 2201 :  38 - 0x26
      12'h89A: dout <= 8'b00010000; // 2202 :  16 - 0x10
      12'h89B: dout <= 8'b00001100; // 2203 :  12 - 0xc
      12'h89C: dout <= 8'b00000011; // 2204 :   3 - 0x3
      12'h89D: dout <= 8'b00000000; // 2205 :   0 - 0x0
      12'h89E: dout <= 8'b00000000; // 2206 :   0 - 0x0
      12'h89F: dout <= 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout <= 8'b00000000; // 2208 :   0 - 0x0 -- Sprite 0x8a
      12'h8A1: dout <= 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout <= 8'b00000000; // 2210 :   0 - 0x0
      12'h8A3: dout <= 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout <= 8'b11000000; // 2212 : 192 - 0xc0
      12'h8A5: dout <= 8'b11110000; // 2213 : 240 - 0xf0
      12'h8A6: dout <= 8'b11111000; // 2214 : 248 - 0xf8
      12'h8A7: dout <= 8'b11111000; // 2215 : 248 - 0xf8
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout <= 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout <= 8'b11000000; // 2219 : 192 - 0xc0
      12'h8AC: dout <= 8'b00110000; // 2220 :  48 - 0x30
      12'h8AD: dout <= 8'b00001000; // 2221 :   8 - 0x8
      12'h8AE: dout <= 8'b11000100; // 2222 : 196 - 0xc4
      12'h8AF: dout <= 8'b10000100; // 2223 : 132 - 0x84
      12'h8B0: dout <= 8'b11111000; // 2224 : 248 - 0xf8 -- Sprite 0x8b
      12'h8B1: dout <= 8'b11111000; // 2225 : 248 - 0xf8
      12'h8B2: dout <= 8'b11110000; // 2226 : 240 - 0xf0
      12'h8B3: dout <= 8'b11000000; // 2227 : 192 - 0xc0
      12'h8B4: dout <= 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout <= 8'b00000000; // 2229 :   0 - 0x0
      12'h8B6: dout <= 8'b00000000; // 2230 :   0 - 0x0
      12'h8B7: dout <= 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout <= 8'b00000100; // 2232 :   4 - 0x4 -- plane 1
      12'h8B9: dout <= 8'b01000100; // 2233 :  68 - 0x44
      12'h8BA: dout <= 8'b00001000; // 2234 :   8 - 0x8
      12'h8BB: dout <= 8'b00110000; // 2235 :  48 - 0x30
      12'h8BC: dout <= 8'b11000000; // 2236 : 192 - 0xc0
      12'h8BD: dout <= 8'b00000000; // 2237 :   0 - 0x0
      12'h8BE: dout <= 8'b00000000; // 2238 :   0 - 0x0
      12'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout <= 8'b00000000; // 2240 :   0 - 0x0 -- Sprite 0x8c
      12'h8C1: dout <= 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout <= 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00000011; // 2244 :   3 - 0x3
      12'h8C5: dout <= 8'b00001111; // 2245 :  15 - 0xf
      12'h8C6: dout <= 8'b00011111; // 2246 :  31 - 0x1f
      12'h8C7: dout <= 8'b00011111; // 2247 :  31 - 0x1f
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000011; // 2251 :   3 - 0x3
      12'h8CC: dout <= 8'b00001100; // 2252 :  12 - 0xc
      12'h8CD: dout <= 8'b00010000; // 2253 :  16 - 0x10
      12'h8CE: dout <= 8'b00100011; // 2254 :  35 - 0x23
      12'h8CF: dout <= 8'b00100001; // 2255 :  33 - 0x21
      12'h8D0: dout <= 8'b00011111; // 2256 :  31 - 0x1f -- Sprite 0x8d
      12'h8D1: dout <= 8'b00011111; // 2257 :  31 - 0x1f
      12'h8D2: dout <= 8'b00001111; // 2258 :  15 - 0xf
      12'h8D3: dout <= 8'b00000011; // 2259 :   3 - 0x3
      12'h8D4: dout <= 8'b00000000; // 2260 :   0 - 0x0
      12'h8D5: dout <= 8'b00000000; // 2261 :   0 - 0x0
      12'h8D6: dout <= 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout <= 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout <= 8'b00100000; // 2264 :  32 - 0x20 -- plane 1
      12'h8D9: dout <= 8'b00100010; // 2265 :  34 - 0x22
      12'h8DA: dout <= 8'b00010000; // 2266 :  16 - 0x10
      12'h8DB: dout <= 8'b00001100; // 2267 :  12 - 0xc
      12'h8DC: dout <= 8'b00000011; // 2268 :   3 - 0x3
      12'h8DD: dout <= 8'b00000000; // 2269 :   0 - 0x0
      12'h8DE: dout <= 8'b00000000; // 2270 :   0 - 0x0
      12'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout <= 8'b00000000; // 2272 :   0 - 0x0 -- Sprite 0x8e
      12'h8E1: dout <= 8'b00000000; // 2273 :   0 - 0x0
      12'h8E2: dout <= 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout <= 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout <= 8'b11000000; // 2276 : 192 - 0xc0
      12'h8E5: dout <= 8'b11110000; // 2277 : 240 - 0xf0
      12'h8E6: dout <= 8'b11111000; // 2278 : 248 - 0xf8
      12'h8E7: dout <= 8'b11111000; // 2279 : 248 - 0xf8
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- plane 1
      12'h8E9: dout <= 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout <= 8'b11000000; // 2283 : 192 - 0xc0
      12'h8EC: dout <= 8'b00110000; // 2284 :  48 - 0x30
      12'h8ED: dout <= 8'b00001000; // 2285 :   8 - 0x8
      12'h8EE: dout <= 8'b00000100; // 2286 :   4 - 0x4
      12'h8EF: dout <= 8'b10000100; // 2287 : 132 - 0x84
      12'h8F0: dout <= 8'b11111000; // 2288 : 248 - 0xf8 -- Sprite 0x8f
      12'h8F1: dout <= 8'b11111000; // 2289 : 248 - 0xf8
      12'h8F2: dout <= 8'b11110000; // 2290 : 240 - 0xf0
      12'h8F3: dout <= 8'b11000000; // 2291 : 192 - 0xc0
      12'h8F4: dout <= 8'b00000000; // 2292 :   0 - 0x0
      12'h8F5: dout <= 8'b00000000; // 2293 :   0 - 0x0
      12'h8F6: dout <= 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout <= 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout <= 8'b11000100; // 2296 : 196 - 0xc4 -- plane 1
      12'h8F9: dout <= 8'b01100100; // 2297 : 100 - 0x64
      12'h8FA: dout <= 8'b00001000; // 2298 :   8 - 0x8
      12'h8FB: dout <= 8'b00110000; // 2299 :  48 - 0x30
      12'h8FC: dout <= 8'b11000000; // 2300 : 192 - 0xc0
      12'h8FD: dout <= 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout <= 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00001111; // 2307 :  15 - 0xf
      12'h904: dout <= 8'b00110000; // 2308 :  48 - 0x30
      12'h905: dout <= 8'b01100000; // 2309 :  96 - 0x60
      12'h906: dout <= 8'b00111111; // 2310 :  63 - 0x3f
      12'h907: dout <= 8'b01111111; // 2311 : 127 - 0x7f
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout <= 8'b00101111; // 2316 :  47 - 0x2f
      12'h90D: dout <= 8'b00111111; // 2317 :  63 - 0x3f
      12'h90E: dout <= 8'b01100000; // 2318 :  96 - 0x60
      12'h90F: dout <= 8'b00100000; // 2319 :  32 - 0x20
      12'h910: dout <= 8'b01111111; // 2320 : 127 - 0x7f -- Sprite 0x91
      12'h911: dout <= 8'b00111111; // 2321 :  63 - 0x3f
      12'h912: dout <= 8'b01100000; // 2322 :  96 - 0x60
      12'h913: dout <= 8'b00110000; // 2323 :  48 - 0x30
      12'h914: dout <= 8'b00001111; // 2324 :  15 - 0xf
      12'h915: dout <= 8'b00000000; // 2325 :   0 - 0x0
      12'h916: dout <= 8'b00000000; // 2326 :   0 - 0x0
      12'h917: dout <= 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout <= 8'b00100000; // 2328 :  32 - 0x20 -- plane 1
      12'h919: dout <= 8'b01100000; // 2329 :  96 - 0x60
      12'h91A: dout <= 8'b00111111; // 2330 :  63 - 0x3f
      12'h91B: dout <= 8'b00101111; // 2331 :  47 - 0x2f
      12'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b00000000; // 2336 :   0 - 0x0 -- Sprite 0x92
      12'h921: dout <= 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout <= 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout <= 8'b11111000; // 2339 : 248 - 0xf8
      12'h924: dout <= 8'b00000110; // 2340 :   6 - 0x6
      12'h925: dout <= 8'b00000011; // 2341 :   3 - 0x3
      12'h926: dout <= 8'b11111110; // 2342 : 254 - 0xfe
      12'h927: dout <= 8'b11111111; // 2343 : 255 - 0xff
      12'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0 -- plane 1
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00000000; // 2346 :   0 - 0x0
      12'h92B: dout <= 8'b00000000; // 2347 :   0 - 0x0
      12'h92C: dout <= 8'b11111010; // 2348 : 250 - 0xfa
      12'h92D: dout <= 8'b11111110; // 2349 : 254 - 0xfe
      12'h92E: dout <= 8'b00000011; // 2350 :   3 - 0x3
      12'h92F: dout <= 8'b00000010; // 2351 :   2 - 0x2
      12'h930: dout <= 8'b11111111; // 2352 : 255 - 0xff -- Sprite 0x93
      12'h931: dout <= 8'b11111110; // 2353 : 254 - 0xfe
      12'h932: dout <= 8'b00000011; // 2354 :   3 - 0x3
      12'h933: dout <= 8'b00000110; // 2355 :   6 - 0x6
      12'h934: dout <= 8'b11111000; // 2356 : 248 - 0xf8
      12'h935: dout <= 8'b00000000; // 2357 :   0 - 0x0
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000010; // 2360 :   2 - 0x2 -- plane 1
      12'h939: dout <= 8'b00000011; // 2361 :   3 - 0x3
      12'h93A: dout <= 8'b11111110; // 2362 : 254 - 0xfe
      12'h93B: dout <= 8'b11111010; // 2363 : 250 - 0xfa
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout <= 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout <= 8'b00101111; // 2372 :  47 - 0x2f
      12'h945: dout <= 8'b00111111; // 2373 :  63 - 0x3f
      12'h946: dout <= 8'b01100000; // 2374 :  96 - 0x60
      12'h947: dout <= 8'b00100000; // 2375 :  32 - 0x20
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- plane 1
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout <= 8'b00001111; // 2379 :  15 - 0xf
      12'h94C: dout <= 8'b00110000; // 2380 :  48 - 0x30
      12'h94D: dout <= 8'b01100000; // 2381 :  96 - 0x60
      12'h94E: dout <= 8'b00111111; // 2382 :  63 - 0x3f
      12'h94F: dout <= 8'b01111111; // 2383 : 127 - 0x7f
      12'h950: dout <= 8'b00100000; // 2384 :  32 - 0x20 -- Sprite 0x95
      12'h951: dout <= 8'b01100000; // 2385 :  96 - 0x60
      12'h952: dout <= 8'b00111111; // 2386 :  63 - 0x3f
      12'h953: dout <= 8'b00101111; // 2387 :  47 - 0x2f
      12'h954: dout <= 8'b00000000; // 2388 :   0 - 0x0
      12'h955: dout <= 8'b00000000; // 2389 :   0 - 0x0
      12'h956: dout <= 8'b00000000; // 2390 :   0 - 0x0
      12'h957: dout <= 8'b00000000; // 2391 :   0 - 0x0
      12'h958: dout <= 8'b01111111; // 2392 : 127 - 0x7f -- plane 1
      12'h959: dout <= 8'b00111111; // 2393 :  63 - 0x3f
      12'h95A: dout <= 8'b01100000; // 2394 :  96 - 0x60
      12'h95B: dout <= 8'b00110000; // 2395 :  48 - 0x30
      12'h95C: dout <= 8'b00001111; // 2396 :  15 - 0xf
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Sprite 0x96
      12'h961: dout <= 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout <= 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout <= 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout <= 8'b11111010; // 2404 : 250 - 0xfa
      12'h965: dout <= 8'b11111110; // 2405 : 254 - 0xfe
      12'h966: dout <= 8'b00000011; // 2406 :   3 - 0x3
      12'h967: dout <= 8'b00000010; // 2407 :   2 - 0x2
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- plane 1
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b00000000; // 2410 :   0 - 0x0
      12'h96B: dout <= 8'b11111000; // 2411 : 248 - 0xf8
      12'h96C: dout <= 8'b00000110; // 2412 :   6 - 0x6
      12'h96D: dout <= 8'b00000011; // 2413 :   3 - 0x3
      12'h96E: dout <= 8'b11111110; // 2414 : 254 - 0xfe
      12'h96F: dout <= 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout <= 8'b00000010; // 2416 :   2 - 0x2 -- Sprite 0x97
      12'h971: dout <= 8'b00000011; // 2417 :   3 - 0x3
      12'h972: dout <= 8'b11111110; // 2418 : 254 - 0xfe
      12'h973: dout <= 8'b11111010; // 2419 : 250 - 0xfa
      12'h974: dout <= 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b11111111; // 2424 : 255 - 0xff -- plane 1
      12'h979: dout <= 8'b11111110; // 2425 : 254 - 0xfe
      12'h97A: dout <= 8'b00000011; // 2426 :   3 - 0x3
      12'h97B: dout <= 8'b00000110; // 2427 :   6 - 0x6
      12'h97C: dout <= 8'b11111000; // 2428 : 248 - 0xf8
      12'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b00000000; // 2432 :   0 - 0x0 -- Sprite 0x98
      12'h981: dout <= 8'b01000100; // 2433 :  68 - 0x44
      12'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout <= 8'b01000001; // 2435 :  65 - 0x41
      12'h984: dout <= 8'b00100000; // 2436 :  32 - 0x20
      12'h985: dout <= 8'b01001011; // 2437 :  75 - 0x4b
      12'h986: dout <= 8'b00100111; // 2438 :  39 - 0x27
      12'h987: dout <= 8'b00011111; // 2439 :  31 - 0x1f
      12'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0 -- plane 1
      12'h989: dout <= 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout <= 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout <= 8'b01000000; // 2443 :  64 - 0x40
      12'h98C: dout <= 8'b00100000; // 2444 :  32 - 0x20
      12'h98D: dout <= 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout <= 8'b00000000; // 2446 :   0 - 0x0
      12'h98F: dout <= 8'b00000001; // 2447 :   1 - 0x1
      12'h990: dout <= 8'b00001111; // 2448 :  15 - 0xf -- Sprite 0x99
      12'h991: dout <= 8'b00011110; // 2449 :  30 - 0x1e
      12'h992: dout <= 8'b00011111; // 2450 :  31 - 0x1f
      12'h993: dout <= 8'b00011111; // 2451 :  31 - 0x1f
      12'h994: dout <= 8'b00011111; // 2452 :  31 - 0x1f
      12'h995: dout <= 8'b00001111; // 2453 :  15 - 0xf
      12'h996: dout <= 8'b00001111; // 2454 :  15 - 0xf
      12'h997: dout <= 8'b00000011; // 2455 :   3 - 0x3
      12'h998: dout <= 8'b00000011; // 2456 :   3 - 0x3 -- plane 1
      12'h999: dout <= 8'b00000111; // 2457 :   7 - 0x7
      12'h99A: dout <= 8'b00000110; // 2458 :   6 - 0x6
      12'h99B: dout <= 8'b00000110; // 2459 :   6 - 0x6
      12'h99C: dout <= 8'b00000111; // 2460 :   7 - 0x7
      12'h99D: dout <= 8'b00000011; // 2461 :   3 - 0x3
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b00000000; // 2464 :   0 - 0x0 -- Sprite 0x9a
      12'h9A1: dout <= 8'b00100000; // 2465 :  32 - 0x20
      12'h9A2: dout <= 8'b01010000; // 2466 :  80 - 0x50
      12'h9A3: dout <= 8'b00100000; // 2467 :  32 - 0x20
      12'h9A4: dout <= 8'b01100000; // 2468 :  96 - 0x60
      12'h9A5: dout <= 8'b01001000; // 2469 :  72 - 0x48
      12'h9A6: dout <= 8'b11100000; // 2470 : 224 - 0xe0
      12'h9A7: dout <= 8'b11110000; // 2471 : 240 - 0xf0
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b01000000; // 2474 :  64 - 0x40
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b00001000; // 2477 :   8 - 0x8
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b01000000; // 2479 :  64 - 0x40
      12'h9B0: dout <= 8'b11111000; // 2480 : 248 - 0xf8 -- Sprite 0x9b
      12'h9B1: dout <= 8'b01111000; // 2481 : 120 - 0x78
      12'h9B2: dout <= 8'b00111100; // 2482 :  60 - 0x3c
      12'h9B3: dout <= 8'b00111100; // 2483 :  60 - 0x3c
      12'h9B4: dout <= 8'b00111100; // 2484 :  60 - 0x3c
      12'h9B5: dout <= 8'b11111100; // 2485 : 252 - 0xfc
      12'h9B6: dout <= 8'b11111000; // 2486 : 248 - 0xf8
      12'h9B7: dout <= 8'b11100000; // 2487 : 224 - 0xe0
      12'h9B8: dout <= 8'b11100000; // 2488 : 224 - 0xe0 -- plane 1
      12'h9B9: dout <= 8'b11110000; // 2489 : 240 - 0xf0
      12'h9BA: dout <= 8'b11010000; // 2490 : 208 - 0xd0
      12'h9BB: dout <= 8'b11010000; // 2491 : 208 - 0xd0
      12'h9BC: dout <= 8'b11110000; // 2492 : 240 - 0xf0
      12'h9BD: dout <= 8'b11100000; // 2493 : 224 - 0xe0
      12'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00010000; // 2496 :  16 - 0x10 -- Sprite 0x9c
      12'h9C1: dout <= 8'b00000001; // 2497 :   1 - 0x1
      12'h9C2: dout <= 8'b00101010; // 2498 :  42 - 0x2a
      12'h9C3: dout <= 8'b00001100; // 2499 :  12 - 0xc
      12'h9C4: dout <= 8'b10100110; // 2500 : 166 - 0xa6
      12'h9C5: dout <= 8'b00010111; // 2501 :  23 - 0x17
      12'h9C6: dout <= 8'b00011111; // 2502 :  31 - 0x1f
      12'h9C7: dout <= 8'b00011111; // 2503 :  31 - 0x1f
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000010; // 2506 :   2 - 0x2
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b10000000; // 2508 : 128 - 0x80
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000011; // 2510 :   3 - 0x3
      12'h9CF: dout <= 8'b00000111; // 2511 :   7 - 0x7
      12'h9D0: dout <= 8'b01011110; // 2512 :  94 - 0x5e -- Sprite 0x9d
      12'h9D1: dout <= 8'b00111100; // 2513 :  60 - 0x3c
      12'h9D2: dout <= 8'b00111101; // 2514 :  61 - 0x3d
      12'h9D3: dout <= 8'b00111101; // 2515 :  61 - 0x3d
      12'h9D4: dout <= 8'b00111110; // 2516 :  62 - 0x3e
      12'h9D5: dout <= 8'b00011111; // 2517 :  31 - 0x1f
      12'h9D6: dout <= 8'b00001111; // 2518 :  15 - 0xf
      12'h9D7: dout <= 8'b00000111; // 2519 :   7 - 0x7
      12'h9D8: dout <= 8'b00000111; // 2520 :   7 - 0x7 -- plane 1
      12'h9D9: dout <= 8'b00001111; // 2521 :  15 - 0xf
      12'h9DA: dout <= 8'b00001110; // 2522 :  14 - 0xe
      12'h9DB: dout <= 8'b00001110; // 2523 :  14 - 0xe
      12'h9DC: dout <= 8'b00001111; // 2524 :  15 - 0xf
      12'h9DD: dout <= 8'b00000111; // 2525 :   7 - 0x7
      12'h9DE: dout <= 8'b00000011; // 2526 :   3 - 0x3
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Sprite 0x9e
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b10000000; // 2530 : 128 - 0x80
      12'h9E3: dout <= 8'b11001000; // 2531 : 200 - 0xc8
      12'h9E4: dout <= 8'b01100000; // 2532 :  96 - 0x60
      12'h9E5: dout <= 8'b11100000; // 2533 : 224 - 0xe0
      12'h9E6: dout <= 8'b11110100; // 2534 : 244 - 0xf4
      12'h9E7: dout <= 8'b11111000; // 2535 : 248 - 0xf8
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00001000; // 2539 :   8 - 0x8
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b10000000; // 2541 : 128 - 0x80
      12'h9EE: dout <= 8'b00100100; // 2542 :  36 - 0x24
      12'h9EF: dout <= 8'b11000000; // 2543 : 192 - 0xc0
      12'h9F0: dout <= 8'b01111100; // 2544 : 124 - 0x7c -- Sprite 0x9f
      12'h9F1: dout <= 8'b00011100; // 2545 :  28 - 0x1c
      12'h9F2: dout <= 8'b00101110; // 2546 :  46 - 0x2e
      12'h9F3: dout <= 8'b00101110; // 2547 :  46 - 0x2e
      12'h9F4: dout <= 8'b00011110; // 2548 :  30 - 0x1e
      12'h9F5: dout <= 8'b11111100; // 2549 : 252 - 0xfc
      12'h9F6: dout <= 8'b11111000; // 2550 : 248 - 0xf8
      12'h9F7: dout <= 8'b11100000; // 2551 : 224 - 0xe0
      12'h9F8: dout <= 8'b11110000; // 2552 : 240 - 0xf0 -- plane 1
      12'h9F9: dout <= 8'b11111000; // 2553 : 248 - 0xf8
      12'h9FA: dout <= 8'b11011000; // 2554 : 216 - 0xd8
      12'h9FB: dout <= 8'b11011000; // 2555 : 216 - 0xd8
      12'h9FC: dout <= 8'b11111000; // 2556 : 248 - 0xf8
      12'h9FD: dout <= 8'b11110000; // 2557 : 240 - 0xf0
      12'h9FE: dout <= 8'b11000000; // 2558 : 192 - 0xc0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b11111111; // 2560 : 255 - 0xff -- Sprite 0xa0
      12'hA01: dout <= 8'b11111111; // 2561 : 255 - 0xff
      12'hA02: dout <= 8'b00111000; // 2562 :  56 - 0x38
      12'hA03: dout <= 8'b01101100; // 2563 : 108 - 0x6c
      12'hA04: dout <= 8'b11000110; // 2564 : 198 - 0xc6
      12'hA05: dout <= 8'b10000011; // 2565 : 131 - 0x83
      12'hA06: dout <= 8'b11111111; // 2566 : 255 - 0xff
      12'hA07: dout <= 8'b11111111; // 2567 : 255 - 0xff
      12'hA08: dout <= 8'b11111111; // 2568 : 255 - 0xff -- plane 1
      12'hA09: dout <= 8'b11111111; // 2569 : 255 - 0xff
      12'hA0A: dout <= 8'b00111000; // 2570 :  56 - 0x38
      12'hA0B: dout <= 8'b01101100; // 2571 : 108 - 0x6c
      12'hA0C: dout <= 8'b11000110; // 2572 : 198 - 0xc6
      12'hA0D: dout <= 8'b10000011; // 2573 : 131 - 0x83
      12'hA0E: dout <= 8'b11111111; // 2574 : 255 - 0xff
      12'hA0F: dout <= 8'b11111111; // 2575 : 255 - 0xff
      12'hA10: dout <= 8'b11111111; // 2576 : 255 - 0xff -- Sprite 0xa1
      12'hA11: dout <= 8'b11111111; // 2577 : 255 - 0xff
      12'hA12: dout <= 8'b00111000; // 2578 :  56 - 0x38
      12'hA13: dout <= 8'b01101100; // 2579 : 108 - 0x6c
      12'hA14: dout <= 8'b11000110; // 2580 : 198 - 0xc6
      12'hA15: dout <= 8'b10000011; // 2581 : 131 - 0x83
      12'hA16: dout <= 8'b11111111; // 2582 : 255 - 0xff
      12'hA17: dout <= 8'b11111111; // 2583 : 255 - 0xff
      12'hA18: dout <= 8'b11111111; // 2584 : 255 - 0xff -- plane 1
      12'hA19: dout <= 8'b11111111; // 2585 : 255 - 0xff
      12'hA1A: dout <= 8'b00111000; // 2586 :  56 - 0x38
      12'hA1B: dout <= 8'b01101100; // 2587 : 108 - 0x6c
      12'hA1C: dout <= 8'b11000110; // 2588 : 198 - 0xc6
      12'hA1D: dout <= 8'b10000011; // 2589 : 131 - 0x83
      12'hA1E: dout <= 8'b11111111; // 2590 : 255 - 0xff
      12'hA1F: dout <= 8'b11111111; // 2591 : 255 - 0xff
      12'hA20: dout <= 8'b10010010; // 2592 : 146 - 0x92 -- Sprite 0xa2
      12'hA21: dout <= 8'b01010100; // 2593 :  84 - 0x54
      12'hA22: dout <= 8'b00111000; // 2594 :  56 - 0x38
      12'hA23: dout <= 8'b11111110; // 2595 : 254 - 0xfe
      12'hA24: dout <= 8'b00111000; // 2596 :  56 - 0x38
      12'hA25: dout <= 8'b01010100; // 2597 :  84 - 0x54
      12'hA26: dout <= 8'b10010010; // 2598 : 146 - 0x92
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b11111111; // 2608 : 255 - 0xff -- Sprite 0xa3
      12'hA31: dout <= 8'b11111111; // 2609 : 255 - 0xff
      12'hA32: dout <= 8'b11111111; // 2610 : 255 - 0xff
      12'hA33: dout <= 8'b11111111; // 2611 : 255 - 0xff
      12'hA34: dout <= 8'b11111111; // 2612 : 255 - 0xff
      12'hA35: dout <= 8'b11111111; // 2613 : 255 - 0xff
      12'hA36: dout <= 8'b11111111; // 2614 : 255 - 0xff
      12'hA37: dout <= 8'b11111111; // 2615 : 255 - 0xff
      12'hA38: dout <= 8'b11111111; // 2616 : 255 - 0xff -- plane 1
      12'hA39: dout <= 8'b11111111; // 2617 : 255 - 0xff
      12'hA3A: dout <= 8'b11111111; // 2618 : 255 - 0xff
      12'hA3B: dout <= 8'b11111111; // 2619 : 255 - 0xff
      12'hA3C: dout <= 8'b11111111; // 2620 : 255 - 0xff
      12'hA3D: dout <= 8'b11111111; // 2621 : 255 - 0xff
      12'hA3E: dout <= 8'b11111111; // 2622 : 255 - 0xff
      12'hA3F: dout <= 8'b11111111; // 2623 : 255 - 0xff
      12'hA40: dout <= 8'b11111111; // 2624 : 255 - 0xff -- Sprite 0xa4
      12'hA41: dout <= 8'b11111111; // 2625 : 255 - 0xff
      12'hA42: dout <= 8'b11111111; // 2626 : 255 - 0xff
      12'hA43: dout <= 8'b11111111; // 2627 : 255 - 0xff
      12'hA44: dout <= 8'b11111111; // 2628 : 255 - 0xff
      12'hA45: dout <= 8'b11111111; // 2629 : 255 - 0xff
      12'hA46: dout <= 8'b11111111; // 2630 : 255 - 0xff
      12'hA47: dout <= 8'b11111111; // 2631 : 255 - 0xff
      12'hA48: dout <= 8'b11111111; // 2632 : 255 - 0xff -- plane 1
      12'hA49: dout <= 8'b11111111; // 2633 : 255 - 0xff
      12'hA4A: dout <= 8'b11111111; // 2634 : 255 - 0xff
      12'hA4B: dout <= 8'b11111111; // 2635 : 255 - 0xff
      12'hA4C: dout <= 8'b11111111; // 2636 : 255 - 0xff
      12'hA4D: dout <= 8'b11111111; // 2637 : 255 - 0xff
      12'hA4E: dout <= 8'b11111111; // 2638 : 255 - 0xff
      12'hA4F: dout <= 8'b11111111; // 2639 : 255 - 0xff
      12'hA50: dout <= 8'b11111111; // 2640 : 255 - 0xff -- Sprite 0xa5
      12'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout <= 8'b11111111; // 2642 : 255 - 0xff
      12'hA53: dout <= 8'b11111111; // 2643 : 255 - 0xff
      12'hA54: dout <= 8'b11111111; // 2644 : 255 - 0xff
      12'hA55: dout <= 8'b11111111; // 2645 : 255 - 0xff
      12'hA56: dout <= 8'b11111111; // 2646 : 255 - 0xff
      12'hA57: dout <= 8'b11111111; // 2647 : 255 - 0xff
      12'hA58: dout <= 8'b11111111; // 2648 : 255 - 0xff -- plane 1
      12'hA59: dout <= 8'b11111111; // 2649 : 255 - 0xff
      12'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      12'hA5B: dout <= 8'b11111111; // 2651 : 255 - 0xff
      12'hA5C: dout <= 8'b11111111; // 2652 : 255 - 0xff
      12'hA5D: dout <= 8'b11111111; // 2653 : 255 - 0xff
      12'hA5E: dout <= 8'b11111111; // 2654 : 255 - 0xff
      12'hA5F: dout <= 8'b11111111; // 2655 : 255 - 0xff
      12'hA60: dout <= 8'b11111111; // 2656 : 255 - 0xff -- Sprite 0xa6
      12'hA61: dout <= 8'b11111111; // 2657 : 255 - 0xff
      12'hA62: dout <= 8'b11111111; // 2658 : 255 - 0xff
      12'hA63: dout <= 8'b11111111; // 2659 : 255 - 0xff
      12'hA64: dout <= 8'b11111111; // 2660 : 255 - 0xff
      12'hA65: dout <= 8'b11111111; // 2661 : 255 - 0xff
      12'hA66: dout <= 8'b11111111; // 2662 : 255 - 0xff
      12'hA67: dout <= 8'b11111111; // 2663 : 255 - 0xff
      12'hA68: dout <= 8'b11111111; // 2664 : 255 - 0xff -- plane 1
      12'hA69: dout <= 8'b11111111; // 2665 : 255 - 0xff
      12'hA6A: dout <= 8'b11111111; // 2666 : 255 - 0xff
      12'hA6B: dout <= 8'b11111111; // 2667 : 255 - 0xff
      12'hA6C: dout <= 8'b11111111; // 2668 : 255 - 0xff
      12'hA6D: dout <= 8'b11111111; // 2669 : 255 - 0xff
      12'hA6E: dout <= 8'b11111111; // 2670 : 255 - 0xff
      12'hA6F: dout <= 8'b11111111; // 2671 : 255 - 0xff
      12'hA70: dout <= 8'b11111111; // 2672 : 255 - 0xff -- Sprite 0xa7
      12'hA71: dout <= 8'b11111111; // 2673 : 255 - 0xff
      12'hA72: dout <= 8'b11111111; // 2674 : 255 - 0xff
      12'hA73: dout <= 8'b11111111; // 2675 : 255 - 0xff
      12'hA74: dout <= 8'b11111111; // 2676 : 255 - 0xff
      12'hA75: dout <= 8'b11111111; // 2677 : 255 - 0xff
      12'hA76: dout <= 8'b11111111; // 2678 : 255 - 0xff
      12'hA77: dout <= 8'b11111111; // 2679 : 255 - 0xff
      12'hA78: dout <= 8'b11111111; // 2680 : 255 - 0xff -- plane 1
      12'hA79: dout <= 8'b11111111; // 2681 : 255 - 0xff
      12'hA7A: dout <= 8'b11111111; // 2682 : 255 - 0xff
      12'hA7B: dout <= 8'b11111111; // 2683 : 255 - 0xff
      12'hA7C: dout <= 8'b11111111; // 2684 : 255 - 0xff
      12'hA7D: dout <= 8'b11111111; // 2685 : 255 - 0xff
      12'hA7E: dout <= 8'b11111111; // 2686 : 255 - 0xff
      12'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout <= 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout <= 8'b00100011; // 2693 :  35 - 0x23
      12'hA86: dout <= 8'b10010111; // 2694 : 151 - 0x97
      12'hA87: dout <= 8'b00101111; // 2695 :  47 - 0x2f
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- plane 1
      12'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout <= 8'b00000001; // 2702 :   1 - 0x1
      12'hA8F: dout <= 8'b00000011; // 2703 :   3 - 0x3
      12'hA90: dout <= 8'b01101110; // 2704 : 110 - 0x6e -- Sprite 0xa9
      12'hA91: dout <= 8'b11101111; // 2705 : 239 - 0xef
      12'hA92: dout <= 8'b11110111; // 2706 : 247 - 0xf7
      12'hA93: dout <= 8'b11111111; // 2707 : 255 - 0xff
      12'hA94: dout <= 8'b01111111; // 2708 : 127 - 0x7f
      12'hA95: dout <= 8'b00111111; // 2709 :  63 - 0x3f
      12'hA96: dout <= 8'b01011111; // 2710 :  95 - 0x5f
      12'hA97: dout <= 8'b00001111; // 2711 :  15 - 0xf
      12'hA98: dout <= 8'b00000111; // 2712 :   7 - 0x7 -- plane 1
      12'hA99: dout <= 8'b00000111; // 2713 :   7 - 0x7
      12'hA9A: dout <= 8'b00000011; // 2714 :   3 - 0x3
      12'hA9B: dout <= 8'b00100111; // 2715 :  39 - 0x27
      12'hA9C: dout <= 8'b00011111; // 2716 :  31 - 0x1f
      12'hA9D: dout <= 8'b00000111; // 2717 :   7 - 0x7
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b00000000; // 2720 :   0 - 0x0 -- Sprite 0xaa
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b11111000; // 2724 : 248 - 0xf8
      12'hAA5: dout <= 8'b11111100; // 2725 : 252 - 0xfc
      12'hAA6: dout <= 8'b11111110; // 2726 : 254 - 0xfe
      12'hAA7: dout <= 8'b01011110; // 2727 :  94 - 0x5e
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b11110000; // 2733 : 240 - 0xf0
      12'hAAE: dout <= 8'b11111000; // 2734 : 248 - 0xf8
      12'hAAF: dout <= 8'b10101100; // 2735 : 172 - 0xac
      12'hAB0: dout <= 8'b01011110; // 2736 :  94 - 0x5e -- Sprite 0xab
      12'hAB1: dout <= 8'b00001100; // 2737 :  12 - 0xc
      12'hAB2: dout <= 8'b10011110; // 2738 : 158 - 0x9e
      12'hAB3: dout <= 8'b11111110; // 2739 : 254 - 0xfe
      12'hAB4: dout <= 8'b11111110; // 2740 : 254 - 0xfe
      12'hAB5: dout <= 8'b11111110; // 2741 : 254 - 0xfe
      12'hAB6: dout <= 8'b11111000; // 2742 : 248 - 0xf8
      12'hAB7: dout <= 8'b11000000; // 2743 : 192 - 0xc0
      12'hAB8: dout <= 8'b10101100; // 2744 : 172 - 0xac -- plane 1
      12'hAB9: dout <= 8'b11111000; // 2745 : 248 - 0xf8
      12'hABA: dout <= 8'b11111000; // 2746 : 248 - 0xf8
      12'hABB: dout <= 8'b11111000; // 2747 : 248 - 0xf8
      12'hABC: dout <= 8'b11110000; // 2748 : 240 - 0xf0
      12'hABD: dout <= 8'b11000000; // 2749 : 192 - 0xc0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout <= 8'b00000011; // 2757 :   3 - 0x3
      12'hAC6: dout <= 8'b00000111; // 2758 :   7 - 0x7
      12'hAC7: dout <= 8'b00101111; // 2759 :  47 - 0x2f
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000001; // 2766 :   1 - 0x1
      12'hACF: dout <= 8'b00000011; // 2767 :   3 - 0x3
      12'hAD0: dout <= 8'b01001110; // 2768 :  78 - 0x4e -- Sprite 0xad
      12'hAD1: dout <= 8'b01101110; // 2769 : 110 - 0x6e
      12'hAD2: dout <= 8'b11111110; // 2770 : 254 - 0xfe
      12'hAD3: dout <= 8'b01111111; // 2771 : 127 - 0x7f
      12'hAD4: dout <= 8'b00111111; // 2772 :  63 - 0x3f
      12'hAD5: dout <= 8'b00011111; // 2773 :  31 - 0x1f
      12'hAD6: dout <= 8'b00001111; // 2774 :  15 - 0xf
      12'hAD7: dout <= 8'b00000011; // 2775 :   3 - 0x3
      12'hAD8: dout <= 8'b00000111; // 2776 :   7 - 0x7 -- plane 1
      12'hAD9: dout <= 8'b00000111; // 2777 :   7 - 0x7
      12'hADA: dout <= 8'b00000111; // 2778 :   7 - 0x7
      12'hADB: dout <= 8'b00100111; // 2779 :  39 - 0x27
      12'hADC: dout <= 8'b00011111; // 2780 :  31 - 0x1f
      12'hADD: dout <= 8'b00000111; // 2781 :   7 - 0x7
      12'hADE: dout <= 8'b00000001; // 2782 :   1 - 0x1
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Sprite 0xae
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00000000; // 2786 :   0 - 0x0
      12'hAE3: dout <= 8'b00000000; // 2787 :   0 - 0x0
      12'hAE4: dout <= 8'b11111000; // 2788 : 248 - 0xf8
      12'hAE5: dout <= 8'b11111100; // 2789 : 252 - 0xfc
      12'hAE6: dout <= 8'b11111110; // 2790 : 254 - 0xfe
      12'hAE7: dout <= 8'b01010110; // 2791 :  86 - 0x56
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b11110000; // 2797 : 240 - 0xf0
      12'hAEE: dout <= 8'b11111000; // 2798 : 248 - 0xf8
      12'hAEF: dout <= 8'b10101100; // 2799 : 172 - 0xac
      12'hAF0: dout <= 8'b01010110; // 2800 :  86 - 0x56 -- Sprite 0xaf
      12'hAF1: dout <= 8'b00001100; // 2801 :  12 - 0xc
      12'hAF2: dout <= 8'b00001110; // 2802 :  14 - 0xe
      12'hAF3: dout <= 8'b00011111; // 2803 :  31 - 0x1f
      12'hAF4: dout <= 8'b11111111; // 2804 : 255 - 0xff
      12'hAF5: dout <= 8'b11111111; // 2805 : 255 - 0xff
      12'hAF6: dout <= 8'b11111110; // 2806 : 254 - 0xfe
      12'hAF7: dout <= 8'b11111000; // 2807 : 248 - 0xf8
      12'hAF8: dout <= 8'b10101100; // 2808 : 172 - 0xac -- plane 1
      12'hAF9: dout <= 8'b11111000; // 2809 : 248 - 0xf8
      12'hAFA: dout <= 8'b11111000; // 2810 : 248 - 0xf8
      12'hAFB: dout <= 8'b11111100; // 2811 : 252 - 0xfc
      12'hAFC: dout <= 8'b11111100; // 2812 : 252 - 0xfc
      12'hAFD: dout <= 8'b11111000; // 2813 : 248 - 0xf8
      12'hAFE: dout <= 8'b11110000; // 2814 : 240 - 0xf0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b11111111; // 2816 : 255 - 0xff -- Sprite 0xb0
      12'hB01: dout <= 8'b11111111; // 2817 : 255 - 0xff
      12'hB02: dout <= 8'b11111111; // 2818 : 255 - 0xff
      12'hB03: dout <= 8'b11111111; // 2819 : 255 - 0xff
      12'hB04: dout <= 8'b11111111; // 2820 : 255 - 0xff
      12'hB05: dout <= 8'b11111111; // 2821 : 255 - 0xff
      12'hB06: dout <= 8'b11111111; // 2822 : 255 - 0xff
      12'hB07: dout <= 8'b11111111; // 2823 : 255 - 0xff
      12'hB08: dout <= 8'b11111111; // 2824 : 255 - 0xff -- plane 1
      12'hB09: dout <= 8'b11111111; // 2825 : 255 - 0xff
      12'hB0A: dout <= 8'b11111111; // 2826 : 255 - 0xff
      12'hB0B: dout <= 8'b11111111; // 2827 : 255 - 0xff
      12'hB0C: dout <= 8'b11111111; // 2828 : 255 - 0xff
      12'hB0D: dout <= 8'b11111111; // 2829 : 255 - 0xff
      12'hB0E: dout <= 8'b11111111; // 2830 : 255 - 0xff
      12'hB0F: dout <= 8'b11111111; // 2831 : 255 - 0xff
      12'hB10: dout <= 8'b11111111; // 2832 : 255 - 0xff -- Sprite 0xb1
      12'hB11: dout <= 8'b11111111; // 2833 : 255 - 0xff
      12'hB12: dout <= 8'b11111111; // 2834 : 255 - 0xff
      12'hB13: dout <= 8'b11111111; // 2835 : 255 - 0xff
      12'hB14: dout <= 8'b11111111; // 2836 : 255 - 0xff
      12'hB15: dout <= 8'b11111111; // 2837 : 255 - 0xff
      12'hB16: dout <= 8'b11111111; // 2838 : 255 - 0xff
      12'hB17: dout <= 8'b11111111; // 2839 : 255 - 0xff
      12'hB18: dout <= 8'b11111111; // 2840 : 255 - 0xff -- plane 1
      12'hB19: dout <= 8'b11111111; // 2841 : 255 - 0xff
      12'hB1A: dout <= 8'b11111111; // 2842 : 255 - 0xff
      12'hB1B: dout <= 8'b11111111; // 2843 : 255 - 0xff
      12'hB1C: dout <= 8'b11111111; // 2844 : 255 - 0xff
      12'hB1D: dout <= 8'b11111111; // 2845 : 255 - 0xff
      12'hB1E: dout <= 8'b11111111; // 2846 : 255 - 0xff
      12'hB1F: dout <= 8'b11111111; // 2847 : 255 - 0xff
      12'hB20: dout <= 8'b11111111; // 2848 : 255 - 0xff -- Sprite 0xb2
      12'hB21: dout <= 8'b11111111; // 2849 : 255 - 0xff
      12'hB22: dout <= 8'b11111111; // 2850 : 255 - 0xff
      12'hB23: dout <= 8'b11111111; // 2851 : 255 - 0xff
      12'hB24: dout <= 8'b11111111; // 2852 : 255 - 0xff
      12'hB25: dout <= 8'b11111111; // 2853 : 255 - 0xff
      12'hB26: dout <= 8'b11111111; // 2854 : 255 - 0xff
      12'hB27: dout <= 8'b11111111; // 2855 : 255 - 0xff
      12'hB28: dout <= 8'b11111111; // 2856 : 255 - 0xff -- plane 1
      12'hB29: dout <= 8'b11111111; // 2857 : 255 - 0xff
      12'hB2A: dout <= 8'b11111111; // 2858 : 255 - 0xff
      12'hB2B: dout <= 8'b11111111; // 2859 : 255 - 0xff
      12'hB2C: dout <= 8'b11111111; // 2860 : 255 - 0xff
      12'hB2D: dout <= 8'b11111111; // 2861 : 255 - 0xff
      12'hB2E: dout <= 8'b11111111; // 2862 : 255 - 0xff
      12'hB2F: dout <= 8'b11111111; // 2863 : 255 - 0xff
      12'hB30: dout <= 8'b11111111; // 2864 : 255 - 0xff -- Sprite 0xb3
      12'hB31: dout <= 8'b11111111; // 2865 : 255 - 0xff
      12'hB32: dout <= 8'b11111111; // 2866 : 255 - 0xff
      12'hB33: dout <= 8'b11111111; // 2867 : 255 - 0xff
      12'hB34: dout <= 8'b11111111; // 2868 : 255 - 0xff
      12'hB35: dout <= 8'b11111111; // 2869 : 255 - 0xff
      12'hB36: dout <= 8'b11111111; // 2870 : 255 - 0xff
      12'hB37: dout <= 8'b11111111; // 2871 : 255 - 0xff
      12'hB38: dout <= 8'b11111111; // 2872 : 255 - 0xff -- plane 1
      12'hB39: dout <= 8'b11111111; // 2873 : 255 - 0xff
      12'hB3A: dout <= 8'b11111111; // 2874 : 255 - 0xff
      12'hB3B: dout <= 8'b11111111; // 2875 : 255 - 0xff
      12'hB3C: dout <= 8'b11111111; // 2876 : 255 - 0xff
      12'hB3D: dout <= 8'b11111111; // 2877 : 255 - 0xff
      12'hB3E: dout <= 8'b11111111; // 2878 : 255 - 0xff
      12'hB3F: dout <= 8'b11111111; // 2879 : 255 - 0xff
      12'hB40: dout <= 8'b11111111; // 2880 : 255 - 0xff -- Sprite 0xb4
      12'hB41: dout <= 8'b11111111; // 2881 : 255 - 0xff
      12'hB42: dout <= 8'b11111111; // 2882 : 255 - 0xff
      12'hB43: dout <= 8'b11111111; // 2883 : 255 - 0xff
      12'hB44: dout <= 8'b11111111; // 2884 : 255 - 0xff
      12'hB45: dout <= 8'b11111111; // 2885 : 255 - 0xff
      12'hB46: dout <= 8'b11111111; // 2886 : 255 - 0xff
      12'hB47: dout <= 8'b11111111; // 2887 : 255 - 0xff
      12'hB48: dout <= 8'b11111111; // 2888 : 255 - 0xff -- plane 1
      12'hB49: dout <= 8'b11111111; // 2889 : 255 - 0xff
      12'hB4A: dout <= 8'b11111111; // 2890 : 255 - 0xff
      12'hB4B: dout <= 8'b11111111; // 2891 : 255 - 0xff
      12'hB4C: dout <= 8'b11111111; // 2892 : 255 - 0xff
      12'hB4D: dout <= 8'b11111111; // 2893 : 255 - 0xff
      12'hB4E: dout <= 8'b11111111; // 2894 : 255 - 0xff
      12'hB4F: dout <= 8'b11111111; // 2895 : 255 - 0xff
      12'hB50: dout <= 8'b11111111; // 2896 : 255 - 0xff -- Sprite 0xb5
      12'hB51: dout <= 8'b11111111; // 2897 : 255 - 0xff
      12'hB52: dout <= 8'b11111111; // 2898 : 255 - 0xff
      12'hB53: dout <= 8'b11111111; // 2899 : 255 - 0xff
      12'hB54: dout <= 8'b11111111; // 2900 : 255 - 0xff
      12'hB55: dout <= 8'b11111111; // 2901 : 255 - 0xff
      12'hB56: dout <= 8'b11111111; // 2902 : 255 - 0xff
      12'hB57: dout <= 8'b11111111; // 2903 : 255 - 0xff
      12'hB58: dout <= 8'b11111111; // 2904 : 255 - 0xff -- plane 1
      12'hB59: dout <= 8'b11111111; // 2905 : 255 - 0xff
      12'hB5A: dout <= 8'b11111111; // 2906 : 255 - 0xff
      12'hB5B: dout <= 8'b11111111; // 2907 : 255 - 0xff
      12'hB5C: dout <= 8'b11111111; // 2908 : 255 - 0xff
      12'hB5D: dout <= 8'b11111111; // 2909 : 255 - 0xff
      12'hB5E: dout <= 8'b11111111; // 2910 : 255 - 0xff
      12'hB5F: dout <= 8'b11111111; // 2911 : 255 - 0xff
      12'hB60: dout <= 8'b11111111; // 2912 : 255 - 0xff -- Sprite 0xb6
      12'hB61: dout <= 8'b11111111; // 2913 : 255 - 0xff
      12'hB62: dout <= 8'b11111111; // 2914 : 255 - 0xff
      12'hB63: dout <= 8'b11111111; // 2915 : 255 - 0xff
      12'hB64: dout <= 8'b11111111; // 2916 : 255 - 0xff
      12'hB65: dout <= 8'b11111111; // 2917 : 255 - 0xff
      12'hB66: dout <= 8'b11111111; // 2918 : 255 - 0xff
      12'hB67: dout <= 8'b11111111; // 2919 : 255 - 0xff
      12'hB68: dout <= 8'b11111111; // 2920 : 255 - 0xff -- plane 1
      12'hB69: dout <= 8'b11111111; // 2921 : 255 - 0xff
      12'hB6A: dout <= 8'b11111111; // 2922 : 255 - 0xff
      12'hB6B: dout <= 8'b11111111; // 2923 : 255 - 0xff
      12'hB6C: dout <= 8'b11111111; // 2924 : 255 - 0xff
      12'hB6D: dout <= 8'b11111111; // 2925 : 255 - 0xff
      12'hB6E: dout <= 8'b11111111; // 2926 : 255 - 0xff
      12'hB6F: dout <= 8'b11111111; // 2927 : 255 - 0xff
      12'hB70: dout <= 8'b11111111; // 2928 : 255 - 0xff -- Sprite 0xb7
      12'hB71: dout <= 8'b11111111; // 2929 : 255 - 0xff
      12'hB72: dout <= 8'b11111111; // 2930 : 255 - 0xff
      12'hB73: dout <= 8'b11111111; // 2931 : 255 - 0xff
      12'hB74: dout <= 8'b11111111; // 2932 : 255 - 0xff
      12'hB75: dout <= 8'b11111111; // 2933 : 255 - 0xff
      12'hB76: dout <= 8'b11111111; // 2934 : 255 - 0xff
      12'hB77: dout <= 8'b11111111; // 2935 : 255 - 0xff
      12'hB78: dout <= 8'b11111111; // 2936 : 255 - 0xff -- plane 1
      12'hB79: dout <= 8'b11111111; // 2937 : 255 - 0xff
      12'hB7A: dout <= 8'b11111111; // 2938 : 255 - 0xff
      12'hB7B: dout <= 8'b11111111; // 2939 : 255 - 0xff
      12'hB7C: dout <= 8'b11111111; // 2940 : 255 - 0xff
      12'hB7D: dout <= 8'b11111111; // 2941 : 255 - 0xff
      12'hB7E: dout <= 8'b11111111; // 2942 : 255 - 0xff
      12'hB7F: dout <= 8'b11111111; // 2943 : 255 - 0xff
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Sprite 0xb8
      12'hB81: dout <= 8'b00000111; // 2945 :   7 - 0x7
      12'hB82: dout <= 8'b00001000; // 2946 :   8 - 0x8
      12'hB83: dout <= 8'b00010000; // 2947 :  16 - 0x10
      12'hB84: dout <= 8'b00010000; // 2948 :  16 - 0x10
      12'hB85: dout <= 8'b00100000; // 2949 :  32 - 0x20
      12'hB86: dout <= 8'b00100000; // 2950 :  32 - 0x20
      12'hB87: dout <= 8'b00100000; // 2951 :  32 - 0x20
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout <= 8'b00000111; // 2953 :   7 - 0x7
      12'hB8A: dout <= 8'b00001000; // 2954 :   8 - 0x8
      12'hB8B: dout <= 8'b00010000; // 2955 :  16 - 0x10
      12'hB8C: dout <= 8'b00010000; // 2956 :  16 - 0x10
      12'hB8D: dout <= 8'b00100000; // 2957 :  32 - 0x20
      12'hB8E: dout <= 8'b00100000; // 2958 :  32 - 0x20
      12'hB8F: dout <= 8'b00100000; // 2959 :  32 - 0x20
      12'hB90: dout <= 8'b00011111; // 2960 :  31 - 0x1f -- Sprite 0xb9
      12'hB91: dout <= 8'b00101111; // 2961 :  47 - 0x2f
      12'hB92: dout <= 8'b00110111; // 2962 :  55 - 0x37
      12'hB93: dout <= 8'b00111010; // 2963 :  58 - 0x3a
      12'hB94: dout <= 8'b00111101; // 2964 :  61 - 0x3d
      12'hB95: dout <= 8'b00111110; // 2965 :  62 - 0x3e
      12'hB96: dout <= 8'b00111111; // 2966 :  63 - 0x3f
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00011111; // 2968 :  31 - 0x1f -- plane 1
      12'hB99: dout <= 8'b00111111; // 2969 :  63 - 0x3f
      12'hB9A: dout <= 8'b00111111; // 2970 :  63 - 0x3f
      12'hB9B: dout <= 8'b00111111; // 2971 :  63 - 0x3f
      12'hB9C: dout <= 8'b00111110; // 2972 :  62 - 0x3e
      12'hB9D: dout <= 8'b00111111; // 2973 :  63 - 0x3f
      12'hB9E: dout <= 8'b00111111; // 2974 :  63 - 0x3f
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Sprite 0xba
      12'hBA1: dout <= 8'b00000101; // 2977 :   5 - 0x5
      12'hBA2: dout <= 8'b00011001; // 2978 :  25 - 0x19
      12'hBA3: dout <= 8'b00110011; // 2979 :  51 - 0x33
      12'hBA4: dout <= 8'b01100011; // 2980 :  99 - 0x63
      12'hBA5: dout <= 8'b11000111; // 2981 : 199 - 0xc7
      12'hBA6: dout <= 8'b11000111; // 2982 : 199 - 0xc7
      12'hBA7: dout <= 8'b11000100; // 2983 : 196 - 0xc4
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout <= 8'b00000111; // 2985 :   7 - 0x7
      12'hBAA: dout <= 8'b00011111; // 2986 :  31 - 0x1f
      12'hBAB: dout <= 8'b00111111; // 2987 :  63 - 0x3f
      12'hBAC: dout <= 8'b01111111; // 2988 : 127 - 0x7f
      12'hBAD: dout <= 8'b11111111; // 2989 : 255 - 0xff
      12'hBAE: dout <= 8'b11111111; // 2990 : 255 - 0xff
      12'hBAF: dout <= 8'b11011101; // 2991 : 221 - 0xdd
      12'hBB0: dout <= 8'b10000000; // 2992 : 128 - 0x80 -- Sprite 0xbb
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000011; // 2997 :   3 - 0x3
      12'hBB6: dout <= 8'b00000011; // 2998 :   3 - 0x3
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b10001001; // 3000 : 137 - 0x89 -- plane 1
      12'hBB9: dout <= 8'b00000001; // 3001 :   1 - 0x1
      12'hBBA: dout <= 8'b00000001; // 3002 :   1 - 0x1
      12'hBBB: dout <= 8'b00000001; // 3003 :   1 - 0x1
      12'hBBC: dout <= 8'b00000001; // 3004 :   1 - 0x1
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Sprite 0xbc
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- plane 1
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000011; // 3022 :   3 - 0x3
      12'hBCF: dout <= 8'b00000111; // 3023 :   7 - 0x7
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00001111; // 3026 :  15 - 0xf
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b10000000; // 3028 : 128 - 0x80
      12'hBD5: dout <= 8'b01100011; // 3029 :  99 - 0x63
      12'hBD6: dout <= 8'b00011110; // 3030 :  30 - 0x1e
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00001111; // 3032 :  15 - 0xf -- plane 1
      12'hBD9: dout <= 8'b00001111; // 3033 :  15 - 0xf
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00011111; // 3035 :  31 - 0x1f
      12'hBDC: dout <= 8'b01111111; // 3036 : 127 - 0x7f
      12'hBDD: dout <= 8'b00011100; // 3037 :  28 - 0x1c
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000001; // 3040 :   1 - 0x1 -- Sprite 0xbe
      12'hBE1: dout <= 8'b00000011; // 3041 :   3 - 0x3
      12'hBE2: dout <= 8'b00011001; // 3042 :  25 - 0x19
      12'hBE3: dout <= 8'b00111100; // 3043 :  60 - 0x3c
      12'hBE4: dout <= 8'b00011001; // 3044 :  25 - 0x19
      12'hBE5: dout <= 8'b00100011; // 3045 :  35 - 0x23
      12'hBE6: dout <= 8'b01010001; // 3046 :  81 - 0x51
      12'hBE7: dout <= 8'b00100000; // 3047 :  32 - 0x20
      12'hBE8: dout <= 8'b00000001; // 3048 :   1 - 0x1 -- plane 1
      12'hBE9: dout <= 8'b00000010; // 3049 :   2 - 0x2
      12'hBEA: dout <= 8'b00011001; // 3050 :  25 - 0x19
      12'hBEB: dout <= 8'b00100100; // 3051 :  36 - 0x24
      12'hBEC: dout <= 8'b00011001; // 3052 :  25 - 0x19
      12'hBED: dout <= 8'b00100010; // 3053 :  34 - 0x22
      12'hBEE: dout <= 8'b00010001; // 3054 :  17 - 0x11
      12'hBEF: dout <= 8'b00101100; // 3055 :  44 - 0x2c
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00011111; // 3064 :  31 - 0x1f -- plane 1
      12'hBF9: dout <= 8'b00000111; // 3065 :   7 - 0x7
      12'hBFA: dout <= 8'b00000011; // 3066 :   3 - 0x3
      12'hBFB: dout <= 8'b00000011; // 3067 :   3 - 0x3
      12'hBFC: dout <= 8'b00000001; // 3068 :   1 - 0x1
      12'hBFD: dout <= 8'b00000001; // 3069 :   1 - 0x1
      12'hBFE: dout <= 8'b00000001; // 3070 :   1 - 0x1
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      12'hC01: dout <= 8'b00111111; // 3073 :  63 - 0x3f
      12'hC02: dout <= 8'b00011111; // 3074 :  31 - 0x1f
      12'hC03: dout <= 8'b00000000; // 3075 :   0 - 0x0
      12'hC04: dout <= 8'b00000001; // 3076 :   1 - 0x1
      12'hC05: dout <= 8'b00000000; // 3077 :   0 - 0x0
      12'hC06: dout <= 8'b00000001; // 3078 :   1 - 0x1
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000001; // 3083 :   1 - 0x1
      12'hC0C: dout <= 8'b00000011; // 3084 :   3 - 0x3
      12'hC0D: dout <= 8'b00000111; // 3085 :   7 - 0x7
      12'hC0E: dout <= 8'b00001101; // 3086 :  13 - 0xd
      12'hC0F: dout <= 8'b00011001; // 3087 :  25 - 0x19
      12'hC10: dout <= 8'b00010001; // 3088 :  17 - 0x11 -- Sprite 0xc1
      12'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout <= 8'b00000001; // 3090 :   1 - 0x1
      12'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout <= 8'b00000001; // 3092 :   1 - 0x1
      12'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout <= 8'b00011111; // 3094 :  31 - 0x1f
      12'hC17: dout <= 8'b00111111; // 3095 :  63 - 0x3f
      12'hC18: dout <= 8'b00101001; // 3096 :  41 - 0x29 -- plane 1
      12'hC19: dout <= 8'b00011001; // 3097 :  25 - 0x19
      12'hC1A: dout <= 8'b00001101; // 3098 :  13 - 0xd
      12'hC1B: dout <= 8'b00000111; // 3099 :   7 - 0x7
      12'hC1C: dout <= 8'b00000011; // 3100 :   3 - 0x3
      12'hC1D: dout <= 8'b00000001; // 3101 :   1 - 0x1
      12'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      12'hC21: dout <= 8'b11111100; // 3105 : 252 - 0xfc
      12'hC22: dout <= 8'b11111000; // 3106 : 248 - 0xf8
      12'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout <= 8'b10000000; // 3108 : 128 - 0x80
      12'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout <= 8'b10000000; // 3110 : 128 - 0x80
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b10000000; // 3115 : 128 - 0x80
      12'hC2C: dout <= 8'b11000000; // 3116 : 192 - 0xc0
      12'hC2D: dout <= 8'b11100000; // 3117 : 224 - 0xe0
      12'hC2E: dout <= 8'b10110000; // 3118 : 176 - 0xb0
      12'hC2F: dout <= 8'b10011000; // 3119 : 152 - 0x98
      12'hC30: dout <= 8'b10001000; // 3120 : 136 - 0x88 -- Sprite 0xc3
      12'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout <= 8'b10000000; // 3122 : 128 - 0x80
      12'hC33: dout <= 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout <= 8'b10000000; // 3124 : 128 - 0x80
      12'hC35: dout <= 8'b00000000; // 3125 :   0 - 0x0
      12'hC36: dout <= 8'b11111000; // 3126 : 248 - 0xf8
      12'hC37: dout <= 8'b11111100; // 3127 : 252 - 0xfc
      12'hC38: dout <= 8'b10010100; // 3128 : 148 - 0x94 -- plane 1
      12'hC39: dout <= 8'b10011000; // 3129 : 152 - 0x98
      12'hC3A: dout <= 8'b10110000; // 3130 : 176 - 0xb0
      12'hC3B: dout <= 8'b11100000; // 3131 : 224 - 0xe0
      12'hC3C: dout <= 8'b11000000; // 3132 : 192 - 0xc0
      12'hC3D: dout <= 8'b10000000; // 3133 : 128 - 0x80
      12'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      12'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout <= 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout <= 8'b00000000; // 3139 :   0 - 0x0
      12'hC44: dout <= 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout <= 8'b00111111; // 3141 :  63 - 0x3f
      12'hC46: dout <= 8'b00011111; // 3142 :  31 - 0x1f
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      12'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout <= 8'b00000001; // 3151 :   1 - 0x1
      12'hC50: dout <= 8'b00000001; // 3152 :   1 - 0x1 -- Sprite 0xc5
      12'hC51: dout <= 8'b00000001; // 3153 :   1 - 0x1
      12'hC52: dout <= 8'b01000001; // 3154 :  65 - 0x41
      12'hC53: dout <= 8'b00000001; // 3155 :   1 - 0x1
      12'hC54: dout <= 8'b00000001; // 3156 :   1 - 0x1
      12'hC55: dout <= 8'b00000000; // 3157 :   0 - 0x0
      12'hC56: dout <= 8'b00011111; // 3158 :  31 - 0x1f
      12'hC57: dout <= 8'b00111111; // 3159 :  63 - 0x3f
      12'hC58: dout <= 8'b00001111; // 3160 :  15 - 0xf -- plane 1
      12'hC59: dout <= 8'b01111001; // 3161 : 121 - 0x79
      12'hC5A: dout <= 8'b10100001; // 3162 : 161 - 0xa1
      12'hC5B: dout <= 8'b01111001; // 3163 : 121 - 0x79
      12'hC5C: dout <= 8'b00001111; // 3164 :  15 - 0xf
      12'hC5D: dout <= 8'b00000001; // 3165 :   1 - 0x1
      12'hC5E: dout <= 8'b00000000; // 3166 :   0 - 0x0
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b00000000; // 3168 :   0 - 0x0 -- Sprite 0xc6
      12'hC61: dout <= 8'b00000000; // 3169 :   0 - 0x0
      12'hC62: dout <= 8'b00000000; // 3170 :   0 - 0x0
      12'hC63: dout <= 8'b00000000; // 3171 :   0 - 0x0
      12'hC64: dout <= 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout <= 8'b11111100; // 3173 : 252 - 0xfc
      12'hC66: dout <= 8'b11111000; // 3174 : 248 - 0xf8
      12'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout <= 8'b00000000; // 3177 :   0 - 0x0
      12'hC6A: dout <= 8'b00000000; // 3178 :   0 - 0x0
      12'hC6B: dout <= 8'b00000000; // 3179 :   0 - 0x0
      12'hC6C: dout <= 8'b00000000; // 3180 :   0 - 0x0
      12'hC6D: dout <= 8'b00000000; // 3181 :   0 - 0x0
      12'hC6E: dout <= 8'b00000000; // 3182 :   0 - 0x0
      12'hC6F: dout <= 8'b10000000; // 3183 : 128 - 0x80
      12'hC70: dout <= 8'b10000000; // 3184 : 128 - 0x80 -- Sprite 0xc7
      12'hC71: dout <= 8'b10000000; // 3185 : 128 - 0x80
      12'hC72: dout <= 8'b10000010; // 3186 : 130 - 0x82
      12'hC73: dout <= 8'b10000000; // 3187 : 128 - 0x80
      12'hC74: dout <= 8'b10000000; // 3188 : 128 - 0x80
      12'hC75: dout <= 8'b00000000; // 3189 :   0 - 0x0
      12'hC76: dout <= 8'b11111000; // 3190 : 248 - 0xf8
      12'hC77: dout <= 8'b11111100; // 3191 : 252 - 0xfc
      12'hC78: dout <= 8'b11110000; // 3192 : 240 - 0xf0 -- plane 1
      12'hC79: dout <= 8'b10011110; // 3193 : 158 - 0x9e
      12'hC7A: dout <= 8'b10000101; // 3194 : 133 - 0x85
      12'hC7B: dout <= 8'b10011110; // 3195 : 158 - 0x9e
      12'hC7C: dout <= 8'b11110000; // 3196 : 240 - 0xf0
      12'hC7D: dout <= 8'b10000000; // 3197 : 128 - 0x80
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00011110; // 3203 :  30 - 0x1e
      12'hC84: dout <= 8'b00111111; // 3204 :  63 - 0x3f
      12'hC85: dout <= 8'b00111111; // 3205 :  63 - 0x3f
      12'hC86: dout <= 8'b00111111; // 3206 :  63 - 0x3f
      12'hC87: dout <= 8'b00111111; // 3207 :  63 - 0x3f
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout <= 8'b00011110; // 3211 :  30 - 0x1e
      12'hC8C: dout <= 8'b00111111; // 3212 :  63 - 0x3f
      12'hC8D: dout <= 8'b00111111; // 3213 :  63 - 0x3f
      12'hC8E: dout <= 8'b00111111; // 3214 :  63 - 0x3f
      12'hC8F: dout <= 8'b00111111; // 3215 :  63 - 0x3f
      12'hC90: dout <= 8'b00011111; // 3216 :  31 - 0x1f -- Sprite 0xc9
      12'hC91: dout <= 8'b00001111; // 3217 :  15 - 0xf
      12'hC92: dout <= 8'b00000111; // 3218 :   7 - 0x7
      12'hC93: dout <= 8'b00000011; // 3219 :   3 - 0x3
      12'hC94: dout <= 8'b00000001; // 3220 :   1 - 0x1
      12'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      12'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b00011111; // 3224 :  31 - 0x1f -- plane 1
      12'hC99: dout <= 8'b00001111; // 3225 :  15 - 0xf
      12'hC9A: dout <= 8'b00000111; // 3226 :   7 - 0x7
      12'hC9B: dout <= 8'b00000011; // 3227 :   3 - 0x3
      12'hC9C: dout <= 8'b00000001; // 3228 :   1 - 0x1
      12'hC9D: dout <= 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      12'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout <= 8'b00000000; // 3234 :   0 - 0x0
      12'hCA3: dout <= 8'b00111100; // 3235 :  60 - 0x3c
      12'hCA4: dout <= 8'b01111110; // 3236 : 126 - 0x7e
      12'hCA5: dout <= 8'b11111110; // 3237 : 254 - 0xfe
      12'hCA6: dout <= 8'b11111110; // 3238 : 254 - 0xfe
      12'hCA7: dout <= 8'b11111110; // 3239 : 254 - 0xfe
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      12'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      12'hCAB: dout <= 8'b00111100; // 3243 :  60 - 0x3c
      12'hCAC: dout <= 8'b01111110; // 3244 : 126 - 0x7e
      12'hCAD: dout <= 8'b11111110; // 3245 : 254 - 0xfe
      12'hCAE: dout <= 8'b11111110; // 3246 : 254 - 0xfe
      12'hCAF: dout <= 8'b11111110; // 3247 : 254 - 0xfe
      12'hCB0: dout <= 8'b11111100; // 3248 : 252 - 0xfc -- Sprite 0xcb
      12'hCB1: dout <= 8'b11111000; // 3249 : 248 - 0xf8
      12'hCB2: dout <= 8'b11110000; // 3250 : 240 - 0xf0
      12'hCB3: dout <= 8'b11100000; // 3251 : 224 - 0xe0
      12'hCB4: dout <= 8'b11000000; // 3252 : 192 - 0xc0
      12'hCB5: dout <= 8'b10000000; // 3253 : 128 - 0x80
      12'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      12'hCB8: dout <= 8'b11111100; // 3256 : 252 - 0xfc -- plane 1
      12'hCB9: dout <= 8'b11111000; // 3257 : 248 - 0xf8
      12'hCBA: dout <= 8'b11110000; // 3258 : 240 - 0xf0
      12'hCBB: dout <= 8'b11100000; // 3259 : 224 - 0xe0
      12'hCBC: dout <= 8'b11000000; // 3260 : 192 - 0xc0
      12'hCBD: dout <= 8'b10000000; // 3261 : 128 - 0x80
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b11111111; // 3264 : 255 - 0xff -- Sprite 0xcc
      12'hCC1: dout <= 8'b11111111; // 3265 : 255 - 0xff
      12'hCC2: dout <= 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout <= 8'b11111111; // 3267 : 255 - 0xff
      12'hCC4: dout <= 8'b11111111; // 3268 : 255 - 0xff
      12'hCC5: dout <= 8'b11111111; // 3269 : 255 - 0xff
      12'hCC6: dout <= 8'b11111111; // 3270 : 255 - 0xff
      12'hCC7: dout <= 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout <= 8'b11111111; // 3272 : 255 - 0xff -- plane 1
      12'hCC9: dout <= 8'b11111111; // 3273 : 255 - 0xff
      12'hCCA: dout <= 8'b11111111; // 3274 : 255 - 0xff
      12'hCCB: dout <= 8'b11111111; // 3275 : 255 - 0xff
      12'hCCC: dout <= 8'b11111111; // 3276 : 255 - 0xff
      12'hCCD: dout <= 8'b11111111; // 3277 : 255 - 0xff
      12'hCCE: dout <= 8'b11111111; // 3278 : 255 - 0xff
      12'hCCF: dout <= 8'b11111111; // 3279 : 255 - 0xff
      12'hCD0: dout <= 8'b11111111; // 3280 : 255 - 0xff -- Sprite 0xcd
      12'hCD1: dout <= 8'b11111111; // 3281 : 255 - 0xff
      12'hCD2: dout <= 8'b11111111; // 3282 : 255 - 0xff
      12'hCD3: dout <= 8'b11111111; // 3283 : 255 - 0xff
      12'hCD4: dout <= 8'b11111111; // 3284 : 255 - 0xff
      12'hCD5: dout <= 8'b11111111; // 3285 : 255 - 0xff
      12'hCD6: dout <= 8'b11111111; // 3286 : 255 - 0xff
      12'hCD7: dout <= 8'b11111111; // 3287 : 255 - 0xff
      12'hCD8: dout <= 8'b11111111; // 3288 : 255 - 0xff -- plane 1
      12'hCD9: dout <= 8'b11111111; // 3289 : 255 - 0xff
      12'hCDA: dout <= 8'b11111111; // 3290 : 255 - 0xff
      12'hCDB: dout <= 8'b11111111; // 3291 : 255 - 0xff
      12'hCDC: dout <= 8'b11111111; // 3292 : 255 - 0xff
      12'hCDD: dout <= 8'b11111111; // 3293 : 255 - 0xff
      12'hCDE: dout <= 8'b11111111; // 3294 : 255 - 0xff
      12'hCDF: dout <= 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout <= 8'b11111111; // 3296 : 255 - 0xff -- Sprite 0xce
      12'hCE1: dout <= 8'b11111111; // 3297 : 255 - 0xff
      12'hCE2: dout <= 8'b11111111; // 3298 : 255 - 0xff
      12'hCE3: dout <= 8'b11111111; // 3299 : 255 - 0xff
      12'hCE4: dout <= 8'b11111111; // 3300 : 255 - 0xff
      12'hCE5: dout <= 8'b11111111; // 3301 : 255 - 0xff
      12'hCE6: dout <= 8'b11111111; // 3302 : 255 - 0xff
      12'hCE7: dout <= 8'b11111111; // 3303 : 255 - 0xff
      12'hCE8: dout <= 8'b11111111; // 3304 : 255 - 0xff -- plane 1
      12'hCE9: dout <= 8'b11111111; // 3305 : 255 - 0xff
      12'hCEA: dout <= 8'b11111111; // 3306 : 255 - 0xff
      12'hCEB: dout <= 8'b11111111; // 3307 : 255 - 0xff
      12'hCEC: dout <= 8'b11111111; // 3308 : 255 - 0xff
      12'hCED: dout <= 8'b11111111; // 3309 : 255 - 0xff
      12'hCEE: dout <= 8'b11111111; // 3310 : 255 - 0xff
      12'hCEF: dout <= 8'b11111111; // 3311 : 255 - 0xff
      12'hCF0: dout <= 8'b11111111; // 3312 : 255 - 0xff -- Sprite 0xcf
      12'hCF1: dout <= 8'b11111111; // 3313 : 255 - 0xff
      12'hCF2: dout <= 8'b11111111; // 3314 : 255 - 0xff
      12'hCF3: dout <= 8'b11111111; // 3315 : 255 - 0xff
      12'hCF4: dout <= 8'b11111111; // 3316 : 255 - 0xff
      12'hCF5: dout <= 8'b11111111; // 3317 : 255 - 0xff
      12'hCF6: dout <= 8'b11111111; // 3318 : 255 - 0xff
      12'hCF7: dout <= 8'b11111111; // 3319 : 255 - 0xff
      12'hCF8: dout <= 8'b11111111; // 3320 : 255 - 0xff -- plane 1
      12'hCF9: dout <= 8'b11111111; // 3321 : 255 - 0xff
      12'hCFA: dout <= 8'b11111111; // 3322 : 255 - 0xff
      12'hCFB: dout <= 8'b11111111; // 3323 : 255 - 0xff
      12'hCFC: dout <= 8'b11111111; // 3324 : 255 - 0xff
      12'hCFD: dout <= 8'b11111111; // 3325 : 255 - 0xff
      12'hCFE: dout <= 8'b11111111; // 3326 : 255 - 0xff
      12'hCFF: dout <= 8'b11111111; // 3327 : 255 - 0xff
      12'hD00: dout <= 8'b00001000; // 3328 :   8 - 0x8 -- Sprite 0xd0
      12'hD01: dout <= 8'b00011001; // 3329 :  25 - 0x19
      12'hD02: dout <= 8'b00001001; // 3330 :   9 - 0x9
      12'hD03: dout <= 8'b00001001; // 3331 :   9 - 0x9
      12'hD04: dout <= 8'b00001001; // 3332 :   9 - 0x9
      12'hD05: dout <= 8'b00001001; // 3333 :   9 - 0x9
      12'hD06: dout <= 8'b00011100; // 3334 :  28 - 0x1c
      12'hD07: dout <= 8'b00000000; // 3335 :   0 - 0x0
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b00000000; // 3338 :   0 - 0x0
      12'hD0B: dout <= 8'b00000000; // 3339 :   0 - 0x0
      12'hD0C: dout <= 8'b00000000; // 3340 :   0 - 0x0
      12'hD0D: dout <= 8'b00000000; // 3341 :   0 - 0x0
      12'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00111000; // 3344 :  56 - 0x38 -- Sprite 0xd1
      12'hD11: dout <= 8'b00000101; // 3345 :   5 - 0x5
      12'hD12: dout <= 8'b00000101; // 3346 :   5 - 0x5
      12'hD13: dout <= 8'b00011001; // 3347 :  25 - 0x19
      12'hD14: dout <= 8'b00000101; // 3348 :   5 - 0x5
      12'hD15: dout <= 8'b00000101; // 3349 :   5 - 0x5
      12'hD16: dout <= 8'b00111000; // 3350 :  56 - 0x38
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout <= 8'b00000000; // 3354 :   0 - 0x0
      12'hD1B: dout <= 8'b00000000; // 3355 :   0 - 0x0
      12'hD1C: dout <= 8'b00000000; // 3356 :   0 - 0x0
      12'hD1D: dout <= 8'b00000000; // 3357 :   0 - 0x0
      12'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00111100; // 3360 :  60 - 0x3c -- Sprite 0xd2
      12'hD21: dout <= 8'b00100001; // 3361 :  33 - 0x21
      12'hD22: dout <= 8'b00100001; // 3362 :  33 - 0x21
      12'hD23: dout <= 8'b00111101; // 3363 :  61 - 0x3d
      12'hD24: dout <= 8'b00000101; // 3364 :   5 - 0x5
      12'hD25: dout <= 8'b00000101; // 3365 :   5 - 0x5
      12'hD26: dout <= 8'b00111000; // 3366 :  56 - 0x38
      12'hD27: dout <= 8'b00000000; // 3367 :   0 - 0x0
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout <= 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout <= 8'b00000000; // 3372 :   0 - 0x0
      12'hD2D: dout <= 8'b00000000; // 3373 :   0 - 0x0
      12'hD2E: dout <= 8'b00000000; // 3374 :   0 - 0x0
      12'hD2F: dout <= 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout <= 8'b00011000; // 3376 :  24 - 0x18 -- Sprite 0xd3
      12'hD31: dout <= 8'b00100101; // 3377 :  37 - 0x25
      12'hD32: dout <= 8'b00100101; // 3378 :  37 - 0x25
      12'hD33: dout <= 8'b00011001; // 3379 :  25 - 0x19
      12'hD34: dout <= 8'b00100101; // 3380 :  37 - 0x25
      12'hD35: dout <= 8'b00100101; // 3381 :  37 - 0x25
      12'hD36: dout <= 8'b00011000; // 3382 :  24 - 0x18
      12'hD37: dout <= 8'b00000000; // 3383 :   0 - 0x0
      12'hD38: dout <= 8'b00000000; // 3384 :   0 - 0x0 -- plane 1
      12'hD39: dout <= 8'b00000000; // 3385 :   0 - 0x0
      12'hD3A: dout <= 8'b00000000; // 3386 :   0 - 0x0
      12'hD3B: dout <= 8'b00000000; // 3387 :   0 - 0x0
      12'hD3C: dout <= 8'b00000000; // 3388 :   0 - 0x0
      12'hD3D: dout <= 8'b00000000; // 3389 :   0 - 0x0
      12'hD3E: dout <= 8'b00000000; // 3390 :   0 - 0x0
      12'hD3F: dout <= 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout <= 8'b11000110; // 3392 : 198 - 0xc6 -- Sprite 0xd4
      12'hD41: dout <= 8'b00101001; // 3393 :  41 - 0x29
      12'hD42: dout <= 8'b00101001; // 3394 :  41 - 0x29
      12'hD43: dout <= 8'b00101001; // 3395 :  41 - 0x29
      12'hD44: dout <= 8'b00101001; // 3396 :  41 - 0x29
      12'hD45: dout <= 8'b00101001; // 3397 :  41 - 0x29
      12'hD46: dout <= 8'b11000110; // 3398 : 198 - 0xc6
      12'hD47: dout <= 8'b00000000; // 3399 :   0 - 0x0
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      12'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      12'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b00000000; // 3408 :   0 - 0x0 -- Sprite 0xd5
      12'hD51: dout <= 8'b00000000; // 3409 :   0 - 0x0
      12'hD52: dout <= 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      12'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout <= 8'b00000000; // 3413 :   0 - 0x0
      12'hD56: dout <= 8'b00000000; // 3414 :   0 - 0x0
      12'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout <= 8'b00000001; // 3419 :   1 - 0x1
      12'hD5C: dout <= 8'b00000011; // 3420 :   3 - 0x3
      12'hD5D: dout <= 8'b01100011; // 3421 :  99 - 0x63
      12'hD5E: dout <= 8'b00110001; // 3422 :  49 - 0x31
      12'hD5F: dout <= 8'b00011111; // 3423 :  31 - 0x1f
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout <= 8'b00000000; // 3427 :   0 - 0x0
      12'hD64: dout <= 8'b00111100; // 3428 :  60 - 0x3c
      12'hD65: dout <= 8'b10110110; // 3429 : 182 - 0xb6
      12'hD66: dout <= 8'b01111100; // 3430 : 124 - 0x7c
      12'hD67: dout <= 8'b11111000; // 3431 : 248 - 0xf8
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b11111100; // 3434 : 252 - 0xfc
      12'hD6B: dout <= 8'b11111110; // 3435 : 254 - 0xfe
      12'hD6C: dout <= 8'b11000000; // 3436 : 192 - 0xc0
      12'hD6D: dout <= 8'b01000000; // 3437 :  64 - 0x40
      12'hD6E: dout <= 8'b10000000; // 3438 : 128 - 0x80
      12'hD6F: dout <= 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout <= 8'b00000011; // 3440 :   3 - 0x3 -- Sprite 0xd7
      12'hD71: dout <= 8'b00000011; // 3441 :   3 - 0x3
      12'hD72: dout <= 8'b00000011; // 3442 :   3 - 0x3
      12'hD73: dout <= 8'b00000111; // 3443 :   7 - 0x7
      12'hD74: dout <= 8'b00001100; // 3444 :  12 - 0xc
      12'hD75: dout <= 8'b00011011; // 3445 :  27 - 0x1b
      12'hD76: dout <= 8'b01110111; // 3446 : 119 - 0x77
      12'hD77: dout <= 8'b00000111; // 3447 :   7 - 0x7
      12'hD78: dout <= 8'b01111111; // 3448 : 127 - 0x7f -- plane 1
      12'hD79: dout <= 8'b00111111; // 3449 :  63 - 0x3f
      12'hD7A: dout <= 8'b01010011; // 3450 :  83 - 0x53
      12'hD7B: dout <= 8'b00000111; // 3451 :   7 - 0x7
      12'hD7C: dout <= 8'b00001100; // 3452 :  12 - 0xc
      12'hD7D: dout <= 8'b00011011; // 3453 :  27 - 0x1b
      12'hD7E: dout <= 8'b00000111; // 3454 :   7 - 0x7
      12'hD7F: dout <= 8'b00000111; // 3455 :   7 - 0x7
      12'hD80: dout <= 8'b00001111; // 3456 :  15 - 0xf -- Sprite 0xd8
      12'hD81: dout <= 8'b00001111; // 3457 :  15 - 0xf
      12'hD82: dout <= 8'b00011111; // 3458 :  31 - 0x1f
      12'hD83: dout <= 8'b00111111; // 3459 :  63 - 0x3f
      12'hD84: dout <= 8'b01111111; // 3460 : 127 - 0x7f
      12'hD85: dout <= 8'b00111111; // 3461 :  63 - 0x3f
      12'hD86: dout <= 8'b00000000; // 3462 :   0 - 0x0
      12'hD87: dout <= 8'b00000000; // 3463 :   0 - 0x0
      12'hD88: dout <= 8'b00001111; // 3464 :  15 - 0xf -- plane 1
      12'hD89: dout <= 8'b00001111; // 3465 :  15 - 0xf
      12'hD8A: dout <= 8'b00000011; // 3466 :   3 - 0x3
      12'hD8B: dout <= 8'b00111000; // 3467 :  56 - 0x38
      12'hD8C: dout <= 8'b00111111; // 3468 :  63 - 0x3f
      12'hD8D: dout <= 8'b00001110; // 3469 :  14 - 0xe
      12'hD8E: dout <= 8'b00011100; // 3470 :  28 - 0x1c
      12'hD8F: dout <= 8'b00001110; // 3471 :  14 - 0xe
      12'hD90: dout <= 8'b11100000; // 3472 : 224 - 0xe0 -- Sprite 0xd9
      12'hD91: dout <= 8'b11110000; // 3473 : 240 - 0xf0
      12'hD92: dout <= 8'b11110000; // 3474 : 240 - 0xf0
      12'hD93: dout <= 8'b11110000; // 3475 : 240 - 0xf0
      12'hD94: dout <= 8'b00011000; // 3476 :  24 - 0x18
      12'hD95: dout <= 8'b11111100; // 3477 : 252 - 0xfc
      12'hD96: dout <= 8'b11111100; // 3478 : 252 - 0xfc
      12'hD97: dout <= 8'b11111100; // 3479 : 252 - 0xfc
      12'hD98: dout <= 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout <= 8'b10010000; // 3481 : 144 - 0x90
      12'hD9A: dout <= 8'b11110000; // 3482 : 240 - 0xf0
      12'hD9B: dout <= 8'b11110000; // 3483 : 240 - 0xf0
      12'hD9C: dout <= 8'b00011000; // 3484 :  24 - 0x18
      12'hD9D: dout <= 8'b11111100; // 3485 : 252 - 0xfc
      12'hD9E: dout <= 8'b11110000; // 3486 : 240 - 0xf0
      12'hD9F: dout <= 8'b11111000; // 3487 : 248 - 0xf8
      12'hDA0: dout <= 8'b11111000; // 3488 : 248 - 0xf8 -- Sprite 0xda
      12'hDA1: dout <= 8'b11111100; // 3489 : 252 - 0xfc
      12'hDA2: dout <= 8'b11111111; // 3490 : 255 - 0xff
      12'hDA3: dout <= 8'b11111111; // 3491 : 255 - 0xff
      12'hDA4: dout <= 8'b11111110; // 3492 : 254 - 0xfe
      12'hDA5: dout <= 8'b11110000; // 3493 : 240 - 0xf0
      12'hDA6: dout <= 8'b00000000; // 3494 :   0 - 0x0
      12'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout <= 8'b11111000; // 3496 : 248 - 0xf8 -- plane 1
      12'hDA9: dout <= 8'b11110000; // 3497 : 240 - 0xf0
      12'hDAA: dout <= 8'b10000111; // 3498 : 135 - 0x87
      12'hDAB: dout <= 8'b00111101; // 3499 :  61 - 0x3d
      12'hDAC: dout <= 8'b11111110; // 3500 : 254 - 0xfe
      12'hDAD: dout <= 8'b00011100; // 3501 :  28 - 0x1c
      12'hDAE: dout <= 8'b00001000; // 3502 :   8 - 0x8
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b00000011; // 3504 :   3 - 0x3 -- Sprite 0xdb
      12'hDB1: dout <= 8'b00000011; // 3505 :   3 - 0x3
      12'hDB2: dout <= 8'b00000011; // 3506 :   3 - 0x3
      12'hDB3: dout <= 8'b00000011; // 3507 :   3 - 0x3
      12'hDB4: dout <= 8'b00000001; // 3508 :   1 - 0x1
      12'hDB5: dout <= 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout <= 8'b00000111; // 3510 :   7 - 0x7
      12'hDB7: dout <= 8'b00011111; // 3511 :  31 - 0x1f
      12'hDB8: dout <= 8'b01111111; // 3512 : 127 - 0x7f -- plane 1
      12'hDB9: dout <= 8'b00111111; // 3513 :  63 - 0x3f
      12'hDBA: dout <= 8'b01010011; // 3514 :  83 - 0x53
      12'hDBB: dout <= 8'b00000011; // 3515 :   3 - 0x3
      12'hDBC: dout <= 8'b00000001; // 3516 :   1 - 0x1
      12'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout <= 8'b00000111; // 3518 :   7 - 0x7
      12'hDBF: dout <= 8'b00011111; // 3519 :  31 - 0x1f
      12'hDC0: dout <= 8'b11111111; // 3520 : 255 - 0xff -- Sprite 0xdc
      12'hDC1: dout <= 8'b11111111; // 3521 : 255 - 0xff
      12'hDC2: dout <= 8'b01111111; // 3522 : 127 - 0x7f
      12'hDC3: dout <= 8'b00111111; // 3523 :  63 - 0x3f
      12'hDC4: dout <= 8'b00001111; // 3524 :  15 - 0xf
      12'hDC5: dout <= 8'b00000011; // 3525 :   3 - 0x3
      12'hDC6: dout <= 8'b00000000; // 3526 :   0 - 0x0
      12'hDC7: dout <= 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout <= 8'b11001111; // 3528 : 207 - 0xcf -- plane 1
      12'hDC9: dout <= 8'b01100011; // 3529 :  99 - 0x63
      12'hDCA: dout <= 8'b00111000; // 3530 :  56 - 0x38
      12'hDCB: dout <= 8'b00111110; // 3531 :  62 - 0x3e
      12'hDCC: dout <= 8'b01111011; // 3532 : 123 - 0x7b
      12'hDCD: dout <= 8'b00110000; // 3533 :  48 - 0x30
      12'hDCE: dout <= 8'b00011000; // 3534 :  24 - 0x18
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b11100000; // 3536 : 224 - 0xe0 -- Sprite 0xdd
      12'hDD1: dout <= 8'b11110000; // 3537 : 240 - 0xf0
      12'hDD2: dout <= 8'b11110000; // 3538 : 240 - 0xf0
      12'hDD3: dout <= 8'b11100000; // 3539 : 224 - 0xe0
      12'hDD4: dout <= 8'b11111110; // 3540 : 254 - 0xfe
      12'hDD5: dout <= 8'b00111100; // 3541 :  60 - 0x3c
      12'hDD6: dout <= 8'b11110000; // 3542 : 240 - 0xf0
      12'hDD7: dout <= 8'b11111100; // 3543 : 252 - 0xfc
      12'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0 -- plane 1
      12'hDD9: dout <= 8'b10010000; // 3545 : 144 - 0x90
      12'hDDA: dout <= 8'b11110000; // 3546 : 240 - 0xf0
      12'hDDB: dout <= 8'b11100000; // 3547 : 224 - 0xe0
      12'hDDC: dout <= 8'b11111000; // 3548 : 248 - 0xf8
      12'hDDD: dout <= 8'b00111000; // 3549 :  56 - 0x38
      12'hDDE: dout <= 8'b11110000; // 3550 : 240 - 0xf0
      12'hDDF: dout <= 8'b11110000; // 3551 : 240 - 0xf0
      12'hDE0: dout <= 8'b11111100; // 3552 : 252 - 0xfc -- Sprite 0xde
      12'hDE1: dout <= 8'b11111000; // 3553 : 248 - 0xf8
      12'hDE2: dout <= 8'b11111000; // 3554 : 248 - 0xf8
      12'hDE3: dout <= 8'b11111000; // 3555 : 248 - 0xf8
      12'hDE4: dout <= 8'b11111000; // 3556 : 248 - 0xf8
      12'hDE5: dout <= 8'b11111000; // 3557 : 248 - 0xf8
      12'hDE6: dout <= 8'b11111000; // 3558 : 248 - 0xf8
      12'hDE7: dout <= 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout <= 8'b11111000; // 3560 : 248 - 0xf8 -- plane 1
      12'hDE9: dout <= 8'b11111000; // 3561 : 248 - 0xf8
      12'hDEA: dout <= 8'b11111000; // 3562 : 248 - 0xf8
      12'hDEB: dout <= 8'b00111000; // 3563 :  56 - 0x38
      12'hDEC: dout <= 8'b10000000; // 3564 : 128 - 0x80
      12'hDED: dout <= 8'b11111000; // 3565 : 248 - 0xf8
      12'hDEE: dout <= 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout <= 8'b01011100; // 3567 :  92 - 0x5c
      12'hDF0: dout <= 8'b11111111; // 3568 : 255 - 0xff -- Sprite 0xdf
      12'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout <= 8'b11111111; // 3570 : 255 - 0xff
      12'hDF3: dout <= 8'b11111111; // 3571 : 255 - 0xff
      12'hDF4: dout <= 8'b11111111; // 3572 : 255 - 0xff
      12'hDF5: dout <= 8'b11111111; // 3573 : 255 - 0xff
      12'hDF6: dout <= 8'b11111111; // 3574 : 255 - 0xff
      12'hDF7: dout <= 8'b11111111; // 3575 : 255 - 0xff
      12'hDF8: dout <= 8'b11111111; // 3576 : 255 - 0xff -- plane 1
      12'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      12'hDFA: dout <= 8'b11111111; // 3578 : 255 - 0xff
      12'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout <= 8'b11111111; // 3580 : 255 - 0xff
      12'hDFD: dout <= 8'b11111111; // 3581 : 255 - 0xff
      12'hDFE: dout <= 8'b11111111; // 3582 : 255 - 0xff
      12'hDFF: dout <= 8'b11111111; // 3583 : 255 - 0xff
      12'hE00: dout <= 8'b11111111; // 3584 : 255 - 0xff -- Sprite 0xe0
      12'hE01: dout <= 8'b11111111; // 3585 : 255 - 0xff
      12'hE02: dout <= 8'b11111111; // 3586 : 255 - 0xff
      12'hE03: dout <= 8'b11111111; // 3587 : 255 - 0xff
      12'hE04: dout <= 8'b11111111; // 3588 : 255 - 0xff
      12'hE05: dout <= 8'b11111111; // 3589 : 255 - 0xff
      12'hE06: dout <= 8'b11111111; // 3590 : 255 - 0xff
      12'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      12'hE08: dout <= 8'b11111111; // 3592 : 255 - 0xff -- plane 1
      12'hE09: dout <= 8'b11111111; // 3593 : 255 - 0xff
      12'hE0A: dout <= 8'b11111111; // 3594 : 255 - 0xff
      12'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      12'hE0C: dout <= 8'b11111111; // 3596 : 255 - 0xff
      12'hE0D: dout <= 8'b11111111; // 3597 : 255 - 0xff
      12'hE0E: dout <= 8'b11111111; // 3598 : 255 - 0xff
      12'hE0F: dout <= 8'b11111111; // 3599 : 255 - 0xff
      12'hE10: dout <= 8'b11111111; // 3600 : 255 - 0xff -- Sprite 0xe1
      12'hE11: dout <= 8'b11111111; // 3601 : 255 - 0xff
      12'hE12: dout <= 8'b11111111; // 3602 : 255 - 0xff
      12'hE13: dout <= 8'b11111111; // 3603 : 255 - 0xff
      12'hE14: dout <= 8'b11111111; // 3604 : 255 - 0xff
      12'hE15: dout <= 8'b11111111; // 3605 : 255 - 0xff
      12'hE16: dout <= 8'b11111111; // 3606 : 255 - 0xff
      12'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      12'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout <= 8'b11111111; // 3610 : 255 - 0xff
      12'hE1B: dout <= 8'b11111111; // 3611 : 255 - 0xff
      12'hE1C: dout <= 8'b11111111; // 3612 : 255 - 0xff
      12'hE1D: dout <= 8'b11111111; // 3613 : 255 - 0xff
      12'hE1E: dout <= 8'b11111111; // 3614 : 255 - 0xff
      12'hE1F: dout <= 8'b11111111; // 3615 : 255 - 0xff
      12'hE20: dout <= 8'b11111111; // 3616 : 255 - 0xff -- Sprite 0xe2
      12'hE21: dout <= 8'b11111111; // 3617 : 255 - 0xff
      12'hE22: dout <= 8'b11111111; // 3618 : 255 - 0xff
      12'hE23: dout <= 8'b11111111; // 3619 : 255 - 0xff
      12'hE24: dout <= 8'b11111111; // 3620 : 255 - 0xff
      12'hE25: dout <= 8'b11111111; // 3621 : 255 - 0xff
      12'hE26: dout <= 8'b11111111; // 3622 : 255 - 0xff
      12'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout <= 8'b11111111; // 3624 : 255 - 0xff -- plane 1
      12'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout <= 8'b11111111; // 3626 : 255 - 0xff
      12'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout <= 8'b11111111; // 3628 : 255 - 0xff
      12'hE2D: dout <= 8'b11111111; // 3629 : 255 - 0xff
      12'hE2E: dout <= 8'b11111111; // 3630 : 255 - 0xff
      12'hE2F: dout <= 8'b11111111; // 3631 : 255 - 0xff
      12'hE30: dout <= 8'b11111111; // 3632 : 255 - 0xff -- Sprite 0xe3
      12'hE31: dout <= 8'b11111111; // 3633 : 255 - 0xff
      12'hE32: dout <= 8'b11111111; // 3634 : 255 - 0xff
      12'hE33: dout <= 8'b11111111; // 3635 : 255 - 0xff
      12'hE34: dout <= 8'b11111111; // 3636 : 255 - 0xff
      12'hE35: dout <= 8'b11111111; // 3637 : 255 - 0xff
      12'hE36: dout <= 8'b11111111; // 3638 : 255 - 0xff
      12'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout <= 8'b11111111; // 3640 : 255 - 0xff -- plane 1
      12'hE39: dout <= 8'b11111111; // 3641 : 255 - 0xff
      12'hE3A: dout <= 8'b11111111; // 3642 : 255 - 0xff
      12'hE3B: dout <= 8'b11111111; // 3643 : 255 - 0xff
      12'hE3C: dout <= 8'b11111111; // 3644 : 255 - 0xff
      12'hE3D: dout <= 8'b11111111; // 3645 : 255 - 0xff
      12'hE3E: dout <= 8'b11111111; // 3646 : 255 - 0xff
      12'hE3F: dout <= 8'b11111111; // 3647 : 255 - 0xff
      12'hE40: dout <= 8'b11111111; // 3648 : 255 - 0xff -- Sprite 0xe4
      12'hE41: dout <= 8'b11111111; // 3649 : 255 - 0xff
      12'hE42: dout <= 8'b11111111; // 3650 : 255 - 0xff
      12'hE43: dout <= 8'b11111111; // 3651 : 255 - 0xff
      12'hE44: dout <= 8'b11111111; // 3652 : 255 - 0xff
      12'hE45: dout <= 8'b11111111; // 3653 : 255 - 0xff
      12'hE46: dout <= 8'b11111111; // 3654 : 255 - 0xff
      12'hE47: dout <= 8'b11111111; // 3655 : 255 - 0xff
      12'hE48: dout <= 8'b11111111; // 3656 : 255 - 0xff -- plane 1
      12'hE49: dout <= 8'b11111111; // 3657 : 255 - 0xff
      12'hE4A: dout <= 8'b11111111; // 3658 : 255 - 0xff
      12'hE4B: dout <= 8'b11111111; // 3659 : 255 - 0xff
      12'hE4C: dout <= 8'b11111111; // 3660 : 255 - 0xff
      12'hE4D: dout <= 8'b11111111; // 3661 : 255 - 0xff
      12'hE4E: dout <= 8'b11111111; // 3662 : 255 - 0xff
      12'hE4F: dout <= 8'b11111111; // 3663 : 255 - 0xff
      12'hE50: dout <= 8'b11111111; // 3664 : 255 - 0xff -- Sprite 0xe5
      12'hE51: dout <= 8'b11111111; // 3665 : 255 - 0xff
      12'hE52: dout <= 8'b11111111; // 3666 : 255 - 0xff
      12'hE53: dout <= 8'b11111111; // 3667 : 255 - 0xff
      12'hE54: dout <= 8'b11111111; // 3668 : 255 - 0xff
      12'hE55: dout <= 8'b11111111; // 3669 : 255 - 0xff
      12'hE56: dout <= 8'b11111111; // 3670 : 255 - 0xff
      12'hE57: dout <= 8'b11111111; // 3671 : 255 - 0xff
      12'hE58: dout <= 8'b11111111; // 3672 : 255 - 0xff -- plane 1
      12'hE59: dout <= 8'b11111111; // 3673 : 255 - 0xff
      12'hE5A: dout <= 8'b11111111; // 3674 : 255 - 0xff
      12'hE5B: dout <= 8'b11111111; // 3675 : 255 - 0xff
      12'hE5C: dout <= 8'b11111111; // 3676 : 255 - 0xff
      12'hE5D: dout <= 8'b11111111; // 3677 : 255 - 0xff
      12'hE5E: dout <= 8'b11111111; // 3678 : 255 - 0xff
      12'hE5F: dout <= 8'b11111111; // 3679 : 255 - 0xff
      12'hE60: dout <= 8'b11111111; // 3680 : 255 - 0xff -- Sprite 0xe6
      12'hE61: dout <= 8'b11111111; // 3681 : 255 - 0xff
      12'hE62: dout <= 8'b11111111; // 3682 : 255 - 0xff
      12'hE63: dout <= 8'b11111111; // 3683 : 255 - 0xff
      12'hE64: dout <= 8'b11111111; // 3684 : 255 - 0xff
      12'hE65: dout <= 8'b11111111; // 3685 : 255 - 0xff
      12'hE66: dout <= 8'b11111111; // 3686 : 255 - 0xff
      12'hE67: dout <= 8'b11111111; // 3687 : 255 - 0xff
      12'hE68: dout <= 8'b11111111; // 3688 : 255 - 0xff -- plane 1
      12'hE69: dout <= 8'b11111111; // 3689 : 255 - 0xff
      12'hE6A: dout <= 8'b11111111; // 3690 : 255 - 0xff
      12'hE6B: dout <= 8'b11111111; // 3691 : 255 - 0xff
      12'hE6C: dout <= 8'b11111111; // 3692 : 255 - 0xff
      12'hE6D: dout <= 8'b11111111; // 3693 : 255 - 0xff
      12'hE6E: dout <= 8'b11111111; // 3694 : 255 - 0xff
      12'hE6F: dout <= 8'b11111111; // 3695 : 255 - 0xff
      12'hE70: dout <= 8'b11111111; // 3696 : 255 - 0xff -- Sprite 0xe7
      12'hE71: dout <= 8'b11111111; // 3697 : 255 - 0xff
      12'hE72: dout <= 8'b11111111; // 3698 : 255 - 0xff
      12'hE73: dout <= 8'b11111111; // 3699 : 255 - 0xff
      12'hE74: dout <= 8'b11111111; // 3700 : 255 - 0xff
      12'hE75: dout <= 8'b11111111; // 3701 : 255 - 0xff
      12'hE76: dout <= 8'b11111111; // 3702 : 255 - 0xff
      12'hE77: dout <= 8'b11111111; // 3703 : 255 - 0xff
      12'hE78: dout <= 8'b11111111; // 3704 : 255 - 0xff -- plane 1
      12'hE79: dout <= 8'b11111111; // 3705 : 255 - 0xff
      12'hE7A: dout <= 8'b11111111; // 3706 : 255 - 0xff
      12'hE7B: dout <= 8'b11111111; // 3707 : 255 - 0xff
      12'hE7C: dout <= 8'b11111111; // 3708 : 255 - 0xff
      12'hE7D: dout <= 8'b11111111; // 3709 : 255 - 0xff
      12'hE7E: dout <= 8'b11111111; // 3710 : 255 - 0xff
      12'hE7F: dout <= 8'b11111111; // 3711 : 255 - 0xff
      12'hE80: dout <= 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      12'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      12'hE83: dout <= 8'b11111111; // 3715 : 255 - 0xff
      12'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      12'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout <= 8'b11111111; // 3720 : 255 - 0xff -- plane 1
      12'hE89: dout <= 8'b11111111; // 3721 : 255 - 0xff
      12'hE8A: dout <= 8'b11111111; // 3722 : 255 - 0xff
      12'hE8B: dout <= 8'b11111111; // 3723 : 255 - 0xff
      12'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      12'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      12'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      12'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      12'hE90: dout <= 8'b11111111; // 3728 : 255 - 0xff -- Sprite 0xe9
      12'hE91: dout <= 8'b11111111; // 3729 : 255 - 0xff
      12'hE92: dout <= 8'b11111111; // 3730 : 255 - 0xff
      12'hE93: dout <= 8'b11111111; // 3731 : 255 - 0xff
      12'hE94: dout <= 8'b11111111; // 3732 : 255 - 0xff
      12'hE95: dout <= 8'b11111111; // 3733 : 255 - 0xff
      12'hE96: dout <= 8'b11111111; // 3734 : 255 - 0xff
      12'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff -- plane 1
      12'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout <= 8'b11111111; // 3740 : 255 - 0xff
      12'hE9D: dout <= 8'b11111111; // 3741 : 255 - 0xff
      12'hE9E: dout <= 8'b11111111; // 3742 : 255 - 0xff
      12'hE9F: dout <= 8'b11111111; // 3743 : 255 - 0xff
      12'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      12'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      12'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      12'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      12'hEA4: dout <= 8'b11111111; // 3748 : 255 - 0xff
      12'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      12'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      12'hEA7: dout <= 8'b11111111; // 3751 : 255 - 0xff
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- plane 1
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout <= 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout <= 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Sprite 0xeb
      12'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout <= 8'b11111111; // 3763 : 255 - 0xff
      12'hEB4: dout <= 8'b11111111; // 3764 : 255 - 0xff
      12'hEB5: dout <= 8'b11111111; // 3765 : 255 - 0xff
      12'hEB6: dout <= 8'b11111111; // 3766 : 255 - 0xff
      12'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout <= 8'b11111111; // 3768 : 255 - 0xff -- plane 1
      12'hEB9: dout <= 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout <= 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout <= 8'b11111111; // 3771 : 255 - 0xff
      12'hEBC: dout <= 8'b11111111; // 3772 : 255 - 0xff
      12'hEBD: dout <= 8'b11111111; // 3773 : 255 - 0xff
      12'hEBE: dout <= 8'b11111111; // 3774 : 255 - 0xff
      12'hEBF: dout <= 8'b11111111; // 3775 : 255 - 0xff
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      12'hEC1: dout <= 8'b00000001; // 3777 :   1 - 0x1
      12'hEC2: dout <= 8'b00000011; // 3778 :   3 - 0x3
      12'hEC3: dout <= 8'b00110011; // 3779 :  51 - 0x33
      12'hEC4: dout <= 8'b00011001; // 3780 :  25 - 0x19
      12'hEC5: dout <= 8'b00001111; // 3781 :  15 - 0xf
      12'hEC6: dout <= 8'b00111111; // 3782 :  63 - 0x3f
      12'hEC7: dout <= 8'b00011111; // 3783 :  31 - 0x1f
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b00000001; // 3785 :   1 - 0x1
      12'hECA: dout <= 8'b00000011; // 3786 :   3 - 0x3
      12'hECB: dout <= 8'b00110011; // 3787 :  51 - 0x33
      12'hECC: dout <= 8'b00011001; // 3788 :  25 - 0x19
      12'hECD: dout <= 8'b00001111; // 3789 :  15 - 0xf
      12'hECE: dout <= 8'b00111111; // 3790 :  63 - 0x3f
      12'hECF: dout <= 8'b00011111; // 3791 :  31 - 0x1f
      12'hED0: dout <= 8'b00101011; // 3792 :  43 - 0x2b -- Sprite 0xed
      12'hED1: dout <= 8'b00000111; // 3793 :   7 - 0x7
      12'hED2: dout <= 8'b00000101; // 3794 :   5 - 0x5
      12'hED3: dout <= 8'b00001101; // 3795 :  13 - 0xd
      12'hED4: dout <= 8'b00001011; // 3796 :  11 - 0xb
      12'hED5: dout <= 8'b00011011; // 3797 :  27 - 0x1b
      12'hED6: dout <= 8'b00011011; // 3798 :  27 - 0x1b
      12'hED7: dout <= 8'b00111011; // 3799 :  59 - 0x3b
      12'hED8: dout <= 8'b00101011; // 3800 :  43 - 0x2b -- plane 1
      12'hED9: dout <= 8'b00000111; // 3801 :   7 - 0x7
      12'hEDA: dout <= 8'b00000101; // 3802 :   5 - 0x5
      12'hEDB: dout <= 8'b00001101; // 3803 :  13 - 0xd
      12'hEDC: dout <= 8'b00001011; // 3804 :  11 - 0xb
      12'hEDD: dout <= 8'b00011011; // 3805 :  27 - 0x1b
      12'hEDE: dout <= 8'b00011011; // 3806 :  27 - 0x1b
      12'hEDF: dout <= 8'b00000011; // 3807 :   3 - 0x3
      12'hEE0: dout <= 8'b00001001; // 3808 :   9 - 0x9 -- Sprite 0xee
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000111; // 3810 :   7 - 0x7
      12'hEE3: dout <= 8'b00000111; // 3811 :   7 - 0x7
      12'hEE4: dout <= 8'b00001111; // 3812 :  15 - 0xf
      12'hEE5: dout <= 8'b00001101; // 3813 :  13 - 0xd
      12'hEE6: dout <= 8'b00000001; // 3814 :   1 - 0x1
      12'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      12'hEE8: dout <= 8'b00000001; // 3816 :   1 - 0x1 -- plane 1
      12'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout <= 8'b00000011; // 3818 :   3 - 0x3
      12'hEEB: dout <= 8'b00000101; // 3819 :   5 - 0x5
      12'hEEC: dout <= 8'b00001110; // 3820 :  14 - 0xe
      12'hEED: dout <= 8'b00001101; // 3821 :  13 - 0xd
      12'hEEE: dout <= 8'b00000001; // 3822 :   1 - 0x1
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b11111000; // 3824 : 248 - 0xf8 -- Sprite 0xef
      12'hEF1: dout <= 8'b11111100; // 3825 : 252 - 0xfc
      12'hEF2: dout <= 8'b11111000; // 3826 : 248 - 0xf8
      12'hEF3: dout <= 8'b11101100; // 3827 : 236 - 0xec
      12'hEF4: dout <= 8'b11111000; // 3828 : 248 - 0xf8
      12'hEF5: dout <= 8'b11110000; // 3829 : 240 - 0xf0
      12'hEF6: dout <= 8'b11000000; // 3830 : 192 - 0xc0
      12'hEF7: dout <= 8'b11000000; // 3831 : 192 - 0xc0
      12'hEF8: dout <= 8'b11111000; // 3832 : 248 - 0xf8 -- plane 1
      12'hEF9: dout <= 8'b11111100; // 3833 : 252 - 0xfc
      12'hEFA: dout <= 8'b11000000; // 3834 : 192 - 0xc0
      12'hEFB: dout <= 8'b01000000; // 3835 :  64 - 0x40
      12'hEFC: dout <= 8'b10000000; // 3836 : 128 - 0x80
      12'hEFD: dout <= 8'b10000000; // 3837 : 128 - 0x80
      12'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout <= 8'b10000000; // 3839 : 128 - 0x80
      12'hF00: dout <= 8'b11110000; // 3840 : 240 - 0xf0 -- Sprite 0xf0
      12'hF01: dout <= 8'b11111000; // 3841 : 248 - 0xf8
      12'hF02: dout <= 8'b11111000; // 3842 : 248 - 0xf8
      12'hF03: dout <= 8'b11101000; // 3843 : 232 - 0xe8
      12'hF04: dout <= 8'b11001100; // 3844 : 204 - 0xcc
      12'hF05: dout <= 8'b11100110; // 3845 : 230 - 0xe6
      12'hF06: dout <= 8'b11111011; // 3846 : 251 - 0xfb
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11010000; // 3848 : 208 - 0xd0 -- plane 1
      12'hF09: dout <= 8'b11111000; // 3849 : 248 - 0xf8
      12'hF0A: dout <= 8'b11111000; // 3850 : 248 - 0xf8
      12'hF0B: dout <= 8'b11101000; // 3851 : 232 - 0xe8
      12'hF0C: dout <= 8'b11001100; // 3852 : 204 - 0xcc
      12'hF0D: dout <= 8'b11100110; // 3853 : 230 - 0xe6
      12'hF0E: dout <= 8'b11111000; // 3854 : 248 - 0xf8
      12'hF0F: dout <= 8'b11111110; // 3855 : 254 - 0xfe
      12'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      12'hF11: dout <= 8'b11111110; // 3857 : 254 - 0xfe
      12'hF12: dout <= 8'b11111110; // 3858 : 254 - 0xfe
      12'hF13: dout <= 8'b11111110; // 3859 : 254 - 0xfe
      12'hF14: dout <= 8'b11111110; // 3860 : 254 - 0xfe
      12'hF15: dout <= 8'b10001111; // 3861 : 143 - 0x8f
      12'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b11111110; // 3864 : 254 - 0xfe -- plane 1
      12'hF19: dout <= 8'b11111110; // 3865 : 254 - 0xfe
      12'hF1A: dout <= 8'b00000110; // 3866 :   6 - 0x6
      12'hF1B: dout <= 8'b11111000; // 3867 : 248 - 0xf8
      12'hF1C: dout <= 8'b00001110; // 3868 :  14 - 0xe
      12'hF1D: dout <= 8'b10000000; // 3869 : 128 - 0x80
      12'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout <= 8'b00000001; // 3872 :   1 - 0x1 -- Sprite 0xf2
      12'hF21: dout <= 8'b00001111; // 3873 :  15 - 0xf
      12'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout <= 8'b00000100; // 3876 :   4 - 0x4
      12'hF25: dout <= 8'b00011110; // 3877 :  30 - 0x1e
      12'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout <= 8'b00000011; // 3879 :   3 - 0x3
      12'hF28: dout <= 8'b00000001; // 3880 :   1 - 0x1 -- plane 1
      12'hF29: dout <= 8'b00001111; // 3881 :  15 - 0xf
      12'hF2A: dout <= 8'b00000111; // 3882 :   7 - 0x7
      12'hF2B: dout <= 8'b00011101; // 3883 :  29 - 0x1d
      12'hF2C: dout <= 8'b00111011; // 3884 :  59 - 0x3b
      12'hF2D: dout <= 8'b00000001; // 3885 :   1 - 0x1
      12'hF2E: dout <= 8'b00001111; // 3886 :  15 - 0xf
      12'hF2F: dout <= 8'b00000010; // 3887 :   2 - 0x2
      12'hF30: dout <= 8'b00000111; // 3888 :   7 - 0x7 -- Sprite 0xf3
      12'hF31: dout <= 8'b00001111; // 3889 :  15 - 0xf
      12'hF32: dout <= 8'b00011111; // 3890 :  31 - 0x1f
      12'hF33: dout <= 8'b00001111; // 3891 :  15 - 0xf
      12'hF34: dout <= 8'b00000111; // 3892 :   7 - 0x7
      12'hF35: dout <= 8'b00001111; // 3893 :  15 - 0xf
      12'hF36: dout <= 8'b00001111; // 3894 :  15 - 0xf
      12'hF37: dout <= 8'b00000011; // 3895 :   3 - 0x3
      12'hF38: dout <= 8'b00000010; // 3896 :   2 - 0x2 -- plane 1
      12'hF39: dout <= 8'b00000011; // 3897 :   3 - 0x3
      12'hF3A: dout <= 8'b00000010; // 3898 :   2 - 0x2
      12'hF3B: dout <= 8'b01110111; // 3899 : 119 - 0x77
      12'hF3C: dout <= 8'b00010111; // 3900 :  23 - 0x17
      12'hF3D: dout <= 8'b00000001; // 3901 :   1 - 0x1
      12'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout <= 8'b11100000; // 3904 : 224 - 0xe0 -- Sprite 0xf4
      12'hF41: dout <= 8'b11110000; // 3905 : 240 - 0xf0
      12'hF42: dout <= 8'b11110000; // 3906 : 240 - 0xf0
      12'hF43: dout <= 8'b01001000; // 3907 :  72 - 0x48
      12'hF44: dout <= 8'b11001000; // 3908 : 200 - 0xc8
      12'hF45: dout <= 8'b10011100; // 3909 : 156 - 0x9c
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b11110000; // 3911 : 240 - 0xf0
      12'hF48: dout <= 8'b11100000; // 3912 : 224 - 0xe0 -- plane 1
      12'hF49: dout <= 8'b11110000; // 3913 : 240 - 0xf0
      12'hF4A: dout <= 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout <= 8'b10110000; // 3915 : 176 - 0xb0
      12'hF4C: dout <= 8'b00110000; // 3916 :  48 - 0x30
      12'hF4D: dout <= 8'b01100000; // 3917 :  96 - 0x60
      12'hF4E: dout <= 8'b11110000; // 3918 : 240 - 0xf0
      12'hF4F: dout <= 8'b00010000; // 3919 :  16 - 0x10
      12'hF50: dout <= 8'b11111000; // 3920 : 248 - 0xf8 -- Sprite 0xf5
      12'hF51: dout <= 8'b11111100; // 3921 : 252 - 0xfc
      12'hF52: dout <= 8'b11111100; // 3922 : 252 - 0xfc
      12'hF53: dout <= 8'b11111000; // 3923 : 248 - 0xf8
      12'hF54: dout <= 8'b11111000; // 3924 : 248 - 0xf8
      12'hF55: dout <= 8'b01111000; // 3925 : 120 - 0x78
      12'hF56: dout <= 8'b01110000; // 3926 : 112 - 0x70
      12'hF57: dout <= 8'b01100000; // 3927 :  96 - 0x60
      12'hF58: dout <= 8'b00110000; // 3928 :  48 - 0x30 -- plane 1
      12'hF59: dout <= 8'b11110000; // 3929 : 240 - 0xf0
      12'hF5A: dout <= 8'b11010000; // 3930 : 208 - 0xd0
      12'hF5B: dout <= 8'b11111100; // 3931 : 252 - 0xfc
      12'hF5C: dout <= 8'b11111110; // 3932 : 254 - 0xfe
      12'hF5D: dout <= 8'b00001000; // 3933 :   8 - 0x8
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b01111100; // 3938 : 124 - 0x7c
      12'hF63: dout <= 8'b10001010; // 3939 : 138 - 0x8a
      12'hF64: dout <= 8'b11111110; // 3940 : 254 - 0xfe
      12'hF65: dout <= 8'b11111110; // 3941 : 254 - 0xfe
      12'hF66: dout <= 8'b11111110; // 3942 : 254 - 0xfe
      12'hF67: dout <= 8'b11111110; // 3943 : 254 - 0xfe
      12'hF68: dout <= 8'b00000000; // 3944 :   0 - 0x0 -- plane 1
      12'hF69: dout <= 8'b00010000; // 3945 :  16 - 0x10
      12'hF6A: dout <= 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout <= 8'b01110100; // 3947 : 116 - 0x74
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout <= 8'b11111110; // 3952 : 254 - 0xfe -- Sprite 0xf7
      12'hF71: dout <= 8'b01111100; // 3953 : 124 - 0x7c
      12'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout <= 8'b00000000; // 3960 :   0 - 0x0 -- plane 1
      12'hF79: dout <= 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout <= 8'b00010000; // 3962 :  16 - 0x10
      12'hF7B: dout <= 8'b00010000; // 3963 :  16 - 0x10
      12'hF7C: dout <= 8'b00010000; // 3964 :  16 - 0x10
      12'hF7D: dout <= 8'b00010000; // 3965 :  16 - 0x10
      12'hF7E: dout <= 8'b00010000; // 3966 :  16 - 0x10
      12'hF7F: dout <= 8'b00010000; // 3967 :  16 - 0x10
      12'hF80: dout <= 8'b00000111; // 3968 :   7 - 0x7 -- Sprite 0xf8
      12'hF81: dout <= 8'b00001011; // 3969 :  11 - 0xb
      12'hF82: dout <= 8'b00001111; // 3970 :  15 - 0xf
      12'hF83: dout <= 8'b00001011; // 3971 :  11 - 0xb
      12'hF84: dout <= 8'b00001011; // 3972 :  11 - 0xb
      12'hF85: dout <= 8'b00001011; // 3973 :  11 - 0xb
      12'hF86: dout <= 8'b00001011; // 3974 :  11 - 0xb
      12'hF87: dout <= 8'b00000111; // 3975 :   7 - 0x7
      12'hF88: dout <= 8'b00000000; // 3976 :   0 - 0x0 -- plane 1
      12'hF89: dout <= 8'b00000100; // 3977 :   4 - 0x4
      12'hF8A: dout <= 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout <= 8'b00010100; // 3979 :  20 - 0x14
      12'hF8C: dout <= 8'b00000100; // 3980 :   4 - 0x4
      12'hF8D: dout <= 8'b00000100; // 3981 :   4 - 0x4
      12'hF8E: dout <= 8'b00000100; // 3982 :   4 - 0x4
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b11000000; // 3984 : 192 - 0xc0 -- Sprite 0xf9
      12'hF91: dout <= 8'b11100000; // 3985 : 224 - 0xe0
      12'hF92: dout <= 8'b11100000; // 3986 : 224 - 0xe0
      12'hF93: dout <= 8'b11100000; // 3987 : 224 - 0xe0
      12'hF94: dout <= 8'b11100000; // 3988 : 224 - 0xe0
      12'hF95: dout <= 8'b11100000; // 3989 : 224 - 0xe0
      12'hF96: dout <= 8'b11100000; // 3990 : 224 - 0xe0
      12'hF97: dout <= 8'b11000000; // 3991 : 192 - 0xc0
      12'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0 -- plane 1
      12'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout <= 8'b00011111; // 3995 :  31 - 0x1f
      12'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b00000011; // 4000 :   3 - 0x3 -- Sprite 0xfa
      12'hFA1: dout <= 8'b00000111; // 4001 :   7 - 0x7
      12'hFA2: dout <= 8'b00000111; // 4002 :   7 - 0x7
      12'hFA3: dout <= 8'b00000111; // 4003 :   7 - 0x7
      12'hFA4: dout <= 8'b00000111; // 4004 :   7 - 0x7
      12'hFA5: dout <= 8'b00000111; // 4005 :   7 - 0x7
      12'hFA6: dout <= 8'b00000111; // 4006 :   7 - 0x7
      12'hFA7: dout <= 8'b00000011; // 4007 :   3 - 0x3
      12'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0 -- plane 1
      12'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout <= 8'b11111000; // 4011 : 248 - 0xf8
      12'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b11100000; // 4016 : 224 - 0xe0 -- Sprite 0xfb
      12'hFB1: dout <= 8'b11010000; // 4017 : 208 - 0xd0
      12'hFB2: dout <= 8'b11010000; // 4018 : 208 - 0xd0
      12'hFB3: dout <= 8'b11010000; // 4019 : 208 - 0xd0
      12'hFB4: dout <= 8'b11010000; // 4020 : 208 - 0xd0
      12'hFB5: dout <= 8'b11110000; // 4021 : 240 - 0xf0
      12'hFB6: dout <= 8'b11010000; // 4022 : 208 - 0xd0
      12'hFB7: dout <= 8'b11100000; // 4023 : 224 - 0xe0
      12'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout <= 8'b00100000; // 4025 :  32 - 0x20
      12'hFBA: dout <= 8'b00100000; // 4026 :  32 - 0x20
      12'hFBB: dout <= 8'b00101000; // 4027 :  40 - 0x28
      12'hFBC: dout <= 8'b00100000; // 4028 :  32 - 0x20
      12'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout <= 8'b00100000; // 4030 :  32 - 0x20
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      12'hFC1: dout <= 8'b00000001; // 4033 :   1 - 0x1
      12'hFC2: dout <= 8'b00010011; // 4034 :  19 - 0x13
      12'hFC3: dout <= 8'b00110111; // 4035 :  55 - 0x37
      12'hFC4: dout <= 8'b00111011; // 4036 :  59 - 0x3b
      12'hFC5: dout <= 8'b01110100; // 4037 : 116 - 0x74
      12'hFC6: dout <= 8'b01111010; // 4038 : 122 - 0x7a
      12'hFC7: dout <= 8'b00111110; // 4039 :  62 - 0x3e
      12'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0 -- plane 1
      12'hFC9: dout <= 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout <= 8'b00001000; // 4042 :   8 - 0x8
      12'hFCB: dout <= 8'b00100101; // 4043 :  37 - 0x25
      12'hFCC: dout <= 8'b00010010; // 4044 :  18 - 0x12
      12'hFCD: dout <= 8'b01010011; // 4045 :  83 - 0x53
      12'hFCE: dout <= 8'b00110011; // 4046 :  51 - 0x33
      12'hFCF: dout <= 8'b00111001; // 4047 :  57 - 0x39
      12'hFD0: dout <= 8'b11011000; // 4048 : 216 - 0xd8 -- Sprite 0xfd
      12'hFD1: dout <= 8'b10011000; // 4049 : 152 - 0x98
      12'hFD2: dout <= 8'b10101000; // 4050 : 168 - 0xa8
      12'hFD3: dout <= 8'b11011000; // 4051 : 216 - 0xd8
      12'hFD4: dout <= 8'b11011010; // 4052 : 218 - 0xda
      12'hFD5: dout <= 8'b01110100; // 4053 : 116 - 0x74
      12'hFD6: dout <= 8'b00101000; // 4054 :  40 - 0x28
      12'hFD7: dout <= 8'b11001000; // 4055 : 200 - 0xc8
      12'hFD8: dout <= 8'b00001000; // 4056 :   8 - 0x8 -- plane 1
      12'hFD9: dout <= 8'b10000000; // 4057 : 128 - 0x80
      12'hFDA: dout <= 8'b00110000; // 4058 :  48 - 0x30
      12'hFDB: dout <= 8'b10011100; // 4059 : 156 - 0x9c
      12'hFDC: dout <= 8'b11001010; // 4060 : 202 - 0xca
      12'hFDD: dout <= 8'b10111000; // 4061 : 184 - 0xb8
      12'hFDE: dout <= 8'b10011000; // 4062 : 152 - 0x98
      12'hFDF: dout <= 8'b01111000; // 4063 : 120 - 0x78
      12'hFE0: dout <= 8'b00001000; // 4064 :   8 - 0x8 -- Sprite 0xfe
      12'hFE1: dout <= 8'b01011001; // 4065 :  89 - 0x59
      12'hFE2: dout <= 8'b00110000; // 4066 :  48 - 0x30
      12'hFE3: dout <= 8'b01110001; // 4067 : 113 - 0x71
      12'hFE4: dout <= 8'b01111001; // 4068 : 121 - 0x79
      12'hFE5: dout <= 8'b00101011; // 4069 :  43 - 0x2b
      12'hFE6: dout <= 8'b00110110; // 4070 :  54 - 0x36
      12'hFE7: dout <= 8'b00010110; // 4071 :  22 - 0x16
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- plane 1
      12'hFE9: dout <= 8'b00001000; // 4073 :   8 - 0x8
      12'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout <= 8'b01000000; // 4075 :  64 - 0x40
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b00110001; // 4077 :  49 - 0x31
      12'hFEE: dout <= 8'b00111101; // 4078 :  61 - 0x3d
      12'hFEF: dout <= 8'b00011001; // 4079 :  25 - 0x19
      12'hFF0: dout <= 8'b11000110; // 4080 : 198 - 0xc6 -- Sprite 0xff
      12'hFF1: dout <= 8'b11000100; // 4081 : 196 - 0xc4
      12'hFF2: dout <= 8'b11001100; // 4082 : 204 - 0xcc
      12'hFF3: dout <= 8'b11001100; // 4083 : 204 - 0xcc
      12'hFF4: dout <= 8'b10111000; // 4084 : 184 - 0xb8
      12'hFF5: dout <= 8'b01111100; // 4085 : 124 - 0x7c
      12'hFF6: dout <= 8'b11101100; // 4086 : 236 - 0xec
      12'hFF7: dout <= 8'b11001000; // 4087 : 200 - 0xc8
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout <= 8'b10000000; // 4089 : 128 - 0x80
      12'hFFA: dout <= 8'b11000000; // 4090 : 192 - 0xc0
      12'hFFB: dout <= 8'b11000000; // 4091 : 192 - 0xc0
      12'hFFC: dout <= 8'b11000000; // 4092 : 192 - 0xc0
      12'hFFD: dout <= 8'b10001000; // 4093 : 136 - 0x88
      12'hFFE: dout <= 8'b10111000; // 4094 : 184 - 0xb8
      12'hFFF: dout <= 8'b10111000; // 4095 : 184 - 0xb8
    endcase
  end

endmodule
